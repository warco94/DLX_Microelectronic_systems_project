
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_syn is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_syn;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SNPS_CLOCK_GATE_HIGH_IF_ID is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic;  TE : in std_logic);

end SNPS_CLOCK_GATE_HIGH_IF_ID;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_IF_ID is

   component CLKGATETST_X1
      port( CK, E, SE : in std_logic;  GCK : out std_logic);
   end component;

begin
   
   latch : CLKGATETST_X1 port map( CK => CLK, E => EN, SE => TE, GCK => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor is

   port( RST : in std_logic;  PC_IN, PC_FAIL, IR_IN : in std_logic_vector (31 
         downto 0);  IR_FAIL : in std_logic_vector (15 downto 0);  WRONG_PRE, 
         RIGHT_PRE : in std_logic;  NPC_OUT, LINK_ADD : out std_logic_vector 
         (31 downto 0);  SEL, TAKEN : out std_logic);

end branch_predictor;

architecture SYN_Behavioral of branch_predictor is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal CACHE_mem_0_1_port, CACHE_mem_0_0_port, CACHE_mem_1_1_port, 
      CACHE_mem_1_0_port, CACHE_mem_2_1_port, CACHE_mem_2_0_port, 
      CACHE_mem_3_1_port, CACHE_mem_3_0_port, CACHE_mem_4_1_port, 
      CACHE_mem_4_0_port, CACHE_mem_5_1_port, CACHE_mem_5_0_port, 
      CACHE_mem_6_1_port, CACHE_mem_6_0_port, CACHE_mem_7_1_port, 
      CACHE_mem_7_0_port, CACHE_mem_8_1_port, CACHE_mem_8_0_port, 
      CACHE_mem_9_1_port, CACHE_mem_9_0_port, CACHE_mem_10_1_port, 
      CACHE_mem_10_0_port, CACHE_mem_11_1_port, CACHE_mem_11_0_port, 
      CACHE_mem_12_1_port, CACHE_mem_12_0_port, CACHE_mem_13_1_port, 
      CACHE_mem_13_0_port, CACHE_mem_14_1_port, CACHE_mem_14_0_port, 
      CACHE_mem_15_1_port, CACHE_mem_15_0_port, CACHE_mem_16_1_port, 
      CACHE_mem_16_0_port, CACHE_mem_17_1_port, CACHE_mem_17_0_port, 
      CACHE_mem_18_1_port, CACHE_mem_18_0_port, CACHE_mem_19_1_port, 
      CACHE_mem_19_0_port, CACHE_mem_20_1_port, CACHE_mem_20_0_port, 
      CACHE_mem_21_1_port, CACHE_mem_21_0_port, CACHE_mem_22_1_port, 
      CACHE_mem_22_0_port, CACHE_mem_23_1_port, CACHE_mem_23_0_port, 
      CACHE_mem_24_1_port, CACHE_mem_24_0_port, CACHE_mem_25_1_port, 
      CACHE_mem_25_0_port, CACHE_mem_26_1_port, CACHE_mem_26_0_port, 
      CACHE_mem_27_1_port, CACHE_mem_27_0_port, CACHE_mem_28_1_port, 
      CACHE_mem_28_0_port, CACHE_mem_29_1_port, CACHE_mem_29_0_port, 
      CACHE_mem_30_1_port, CACHE_mem_30_0_port, CACHE_mem_31_1_port, 
      CACHE_mem_31_0_port, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, 
      N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71
      , N72, N73, N74, N75, N76, N77, N82, N83, N84, N85, N86, N87, N88, N89, 
      N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
      N104, N105, N106, N107, N108, N109, N110, N111, N112, N220, N221, N222, 
      N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, 
      N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, 
      N247, N248, N249, N250, N323, N356, N357, N358, N362, N387, N388, N612, 
      N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, 
      N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, 
      N637, N638, N639, N640, N641, N642, N643, N644, N645, n5, n6, n7, n8, n9,
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n60_port, 
      add_65_carry_2_port, add_65_carry_3_port, add_65_carry_4_port, 
      add_65_carry_5_port, add_65_carry_6_port, add_65_carry_7_port, 
      add_65_carry_8_port, add_65_carry_9_port, add_65_carry_10_port, 
      add_65_carry_11_port, add_65_carry_12_port, add_65_carry_13_port, 
      add_65_carry_14_port, add_65_carry_15_port, add_65_carry_16_port, 
      add_65_carry_17_port, add_65_carry_18_port, add_65_carry_19_port, 
      add_65_carry_20_port, add_65_carry_21_port, add_65_carry_22_port, 
      add_65_carry_23_port, add_65_carry_24_port, add_65_carry_25_port, 
      add_65_carry_26_port, add_65_carry_27_port, add_65_carry_28_port, 
      add_65_carry_29_port, add_65_carry_30_port, add_65_carry_31_port, 
      add_59_n1, add_59_carry_2_port, add_59_carry_3_port, add_59_carry_4_port,
      add_59_carry_5_port, add_59_carry_6_port, add_59_carry_7_port, 
      add_59_carry_8_port, add_59_carry_9_port, add_59_carry_10_port, 
      add_59_carry_11_port, add_59_carry_12_port, add_59_carry_13_port, 
      add_59_carry_14_port, add_59_carry_15_port, add_59_carry_16_port, 
      add_59_carry_17_port, add_59_carry_18_port, add_59_carry_19_port, 
      add_59_carry_20_port, add_59_carry_21_port, add_59_carry_22_port, 
      add_59_carry_23_port, add_59_carry_24_port, add_59_carry_25_port, 
      add_59_carry_26_port, add_59_carry_27_port, add_59_carry_28_port, 
      add_59_carry_29_port, add_59_carry_30_port, add_59_carry_31_port, 
      add_53_aco_n2, add_53_aco_carry_2_port, add_53_aco_carry_3_port, 
      add_53_aco_carry_4_port, add_53_aco_carry_5_port, add_53_aco_carry_6_port
      , add_53_aco_carry_7_port, add_53_aco_carry_8_port, 
      add_53_aco_carry_9_port, add_53_aco_carry_10_port, 
      add_53_aco_carry_11_port, add_53_aco_carry_12_port, 
      add_53_aco_carry_13_port, add_53_aco_carry_14_port, 
      add_53_aco_carry_15_port, add_53_aco_carry_16_port, 
      add_53_aco_carry_17_port, add_53_aco_carry_18_port, 
      add_53_aco_carry_19_port, add_53_aco_carry_20_port, 
      add_53_aco_carry_21_port, add_53_aco_carry_22_port, 
      add_53_aco_carry_23_port, add_53_aco_carry_24_port, 
      add_53_aco_carry_25_port, add_53_aco_carry_26_port, 
      add_53_aco_carry_27_port, add_53_aco_carry_28_port, 
      add_53_aco_carry_29_port, add_53_aco_carry_30_port, 
      add_53_aco_carry_31_port, n62_port, n286, n291, n59_port, n1, n2, n3, n4,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n280, n281, n282, n283, n284, 
      n285, n287, n288, n289, n290, n292, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, 
      n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, 
      n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, 
      n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, 
      n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, 
      n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, 
      n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
      n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, 
      n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
      n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, 
      n5544, n5545, n5546, n5547, n5548, n5549, n_1001, n_1002, n_1003 : 
      std_logic;

begin
   
   NPC_OUT_reg_31_inst : DLH_X1 port map( G => N323, D => n1, Q => NPC_OUT(31))
                           ;
   NPC_OUT_reg_30_inst : DLH_X1 port map( G => N323, D => n2, Q => NPC_OUT(30))
                           ;
   NPC_OUT_reg_29_inst : DLH_X1 port map( G => N323, D => n3, Q => NPC_OUT(29))
                           ;
   NPC_OUT_reg_28_inst : DLH_X1 port map( G => N323, D => n4, Q => NPC_OUT(28))
                           ;
   NPC_OUT_reg_27_inst : DLH_X1 port map( G => N323, D => n20, Q => NPC_OUT(27)
                           );
   NPC_OUT_reg_26_inst : DLH_X1 port map( G => N323, D => n21, Q => NPC_OUT(26)
                           );
   NPC_OUT_reg_25_inst : DLH_X1 port map( G => N323, D => n22, Q => NPC_OUT(25)
                           );
   NPC_OUT_reg_24_inst : DLH_X1 port map( G => N323, D => n23, Q => NPC_OUT(24)
                           );
   NPC_OUT_reg_23_inst : DLH_X1 port map( G => N323, D => n24, Q => NPC_OUT(23)
                           );
   NPC_OUT_reg_22_inst : DLH_X1 port map( G => N323, D => n25, Q => NPC_OUT(22)
                           );
   NPC_OUT_reg_21_inst : DLH_X1 port map( G => N323, D => n26, Q => NPC_OUT(21)
                           );
   NPC_OUT_reg_20_inst : DLH_X1 port map( G => N323, D => n27, Q => NPC_OUT(20)
                           );
   NPC_OUT_reg_19_inst : DLH_X1 port map( G => N323, D => n28, Q => NPC_OUT(19)
                           );
   NPC_OUT_reg_18_inst : DLH_X1 port map( G => N323, D => n29, Q => NPC_OUT(18)
                           );
   NPC_OUT_reg_17_inst : DLH_X1 port map( G => N323, D => n30, Q => NPC_OUT(17)
                           );
   NPC_OUT_reg_16_inst : DLH_X1 port map( G => N323, D => n31, Q => NPC_OUT(16)
                           );
   NPC_OUT_reg_15_inst : DLH_X1 port map( G => N323, D => n32, Q => NPC_OUT(15)
                           );
   NPC_OUT_reg_14_inst : DLH_X1 port map( G => N323, D => n33, Q => NPC_OUT(14)
                           );
   NPC_OUT_reg_13_inst : DLH_X1 port map( G => N323, D => n34, Q => NPC_OUT(13)
                           );
   NPC_OUT_reg_12_inst : DLH_X1 port map( G => N323, D => n35, Q => NPC_OUT(12)
                           );
   NPC_OUT_reg_11_inst : DLH_X1 port map( G => N323, D => n36, Q => NPC_OUT(11)
                           );
   NPC_OUT_reg_10_inst : DLH_X1 port map( G => N323, D => n37, Q => NPC_OUT(10)
                           );
   NPC_OUT_reg_9_inst : DLH_X1 port map( G => N323, D => n38, Q => NPC_OUT(9));
   NPC_OUT_reg_8_inst : DLH_X1 port map( G => N323, D => n39, Q => NPC_OUT(8));
   NPC_OUT_reg_7_inst : DLH_X1 port map( G => N323, D => n40, Q => NPC_OUT(7));
   NPC_OUT_reg_6_inst : DLH_X1 port map( G => N323, D => n41, Q => NPC_OUT(6));
   NPC_OUT_reg_5_inst : DLH_X1 port map( G => N323, D => n42, Q => NPC_OUT(5));
   NPC_OUT_reg_4_inst : DLH_X1 port map( G => N323, D => n43, Q => NPC_OUT(4));
   NPC_OUT_reg_3_inst : DLH_X1 port map( G => N323, D => n44, Q => NPC_OUT(3));
   NPC_OUT_reg_2_inst : DLH_X1 port map( G => N323, D => n45, Q => NPC_OUT(2));
   NPC_OUT_reg_1_inst : DLH_X1 port map( G => N323, D => n46, Q => NPC_OUT(1));
   NPC_OUT_reg_0_inst : DLH_X1 port map( G => N323, D => n60_port, Q => 
                           NPC_OUT(0));
   LINK_ADD_reg_31_inst : DLH_X1 port map( G => N356, D => N388, Q => 
                           LINK_ADD(31));
   LINK_ADD_reg_30_inst : DLH_X1 port map( G => N356, D => N387, Q => 
                           LINK_ADD(30));
   LINK_ADD_reg_29_inst : DLH_X1 port map( G => n5323, D => n58_port, Q => 
                           LINK_ADD(29));
   LINK_ADD_reg_28_inst : DLH_X1 port map( G => n5323, D => n282, Q => 
                           LINK_ADD(28));
   LINK_ADD_reg_27_inst : DLH_X1 port map( G => n5323, D => n57_port, Q => 
                           LINK_ADD(27));
   LINK_ADD_reg_26_inst : DLH_X1 port map( G => n5323, D => n288, Q => 
                           LINK_ADD(26));
   LINK_ADD_reg_25_inst : DLH_X1 port map( G => n5323, D => n56_port, Q => 
                           LINK_ADD(25));
   LINK_ADD_reg_24_inst : DLH_X1 port map( G => n5323, D => n287, Q => 
                           LINK_ADD(24));
   LINK_ADD_reg_23_inst : DLH_X1 port map( G => n5323, D => n55_port, Q => 
                           LINK_ADD(23));
   LINK_ADD_reg_22_inst : DLH_X1 port map( G => n5323, D => n292, Q => 
                           LINK_ADD(22));
   LINK_ADD_reg_21_inst : DLH_X1 port map( G => n5323, D => n54_port, Q => 
                           LINK_ADD(21));
   LINK_ADD_reg_20_inst : DLH_X1 port map( G => n5323, D => n290, Q => 
                           LINK_ADD(20));
   LINK_ADD_reg_19_inst : DLH_X1 port map( G => n5323, D => n53_port, Q => 
                           LINK_ADD(19));
   LINK_ADD_reg_18_inst : DLH_X1 port map( G => n5323, D => n283, Q => 
                           LINK_ADD(18));
   LINK_ADD_reg_17_inst : DLH_X1 port map( G => n5323, D => n52_port, Q => 
                           LINK_ADD(17));
   LINK_ADD_reg_16_inst : DLH_X1 port map( G => n5323, D => n289, Q => 
                           LINK_ADD(16));
   LINK_ADD_reg_15_inst : DLH_X1 port map( G => n5323, D => n51_port, Q => 
                           LINK_ADD(15));
   LINK_ADD_reg_14_inst : DLH_X1 port map( G => n5323, D => n281, Q => 
                           LINK_ADD(14));
   LINK_ADD_reg_13_inst : DLH_X1 port map( G => n5323, D => n50_port, Q => 
                           LINK_ADD(13));
   LINK_ADD_reg_12_inst : DLH_X1 port map( G => n5323, D => n284, Q => 
                           LINK_ADD(12));
   LINK_ADD_reg_11_inst : DLH_X1 port map( G => n5323, D => n49_port, Q => 
                           LINK_ADD(11));
   LINK_ADD_reg_10_inst : DLH_X1 port map( G => n5323, D => n285, Q => 
                           LINK_ADD(10));
   LINK_ADD_reg_9_inst : DLH_X1 port map( G => n5323, D => n48_port, Q => 
                           LINK_ADD(9));
   LINK_ADD_reg_8_inst : DLH_X1 port map( G => n5323, D => n280, Q => 
                           LINK_ADD(8));
   LINK_ADD_reg_7_inst : DLH_X1 port map( G => N356, D => n47_port, Q => 
                           LINK_ADD(7));
   LINK_ADD_reg_6_inst : DLH_X1 port map( G => N356, D => n291, Q => 
                           LINK_ADD(6));
   LINK_ADD_reg_5_inst : DLH_X1 port map( G => N356, D => N362, Q => 
                           LINK_ADD(5));
   LINK_ADD_reg_4_inst : DLH_X1 port map( G => N356, D => n286, Q => 
                           LINK_ADD(4));
   LINK_ADD_reg_3_inst : DLH_X1 port map( G => N356, D => n59_port, Q => 
                           LINK_ADD(3));
   LINK_ADD_reg_2_inst : DLH_X1 port map( G => N356, D => n62_port, Q => 
                           LINK_ADD(2));
   LINK_ADD_reg_1_inst : DLH_X1 port map( G => N356, D => N358, Q => 
                           LINK_ADD(1));
   LINK_ADD_reg_0_inst : DLH_X1 port map( G => N356, D => N357, Q => 
                           LINK_ADD(0));
   CACHE_mem_reg_0_1_inst : DLH_X1 port map( G => N643, D => N645, Q => 
                           CACHE_mem_0_1_port);
   CACHE_mem_reg_0_0_inst : DLH_X1 port map( G => N643, D => N644, Q => 
                           CACHE_mem_0_0_port);
   CACHE_mem_reg_1_1_inst : DLH_X1 port map( G => N642, D => N645, Q => 
                           CACHE_mem_1_1_port);
   CACHE_mem_reg_1_0_inst : DLH_X1 port map( G => N642, D => N644, Q => 
                           CACHE_mem_1_0_port);
   CACHE_mem_reg_2_1_inst : DLH_X1 port map( G => N641, D => N645, Q => 
                           CACHE_mem_2_1_port);
   CACHE_mem_reg_2_0_inst : DLH_X1 port map( G => N641, D => N644, Q => 
                           CACHE_mem_2_0_port);
   CACHE_mem_reg_3_1_inst : DLH_X1 port map( G => N640, D => N645, Q => 
                           CACHE_mem_3_1_port);
   CACHE_mem_reg_3_0_inst : DLH_X1 port map( G => N640, D => N644, Q => 
                           CACHE_mem_3_0_port);
   CACHE_mem_reg_4_1_inst : DLH_X1 port map( G => N639, D => N645, Q => 
                           CACHE_mem_4_1_port);
   CACHE_mem_reg_4_0_inst : DLH_X1 port map( G => N639, D => N644, Q => 
                           CACHE_mem_4_0_port);
   CACHE_mem_reg_5_1_inst : DLH_X1 port map( G => N638, D => N645, Q => 
                           CACHE_mem_5_1_port);
   CACHE_mem_reg_5_0_inst : DLH_X1 port map( G => N638, D => N644, Q => 
                           CACHE_mem_5_0_port);
   CACHE_mem_reg_6_1_inst : DLH_X1 port map( G => N637, D => N645, Q => 
                           CACHE_mem_6_1_port);
   CACHE_mem_reg_6_0_inst : DLH_X1 port map( G => N637, D => N644, Q => 
                           CACHE_mem_6_0_port);
   CACHE_mem_reg_7_1_inst : DLH_X1 port map( G => N636, D => N645, Q => 
                           CACHE_mem_7_1_port);
   CACHE_mem_reg_7_0_inst : DLH_X1 port map( G => N636, D => N644, Q => 
                           CACHE_mem_7_0_port);
   CACHE_mem_reg_8_1_inst : DLH_X1 port map( G => N635, D => N645, Q => 
                           CACHE_mem_8_1_port);
   CACHE_mem_reg_8_0_inst : DLH_X1 port map( G => N635, D => N644, Q => 
                           CACHE_mem_8_0_port);
   CACHE_mem_reg_9_1_inst : DLH_X1 port map( G => N634, D => N645, Q => 
                           CACHE_mem_9_1_port);
   CACHE_mem_reg_9_0_inst : DLH_X1 port map( G => N634, D => N644, Q => 
                           CACHE_mem_9_0_port);
   CACHE_mem_reg_10_1_inst : DLH_X1 port map( G => N633, D => N645, Q => 
                           CACHE_mem_10_1_port);
   CACHE_mem_reg_10_0_inst : DLH_X1 port map( G => N633, D => N644, Q => 
                           CACHE_mem_10_0_port);
   CACHE_mem_reg_11_1_inst : DLH_X1 port map( G => N632, D => N645, Q => 
                           CACHE_mem_11_1_port);
   CACHE_mem_reg_11_0_inst : DLH_X1 port map( G => N632, D => N644, Q => 
                           CACHE_mem_11_0_port);
   CACHE_mem_reg_12_1_inst : DLH_X1 port map( G => N631, D => N645, Q => 
                           CACHE_mem_12_1_port);
   CACHE_mem_reg_12_0_inst : DLH_X1 port map( G => N631, D => N644, Q => 
                           CACHE_mem_12_0_port);
   CACHE_mem_reg_13_1_inst : DLH_X1 port map( G => N630, D => N645, Q => 
                           CACHE_mem_13_1_port);
   CACHE_mem_reg_13_0_inst : DLH_X1 port map( G => N630, D => N644, Q => 
                           CACHE_mem_13_0_port);
   CACHE_mem_reg_14_1_inst : DLH_X1 port map( G => N629, D => N645, Q => 
                           CACHE_mem_14_1_port);
   CACHE_mem_reg_14_0_inst : DLH_X1 port map( G => N629, D => N644, Q => 
                           CACHE_mem_14_0_port);
   CACHE_mem_reg_15_1_inst : DLH_X1 port map( G => N628, D => N645, Q => 
                           CACHE_mem_15_1_port);
   CACHE_mem_reg_15_0_inst : DLH_X1 port map( G => N628, D => N644, Q => 
                           CACHE_mem_15_0_port);
   CACHE_mem_reg_16_1_inst : DLH_X1 port map( G => N627, D => N645, Q => 
                           CACHE_mem_16_1_port);
   CACHE_mem_reg_16_0_inst : DLH_X1 port map( G => N627, D => N644, Q => 
                           CACHE_mem_16_0_port);
   CACHE_mem_reg_17_1_inst : DLH_X1 port map( G => N626, D => N645, Q => 
                           CACHE_mem_17_1_port);
   CACHE_mem_reg_17_0_inst : DLH_X1 port map( G => N626, D => N644, Q => 
                           CACHE_mem_17_0_port);
   CACHE_mem_reg_18_1_inst : DLH_X1 port map( G => N625, D => N645, Q => 
                           CACHE_mem_18_1_port);
   CACHE_mem_reg_18_0_inst : DLH_X1 port map( G => N625, D => N644, Q => 
                           CACHE_mem_18_0_port);
   CACHE_mem_reg_19_1_inst : DLH_X1 port map( G => N624, D => N645, Q => 
                           CACHE_mem_19_1_port);
   CACHE_mem_reg_19_0_inst : DLH_X1 port map( G => N624, D => N644, Q => 
                           CACHE_mem_19_0_port);
   CACHE_mem_reg_20_1_inst : DLH_X1 port map( G => N623, D => N645, Q => 
                           CACHE_mem_20_1_port);
   CACHE_mem_reg_20_0_inst : DLH_X1 port map( G => N623, D => N644, Q => 
                           CACHE_mem_20_0_port);
   CACHE_mem_reg_21_1_inst : DLH_X1 port map( G => N622, D => N645, Q => 
                           CACHE_mem_21_1_port);
   CACHE_mem_reg_21_0_inst : DLH_X1 port map( G => N622, D => N644, Q => 
                           CACHE_mem_21_0_port);
   CACHE_mem_reg_22_1_inst : DLH_X1 port map( G => N621, D => N645, Q => 
                           CACHE_mem_22_1_port);
   CACHE_mem_reg_22_0_inst : DLH_X1 port map( G => N621, D => N644, Q => 
                           CACHE_mem_22_0_port);
   CACHE_mem_reg_23_1_inst : DLH_X1 port map( G => N620, D => N645, Q => 
                           CACHE_mem_23_1_port);
   CACHE_mem_reg_23_0_inst : DLH_X1 port map( G => N620, D => N644, Q => 
                           CACHE_mem_23_0_port);
   CACHE_mem_reg_24_1_inst : DLH_X1 port map( G => N619, D => N645, Q => 
                           CACHE_mem_24_1_port);
   CACHE_mem_reg_24_0_inst : DLH_X1 port map( G => N619, D => N644, Q => 
                           CACHE_mem_24_0_port);
   CACHE_mem_reg_25_1_inst : DLH_X1 port map( G => N618, D => N645, Q => 
                           CACHE_mem_25_1_port);
   CACHE_mem_reg_25_0_inst : DLH_X1 port map( G => N618, D => N644, Q => 
                           CACHE_mem_25_0_port);
   CACHE_mem_reg_26_1_inst : DLH_X1 port map( G => N617, D => N645, Q => 
                           CACHE_mem_26_1_port);
   CACHE_mem_reg_26_0_inst : DLH_X1 port map( G => N617, D => N644, Q => 
                           CACHE_mem_26_0_port);
   CACHE_mem_reg_27_1_inst : DLH_X1 port map( G => N616, D => N645, Q => 
                           CACHE_mem_27_1_port);
   CACHE_mem_reg_27_0_inst : DLH_X1 port map( G => N616, D => N644, Q => 
                           CACHE_mem_27_0_port);
   CACHE_mem_reg_28_1_inst : DLH_X1 port map( G => N615, D => N645, Q => 
                           CACHE_mem_28_1_port);
   CACHE_mem_reg_28_0_inst : DLH_X1 port map( G => N615, D => N644, Q => 
                           CACHE_mem_28_0_port);
   CACHE_mem_reg_29_1_inst : DLH_X1 port map( G => N614, D => N645, Q => 
                           CACHE_mem_29_1_port);
   CACHE_mem_reg_29_0_inst : DLH_X1 port map( G => N614, D => N644, Q => 
                           CACHE_mem_29_0_port);
   CACHE_mem_reg_30_1_inst : DLH_X1 port map( G => N613, D => N645, Q => 
                           CACHE_mem_30_1_port);
   CACHE_mem_reg_30_0_inst : DLH_X1 port map( G => N613, D => N644, Q => 
                           CACHE_mem_30_0_port);
   CACHE_mem_reg_31_1_inst : DLH_X1 port map( G => N612, D => N645, Q => 
                           CACHE_mem_31_1_port);
   CACHE_mem_reg_31_0_inst : DLH_X1 port map( G => N612, D => N644, Q => 
                           CACHE_mem_31_0_port);
   add_65_U1_1 : FA_X1 port map( A => PC_IN(1), B => IR_IN(1), CI => add_59_n1,
                           CO => add_65_carry_2_port, S => N220);
   add_65_U1_2 : FA_X1 port map( A => PC_IN(2), B => IR_IN(2), CI => 
                           add_65_carry_2_port, CO => add_65_carry_3_port, S =>
                           N221);
   add_65_U1_3 : FA_X1 port map( A => PC_IN(3), B => IR_IN(3), CI => 
                           add_65_carry_3_port, CO => add_65_carry_4_port, S =>
                           N222);
   add_65_U1_4 : FA_X1 port map( A => PC_IN(4), B => IR_IN(4), CI => 
                           add_65_carry_4_port, CO => add_65_carry_5_port, S =>
                           N223);
   add_65_U1_5 : FA_X1 port map( A => PC_IN(5), B => IR_IN(5), CI => 
                           add_65_carry_5_port, CO => add_65_carry_6_port, S =>
                           N224);
   add_65_U1_6 : FA_X1 port map( A => PC_IN(6), B => IR_IN(6), CI => 
                           add_65_carry_6_port, CO => add_65_carry_7_port, S =>
                           N225);
   add_65_U1_7 : FA_X1 port map( A => PC_IN(7), B => IR_IN(7), CI => 
                           add_65_carry_7_port, CO => add_65_carry_8_port, S =>
                           N226);
   add_65_U1_8 : FA_X1 port map( A => PC_IN(8), B => IR_IN(8), CI => 
                           add_65_carry_8_port, CO => add_65_carry_9_port, S =>
                           N227);
   add_65_U1_9 : FA_X1 port map( A => PC_IN(9), B => IR_IN(9), CI => 
                           add_65_carry_9_port, CO => add_65_carry_10_port, S 
                           => N228);
   add_65_U1_10 : FA_X1 port map( A => PC_IN(10), B => IR_IN(10), CI => 
                           add_65_carry_10_port, CO => add_65_carry_11_port, S 
                           => N229);
   add_65_U1_11 : FA_X1 port map( A => PC_IN(11), B => IR_IN(11), CI => 
                           add_65_carry_11_port, CO => add_65_carry_12_port, S 
                           => N230);
   add_65_U1_12 : FA_X1 port map( A => PC_IN(12), B => IR_IN(12), CI => 
                           add_65_carry_12_port, CO => add_65_carry_13_port, S 
                           => N231);
   add_65_U1_13 : FA_X1 port map( A => PC_IN(13), B => IR_IN(13), CI => 
                           add_65_carry_13_port, CO => add_65_carry_14_port, S 
                           => N232);
   add_65_U1_14 : FA_X1 port map( A => PC_IN(14), B => IR_IN(14), CI => 
                           add_65_carry_14_port, CO => add_65_carry_15_port, S 
                           => N233);
   add_65_U1_15 : FA_X1 port map( A => PC_IN(15), B => IR_IN(15), CI => 
                           add_65_carry_15_port, CO => add_65_carry_16_port, S 
                           => N234);
   add_65_U1_16 : FA_X1 port map( A => PC_IN(16), B => IR_IN(15), CI => 
                           add_65_carry_16_port, CO => add_65_carry_17_port, S 
                           => N235);
   add_65_U1_17 : FA_X1 port map( A => PC_IN(17), B => IR_IN(15), CI => 
                           add_65_carry_17_port, CO => add_65_carry_18_port, S 
                           => N236);
   add_65_U1_18 : FA_X1 port map( A => PC_IN(18), B => IR_IN(15), CI => 
                           add_65_carry_18_port, CO => add_65_carry_19_port, S 
                           => N237);
   add_65_U1_19 : FA_X1 port map( A => PC_IN(19), B => IR_IN(15), CI => 
                           add_65_carry_19_port, CO => add_65_carry_20_port, S 
                           => N238);
   add_65_U1_20 : FA_X1 port map( A => PC_IN(20), B => IR_IN(15), CI => 
                           add_65_carry_20_port, CO => add_65_carry_21_port, S 
                           => N239);
   add_65_U1_21 : FA_X1 port map( A => PC_IN(21), B => IR_IN(15), CI => 
                           add_65_carry_21_port, CO => add_65_carry_22_port, S 
                           => N240);
   add_65_U1_22 : FA_X1 port map( A => PC_IN(22), B => IR_IN(15), CI => 
                           add_65_carry_22_port, CO => add_65_carry_23_port, S 
                           => N241);
   add_65_U1_23 : FA_X1 port map( A => PC_IN(23), B => IR_IN(15), CI => 
                           add_65_carry_23_port, CO => add_65_carry_24_port, S 
                           => N242);
   add_65_U1_24 : FA_X1 port map( A => PC_IN(24), B => IR_IN(15), CI => 
                           add_65_carry_24_port, CO => add_65_carry_25_port, S 
                           => N243);
   add_65_U1_25 : FA_X1 port map( A => PC_IN(25), B => IR_IN(15), CI => 
                           add_65_carry_25_port, CO => add_65_carry_26_port, S 
                           => N244);
   add_65_U1_26 : FA_X1 port map( A => PC_IN(26), B => IR_IN(15), CI => 
                           add_65_carry_26_port, CO => add_65_carry_27_port, S 
                           => N245);
   add_65_U1_27 : FA_X1 port map( A => PC_IN(27), B => IR_IN(15), CI => 
                           add_65_carry_27_port, CO => add_65_carry_28_port, S 
                           => N246);
   add_65_U1_28 : FA_X1 port map( A => PC_IN(28), B => IR_IN(15), CI => 
                           add_65_carry_28_port, CO => add_65_carry_29_port, S 
                           => N247);
   add_65_U1_29 : FA_X1 port map( A => PC_IN(29), B => IR_IN(15), CI => 
                           add_65_carry_29_port, CO => add_65_carry_30_port, S 
                           => N248);
   add_65_U1_30 : FA_X1 port map( A => PC_IN(30), B => IR_IN(15), CI => 
                           add_65_carry_30_port, CO => add_65_carry_31_port, S 
                           => N249);
   add_65_U1_31 : FA_X1 port map( A => PC_IN(31), B => IR_IN(15), CI => 
                           add_65_carry_31_port, CO => n_1001, S => N250);
   add_59_U1_1 : FA_X1 port map( A => PC_IN(1), B => IR_IN(1), CI => add_59_n1,
                           CO => add_59_carry_2_port, S => N82);
   add_59_U1_2 : FA_X1 port map( A => PC_IN(2), B => IR_IN(2), CI => 
                           add_59_carry_2_port, CO => add_59_carry_3_port, S =>
                           N83);
   add_59_U1_3 : FA_X1 port map( A => PC_IN(3), B => IR_IN(3), CI => 
                           add_59_carry_3_port, CO => add_59_carry_4_port, S =>
                           N84);
   add_59_U1_4 : FA_X1 port map( A => PC_IN(4), B => IR_IN(4), CI => 
                           add_59_carry_4_port, CO => add_59_carry_5_port, S =>
                           N85);
   add_59_U1_5 : FA_X1 port map( A => PC_IN(5), B => IR_IN(5), CI => 
                           add_59_carry_5_port, CO => add_59_carry_6_port, S =>
                           N86);
   add_59_U1_6 : FA_X1 port map( A => PC_IN(6), B => IR_IN(6), CI => 
                           add_59_carry_6_port, CO => add_59_carry_7_port, S =>
                           N87);
   add_59_U1_7 : FA_X1 port map( A => PC_IN(7), B => IR_IN(7), CI => 
                           add_59_carry_7_port, CO => add_59_carry_8_port, S =>
                           N88);
   add_59_U1_8 : FA_X1 port map( A => PC_IN(8), B => IR_IN(8), CI => 
                           add_59_carry_8_port, CO => add_59_carry_9_port, S =>
                           N89);
   add_59_U1_9 : FA_X1 port map( A => PC_IN(9), B => IR_IN(9), CI => 
                           add_59_carry_9_port, CO => add_59_carry_10_port, S 
                           => N90);
   add_59_U1_10 : FA_X1 port map( A => PC_IN(10), B => IR_IN(10), CI => 
                           add_59_carry_10_port, CO => add_59_carry_11_port, S 
                           => N91);
   add_59_U1_11 : FA_X1 port map( A => PC_IN(11), B => IR_IN(11), CI => 
                           add_59_carry_11_port, CO => add_59_carry_12_port, S 
                           => N92);
   add_59_U1_12 : FA_X1 port map( A => PC_IN(12), B => IR_IN(12), CI => 
                           add_59_carry_12_port, CO => add_59_carry_13_port, S 
                           => N93);
   add_59_U1_13 : FA_X1 port map( A => PC_IN(13), B => IR_IN(13), CI => 
                           add_59_carry_13_port, CO => add_59_carry_14_port, S 
                           => N94);
   add_59_U1_14 : FA_X1 port map( A => PC_IN(14), B => IR_IN(14), CI => 
                           add_59_carry_14_port, CO => add_59_carry_15_port, S 
                           => N95);
   add_59_U1_15 : FA_X1 port map( A => PC_IN(15), B => IR_IN(15), CI => 
                           add_59_carry_15_port, CO => add_59_carry_16_port, S 
                           => N96);
   add_59_U1_16 : FA_X1 port map( A => PC_IN(16), B => IR_IN(16), CI => 
                           add_59_carry_16_port, CO => add_59_carry_17_port, S 
                           => N97);
   add_59_U1_17 : FA_X1 port map( A => PC_IN(17), B => IR_IN(17), CI => 
                           add_59_carry_17_port, CO => add_59_carry_18_port, S 
                           => N98);
   add_59_U1_18 : FA_X1 port map( A => PC_IN(18), B => IR_IN(18), CI => 
                           add_59_carry_18_port, CO => add_59_carry_19_port, S 
                           => N99);
   add_59_U1_19 : FA_X1 port map( A => PC_IN(19), B => IR_IN(19), CI => 
                           add_59_carry_19_port, CO => add_59_carry_20_port, S 
                           => N100);
   add_59_U1_20 : FA_X1 port map( A => PC_IN(20), B => IR_IN(20), CI => 
                           add_59_carry_20_port, CO => add_59_carry_21_port, S 
                           => N101);
   add_59_U1_21 : FA_X1 port map( A => PC_IN(21), B => IR_IN(21), CI => 
                           add_59_carry_21_port, CO => add_59_carry_22_port, S 
                           => N102);
   add_59_U1_22 : FA_X1 port map( A => PC_IN(22), B => IR_IN(22), CI => 
                           add_59_carry_22_port, CO => add_59_carry_23_port, S 
                           => N103);
   add_59_U1_23 : FA_X1 port map( A => PC_IN(23), B => IR_IN(23), CI => 
                           add_59_carry_23_port, CO => add_59_carry_24_port, S 
                           => N104);
   add_59_U1_24 : FA_X1 port map( A => PC_IN(24), B => IR_IN(24), CI => 
                           add_59_carry_24_port, CO => add_59_carry_25_port, S 
                           => N105);
   add_59_U1_25 : FA_X1 port map( A => PC_IN(25), B => IR_IN(25), CI => 
                           add_59_carry_25_port, CO => add_59_carry_26_port, S 
                           => N106);
   add_59_U1_26 : FA_X1 port map( A => PC_IN(26), B => IR_IN(25), CI => 
                           add_59_carry_26_port, CO => add_59_carry_27_port, S 
                           => N107);
   add_59_U1_27 : FA_X1 port map( A => PC_IN(27), B => IR_IN(25), CI => 
                           add_59_carry_27_port, CO => add_59_carry_28_port, S 
                           => N108);
   add_59_U1_28 : FA_X1 port map( A => PC_IN(28), B => IR_IN(25), CI => 
                           add_59_carry_28_port, CO => add_59_carry_29_port, S 
                           => N109);
   add_59_U1_29 : FA_X1 port map( A => PC_IN(29), B => IR_IN(25), CI => 
                           add_59_carry_29_port, CO => add_59_carry_30_port, S 
                           => N110);
   add_59_U1_30 : FA_X1 port map( A => PC_IN(30), B => IR_IN(25), CI => 
                           add_59_carry_30_port, CO => add_59_carry_31_port, S 
                           => N111);
   add_59_U1_31 : FA_X1 port map( A => PC_IN(31), B => IR_IN(25), CI => 
                           add_59_carry_31_port, CO => n_1002, S => N112);
   add_53_aco_U1_1 : FA_X1 port map( A => PC_FAIL(1), B => n6, CI => 
                           add_53_aco_n2, CO => add_53_aco_carry_2_port, S => 
                           N47);
   add_53_aco_U1_2 : FA_X1 port map( A => PC_FAIL(2), B => n8, CI => 
                           add_53_aco_carry_2_port, CO => 
                           add_53_aco_carry_3_port, S => N48);
   add_53_aco_U1_3 : FA_X1 port map( A => PC_FAIL(3), B => n9, CI => 
                           add_53_aco_carry_3_port, CO => 
                           add_53_aco_carry_4_port, S => N49);
   add_53_aco_U1_4 : FA_X1 port map( A => PC_FAIL(4), B => n10, CI => 
                           add_53_aco_carry_4_port, CO => 
                           add_53_aco_carry_5_port, S => N50);
   add_53_aco_U1_5 : FA_X1 port map( A => PC_FAIL(5), B => n7, CI => 
                           add_53_aco_carry_5_port, CO => 
                           add_53_aco_carry_6_port, S => N51);
   add_53_aco_U1_6 : FA_X1 port map( A => PC_FAIL(6), B => n11, CI => 
                           add_53_aco_carry_6_port, CO => 
                           add_53_aco_carry_7_port, S => N52);
   add_53_aco_U1_7 : FA_X1 port map( A => PC_FAIL(7), B => n12, CI => 
                           add_53_aco_carry_7_port, CO => 
                           add_53_aco_carry_8_port, S => N53);
   add_53_aco_U1_8 : FA_X1 port map( A => PC_FAIL(8), B => n13, CI => 
                           add_53_aco_carry_8_port, CO => 
                           add_53_aco_carry_9_port, S => N54);
   add_53_aco_U1_9 : FA_X1 port map( A => PC_FAIL(9), B => n14, CI => 
                           add_53_aco_carry_9_port, CO => 
                           add_53_aco_carry_10_port, S => N55);
   add_53_aco_U1_10 : FA_X1 port map( A => PC_FAIL(10), B => n15, CI => 
                           add_53_aco_carry_10_port, CO => 
                           add_53_aco_carry_11_port, S => N56);
   add_53_aco_U1_11 : FA_X1 port map( A => PC_FAIL(11), B => n16, CI => 
                           add_53_aco_carry_11_port, CO => 
                           add_53_aco_carry_12_port, S => N57);
   add_53_aco_U1_12 : FA_X1 port map( A => PC_FAIL(12), B => n17, CI => 
                           add_53_aco_carry_12_port, CO => 
                           add_53_aco_carry_13_port, S => N58);
   add_53_aco_U1_13 : FA_X1 port map( A => PC_FAIL(13), B => n18, CI => 
                           add_53_aco_carry_13_port, CO => 
                           add_53_aco_carry_14_port, S => N59);
   add_53_aco_U1_14 : FA_X1 port map( A => PC_FAIL(14), B => n19, CI => 
                           add_53_aco_carry_14_port, CO => 
                           add_53_aco_carry_15_port, S => N60);
   add_53_aco_U1_15 : FA_X1 port map( A => PC_FAIL(15), B => n5, CI => 
                           add_53_aco_carry_15_port, CO => 
                           add_53_aco_carry_16_port, S => N61);
   add_53_aco_U1_16 : FA_X1 port map( A => PC_FAIL(16), B => n5, CI => 
                           add_53_aco_carry_16_port, CO => 
                           add_53_aco_carry_17_port, S => N62);
   add_53_aco_U1_17 : FA_X1 port map( A => PC_FAIL(17), B => n5, CI => 
                           add_53_aco_carry_17_port, CO => 
                           add_53_aco_carry_18_port, S => N63);
   add_53_aco_U1_18 : FA_X1 port map( A => PC_FAIL(18), B => n5, CI => 
                           add_53_aco_carry_18_port, CO => 
                           add_53_aco_carry_19_port, S => N64);
   add_53_aco_U1_19 : FA_X1 port map( A => PC_FAIL(19), B => n5, CI => 
                           add_53_aco_carry_19_port, CO => 
                           add_53_aco_carry_20_port, S => N65);
   add_53_aco_U1_20 : FA_X1 port map( A => PC_FAIL(20), B => n5, CI => 
                           add_53_aco_carry_20_port, CO => 
                           add_53_aco_carry_21_port, S => N66);
   add_53_aco_U1_21 : FA_X1 port map( A => PC_FAIL(21), B => n5, CI => 
                           add_53_aco_carry_21_port, CO => 
                           add_53_aco_carry_22_port, S => N67);
   add_53_aco_U1_22 : FA_X1 port map( A => PC_FAIL(22), B => n5, CI => 
                           add_53_aco_carry_22_port, CO => 
                           add_53_aco_carry_23_port, S => N68);
   add_53_aco_U1_23 : FA_X1 port map( A => PC_FAIL(23), B => n5, CI => 
                           add_53_aco_carry_23_port, CO => 
                           add_53_aco_carry_24_port, S => N69);
   add_53_aco_U1_24 : FA_X1 port map( A => PC_FAIL(24), B => n5, CI => 
                           add_53_aco_carry_24_port, CO => 
                           add_53_aco_carry_25_port, S => N70);
   add_53_aco_U1_25 : FA_X1 port map( A => PC_FAIL(25), B => n5, CI => 
                           add_53_aco_carry_25_port, CO => 
                           add_53_aco_carry_26_port, S => N71);
   add_53_aco_U1_26 : FA_X1 port map( A => PC_FAIL(26), B => n5, CI => 
                           add_53_aco_carry_26_port, CO => 
                           add_53_aco_carry_27_port, S => N72);
   add_53_aco_U1_27 : FA_X1 port map( A => PC_FAIL(27), B => n5, CI => 
                           add_53_aco_carry_27_port, CO => 
                           add_53_aco_carry_28_port, S => N73);
   add_53_aco_U1_28 : FA_X1 port map( A => PC_FAIL(28), B => n5, CI => 
                           add_53_aco_carry_28_port, CO => 
                           add_53_aco_carry_29_port, S => N74);
   add_53_aco_U1_29 : FA_X1 port map( A => PC_FAIL(29), B => n5, CI => 
                           add_53_aco_carry_29_port, CO => 
                           add_53_aco_carry_30_port, S => N75);
   add_53_aco_U1_30 : FA_X1 port map( A => PC_FAIL(30), B => n5, CI => 
                           add_53_aco_carry_30_port, CO => 
                           add_53_aco_carry_31_port, S => N76);
   add_53_aco_U1_31 : FA_X1 port map( A => PC_FAIL(31), B => n5, CI => 
                           add_53_aco_carry_31_port, CO => n_1003, S => N77);
   U3 : NAND2_X1 port map( A1 => n5320, A2 => n5455, ZN => N323);
   U4 : AOI21_X1 port map( B1 => n5451, B2 => RIGHT_PRE, A => n5548, ZN => 
                           n5400);
   U5 : INV_X1 port map( A => n5516, ZN => n5319);
   U6 : NAND2_X1 port map( A1 => n5515, A2 => n5319, ZN => n5321);
   U7 : NOR2_X2 port map( A1 => n5325, A2 => n5454, ZN => N645);
   U8 : INV_X2 port map( A => n5321, ZN => n5320);
   U9 : NOR2_X2 port map( A1 => n5465, A2 => n5451, ZN => N644);
   U10 : INV_X2 port map( A => n5465, ZN => n5548);
   U11 : NOR3_X2 port map( A1 => n5373, A2 => n5376, A3 => n5375, ZN => n5429);
   U12 : AOI211_X4 port map( C1 => n5449, C2 => n5448, A => n5447, B => n5446, 
                           ZN => n5467);
   U13 : BUF_X1 port map( A => N356, Z => n5323);
   U14 : INV_X1 port map( A => n5429, ZN => n5405);
   U15 : OAI221_X1 port map( B1 => n5324, B2 => n5515, C1 => n5324, C2 => n5455
                           , A => n5465, ZN => SEL);
   U16 : BUF_X1 port map( A => n5547, Z => n5322);
   U17 : NOR2_X1 port map( A1 => n5516, A2 => n5515, ZN => n5547);
   U18 : INV_X1 port map( A => PC_FAIL(2), ZN => n5375);
   U19 : INV_X1 port map( A => PC_FAIL(5), ZN => n5430);
   U20 : INV_X1 port map( A => PC_FAIL(3), ZN => n5376);
   U21 : INV_X1 port map( A => RST, ZN => n5324);
   U22 : INV_X1 port map( A => RST, ZN => n5325);
   U23 : INV_X1 port map( A => IR_IN(28), ZN => n5326);
   U24 : INV_X1 port map( A => n5457, ZN => n5461);
   U25 : AND2_X2 port map( A1 => n5467, A2 => IR_FAIL(15), ZN => n5);
   U26 : INV_X1 port map( A => PC_FAIL(6), ZN => n5431);
   U27 : NOR2_X1 port map( A1 => PC_FAIL(4), A2 => n5374, ZN => n5436);
   U28 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(30), A3 => IR_IN(31), 
                           ZN => n5365);
   U29 : NAND3_X1 port map( A1 => n5365, A2 => IR_IN(27), A3 => n5326, ZN => 
                           n5515);
   U30 : INV_X1 port map( A => WRONG_PRE, ZN => n5453);
   U31 : NAND2_X1 port map( A1 => RST, A2 => n5453, ZN => n5516);
   U32 : NAND2_X1 port map( A1 => PC_IN(3), A2 => PC_IN(2), ZN => n5457);
   U33 : INV_X1 port map( A => PC_IN(4), ZN => n5456);
   U34 : INV_X1 port map( A => PC_IN(5), ZN => n5368);
   U35 : NOR2_X1 port map( A1 => n5456, A2 => n5368, ZN => n5343);
   U36 : NAND2_X1 port map( A1 => n5461, A2 => n5343, ZN => n5460);
   U37 : INV_X1 port map( A => n5460, ZN => n5366);
   U38 : NAND2_X1 port map( A1 => n5366, A2 => PC_IN(6), ZN => n5514);
   U39 : INV_X1 port map( A => n5514, ZN => n5458);
   U40 : AOI21_X1 port map( B1 => CACHE_mem_31_1_port, B2 => n5458, A => 
                           IR_IN(27), ZN => n5364);
   U41 : NOR2_X1 port map( A1 => PC_IN(5), A2 => n5456, ZN => n5351);
   U42 : AND2_X1 port map( A1 => CACHE_mem_21_1_port, A2 => n5351, ZN => n5327)
                           ;
   U43 : INV_X1 port map( A => PC_IN(6), ZN => n5459);
   U44 : AOI211_X1 port map( C1 => n5343, C2 => CACHE_mem_29_1_port, A => n5327
                           , B => n5459, ZN => n5334);
   U45 : NOR2_X1 port map( A1 => PC_IN(4), A2 => n5368, ZN => n5350);
   U46 : NOR2_X1 port map( A1 => PC_IN(4), A2 => PC_IN(5), ZN => n5352);
   U47 : AOI22_X1 port map( A1 => CACHE_mem_25_1_port, A2 => n5350, B1 => 
                           CACHE_mem_17_1_port, B2 => n5352, ZN => n5333);
   U48 : INV_X1 port map( A => CACHE_mem_5_1_port, ZN => n5330);
   U49 : INV_X1 port map( A => n5351, ZN => n5329);
   U50 : AOI22_X1 port map( A1 => n5343, A2 => CACHE_mem_13_1_port, B1 => 
                           CACHE_mem_9_1_port, B2 => n5350, ZN => n5328);
   U51 : OAI211_X1 port map( C1 => n5330, C2 => n5329, A => n5328, B => n5459, 
                           ZN => n5331);
   U52 : AOI21_X1 port map( B1 => CACHE_mem_1_1_port, B2 => n5352, A => n5331, 
                           ZN => n5332);
   U53 : AOI211_X1 port map( C1 => n5334, C2 => n5333, A => PC_IN(3), B => 
                           n5332, ZN => n5362);
   U54 : AOI22_X1 port map( A1 => n5343, A2 => CACHE_mem_14_1_port, B1 => 
                           CACHE_mem_10_1_port, B2 => n5350, ZN => n5336);
   U55 : AOI22_X1 port map( A1 => CACHE_mem_2_1_port, A2 => n5352, B1 => 
                           CACHE_mem_6_1_port, B2 => n5351, ZN => n5335);
   U56 : INV_X1 port map( A => PC_IN(3), ZN => n5463);
   U57 : AOI21_X1 port map( B1 => n5336, B2 => n5335, A => n5463, ZN => n5340);
   U58 : AOI22_X1 port map( A1 => n5343, A2 => CACHE_mem_12_1_port, B1 => 
                           CACHE_mem_8_1_port, B2 => n5350, ZN => n5338);
   U59 : AOI22_X1 port map( A1 => CACHE_mem_0_1_port, A2 => n5352, B1 => 
                           CACHE_mem_4_1_port, B2 => n5351, ZN => n5337);
   U60 : AOI21_X1 port map( B1 => n5338, B2 => n5337, A => PC_IN(3), ZN => 
                           n5339);
   U61 : NOR2_X1 port map( A1 => n5340, A2 => n5339, ZN => n5349);
   U62 : AOI22_X1 port map( A1 => n5343, A2 => CACHE_mem_30_1_port, B1 => 
                           CACHE_mem_26_1_port, B2 => n5350, ZN => n5342);
   U63 : AOI22_X1 port map( A1 => CACHE_mem_18_1_port, A2 => n5352, B1 => 
                           CACHE_mem_22_1_port, B2 => n5351, ZN => n5341);
   U64 : AOI21_X1 port map( B1 => n5342, B2 => n5341, A => n5463, ZN => n5347);
   U65 : AOI22_X1 port map( A1 => n5343, A2 => CACHE_mem_28_1_port, B1 => 
                           CACHE_mem_24_1_port, B2 => n5350, ZN => n5345);
   U66 : AOI22_X1 port map( A1 => CACHE_mem_20_1_port, A2 => n5351, B1 => 
                           CACHE_mem_16_1_port, B2 => n5352, ZN => n5344);
   U67 : AOI21_X1 port map( B1 => n5345, B2 => n5344, A => PC_IN(3), ZN => 
                           n5346);
   U68 : OAI21_X1 port map( B1 => n5347, B2 => n5346, A => PC_IN(6), ZN => 
                           n5348);
   U69 : OAI21_X1 port map( B1 => PC_IN(6), B2 => n5349, A => n5348, ZN => 
                           n5361);
   U70 : INV_X1 port map( A => PC_IN(2), ZN => n5462);
   U71 : AOI21_X1 port map( B1 => CACHE_mem_23_1_port, B2 => n5351, A => n5459,
                           ZN => n5359);
   U72 : AOI22_X1 port map( A1 => CACHE_mem_27_1_port, A2 => n5350, B1 => 
                           CACHE_mem_19_1_port, B2 => n5352, ZN => n5358);
   U73 : INV_X1 port map( A => CACHE_mem_11_1_port, ZN => n5355);
   U74 : INV_X1 port map( A => n5350, ZN => n5354);
   U75 : AOI22_X1 port map( A1 => CACHE_mem_3_1_port, A2 => n5352, B1 => 
                           CACHE_mem_7_1_port, B2 => n5351, ZN => n5353);
   U76 : OAI211_X1 port map( C1 => n5355, C2 => n5354, A => n5353, B => n5459, 
                           ZN => n5356);
   U77 : AOI22_X1 port map( A1 => n5461, A2 => n5356, B1 => n5366, B2 => 
                           CACHE_mem_15_1_port, ZN => n5357);
   U78 : AOI21_X1 port map( B1 => n5359, B2 => n5358, A => n5357, ZN => n5360);
   U79 : AOI221_X1 port map( B1 => n5362, B2 => PC_IN(2), C1 => n5361, C2 => 
                           n5462, A => n5360, ZN => n5363);
   U80 : NAND4_X1 port map( A1 => n5365, A2 => IR_IN(28), A3 => n5364, A4 => 
                           n5363, ZN => n5455);
   U81 : OAI21_X1 port map( B1 => WRONG_PRE, B2 => n5515, A => RST, ZN => N356)
                           ;
   U82 : AND2_X1 port map( A1 => RST, A2 => PC_IN(0), ZN => N357);
   U83 : AND2_X1 port map( A1 => RST, A2 => PC_IN(1), ZN => N358);
   U84 : NAND2_X1 port map( A1 => n5461, A2 => PC_IN(4), ZN => n5367);
   U85 : AOI211_X1 port map( C1 => n5368, C2 => n5367, A => n5366, B => n5325, 
                           ZN => N362);
   U86 : INV_X1 port map( A => PC_IN(7), ZN => n5513);
   U87 : NOR2_X1 port map( A1 => n5514, A2 => n5513, ZN => n5512);
   U88 : NAND2_X1 port map( A1 => n5512, A2 => PC_IN(8), ZN => n5511);
   U89 : INV_X1 port map( A => PC_IN(9), ZN => n5510);
   U90 : NOR2_X1 port map( A1 => n5511, A2 => n5510, ZN => n5509);
   U91 : NAND2_X1 port map( A1 => n5509, A2 => PC_IN(10), ZN => n5508);
   U92 : INV_X1 port map( A => PC_IN(11), ZN => n5507);
   U93 : NOR2_X1 port map( A1 => n5508, A2 => n5507, ZN => n5506);
   U94 : NAND2_X1 port map( A1 => n5506, A2 => PC_IN(12), ZN => n5505);
   U95 : INV_X1 port map( A => PC_IN(13), ZN => n5504);
   U96 : NOR2_X1 port map( A1 => n5505, A2 => n5504, ZN => n5503);
   U97 : NAND2_X1 port map( A1 => n5503, A2 => PC_IN(14), ZN => n5502);
   U98 : INV_X1 port map( A => PC_IN(15), ZN => n5501);
   U99 : NOR2_X1 port map( A1 => n5502, A2 => n5501, ZN => n5500);
   U100 : NAND2_X1 port map( A1 => n5500, A2 => PC_IN(16), ZN => n5499);
   U101 : INV_X1 port map( A => PC_IN(17), ZN => n5498);
   U102 : NOR2_X1 port map( A1 => n5499, A2 => n5498, ZN => n5497);
   U103 : NAND2_X1 port map( A1 => n5497, A2 => PC_IN(18), ZN => n5496);
   U104 : INV_X1 port map( A => PC_IN(19), ZN => n5495);
   U105 : NOR2_X1 port map( A1 => n5496, A2 => n5495, ZN => n5494);
   U106 : NAND2_X1 port map( A1 => n5494, A2 => PC_IN(20), ZN => n5493);
   U107 : INV_X1 port map( A => PC_IN(21), ZN => n5492);
   U108 : NOR2_X1 port map( A1 => n5493, A2 => n5492, ZN => n5491);
   U109 : NAND2_X1 port map( A1 => n5491, A2 => PC_IN(22), ZN => n5490);
   U110 : INV_X1 port map( A => PC_IN(23), ZN => n5489);
   U111 : NOR2_X1 port map( A1 => n5490, A2 => n5489, ZN => n5488);
   U112 : NAND2_X1 port map( A1 => n5488, A2 => PC_IN(24), ZN => n5487);
   U113 : INV_X1 port map( A => PC_IN(25), ZN => n5486);
   U114 : NOR2_X1 port map( A1 => n5487, A2 => n5486, ZN => n5485);
   U115 : NAND2_X1 port map( A1 => n5485, A2 => PC_IN(26), ZN => n5484);
   U116 : INV_X1 port map( A => PC_IN(27), ZN => n5483);
   U117 : NOR2_X1 port map( A1 => n5484, A2 => n5483, ZN => n5482);
   U118 : NAND2_X1 port map( A1 => n5482, A2 => PC_IN(28), ZN => n5481);
   U119 : INV_X1 port map( A => PC_IN(29), ZN => n5480);
   U120 : NOR2_X1 port map( A1 => n5481, A2 => n5480, ZN => n5479);
   U121 : INV_X1 port map( A => n5479, ZN => n5370);
   U122 : INV_X1 port map( A => PC_IN(30), ZN => n5369);
   U123 : NOR2_X1 port map( A1 => n5370, A2 => n5369, ZN => n5372);
   U124 : AOI211_X1 port map( C1 => n5370, C2 => n5369, A => n5372, B => n5324,
                           ZN => N387);
   U125 : OAI21_X1 port map( B1 => PC_IN(31), B2 => n5372, A => RST, ZN => 
                           n5371);
   U126 : AOI21_X1 port map( B1 => PC_IN(31), B2 => n5372, A => n5371, ZN => 
                           N388);
   U127 : INV_X1 port map( A => PC_FAIL(4), ZN => n5373);
   U128 : NAND3_X1 port map( A1 => n5373, A2 => n5376, A3 => n5375, ZN => n5413
                           );
   U129 : INV_X1 port map( A => n5413, ZN => n5434);
   U130 : NAND3_X1 port map( A1 => n5373, A2 => n5376, A3 => PC_FAIL(2), ZN => 
                           n5411);
   U131 : INV_X1 port map( A => n5411, ZN => n5428);
   U132 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_8_0_port, B1 => n5428
                           , B2 => CACHE_mem_9_0_port, ZN => n5380);
   U133 : NAND3_X1 port map( A1 => n5373, A2 => n5375, A3 => PC_FAIL(3), ZN => 
                           n5410);
   U134 : INV_X1 port map( A => n5410, ZN => n5433);
   U135 : NAND2_X1 port map( A1 => PC_FAIL(3), A2 => PC_FAIL(2), ZN => n5374);
   U136 : AOI22_X1 port map( A1 => n5433, A2 => CACHE_mem_10_0_port, B1 => 
                           n5436, B2 => CACHE_mem_11_0_port, ZN => n5379);
   U137 : NAND3_X1 port map( A1 => n5376, A2 => n5375, A3 => PC_FAIL(4), ZN => 
                           n5408);
   U138 : INV_X1 port map( A => n5408, ZN => n5435);
   U139 : NAND3_X1 port map( A1 => n5375, A2 => PC_FAIL(3), A3 => PC_FAIL(4), 
                           ZN => n5406);
   U140 : INV_X1 port map( A => n5406, ZN => n5438);
   U141 : AOI22_X1 port map( A1 => n5435, A2 => CACHE_mem_12_0_port, B1 => 
                           n5438, B2 => CACHE_mem_14_0_port, ZN => n5378);
   U142 : NAND3_X1 port map( A1 => n5376, A2 => PC_FAIL(4), A3 => PC_FAIL(2), 
                           ZN => n5407);
   U143 : INV_X1 port map( A => n5407, ZN => n5437);
   U144 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_15_0_port, B1 => 
                           n5437, B2 => CACHE_mem_13_0_port, ZN => n5377);
   U145 : NAND4_X1 port map( A1 => n5380, A2 => n5379, A3 => n5378, A4 => n5377
                           , ZN => n5386);
   U146 : AOI22_X1 port map( A1 => n5428, A2 => CACHE_mem_1_0_port, B1 => n5433
                           , B2 => CACHE_mem_2_0_port, ZN => n5384);
   U147 : AOI22_X1 port map( A1 => n5436, A2 => CACHE_mem_3_0_port, B1 => n5438
                           , B2 => CACHE_mem_6_0_port, ZN => n5383);
   U148 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_7_0_port, B1 => n5437
                           , B2 => CACHE_mem_5_0_port, ZN => n5382);
   U149 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_0_0_port, B1 => n5435
                           , B2 => CACHE_mem_4_0_port, ZN => n5381);
   U150 : NAND4_X1 port map( A1 => n5384, A2 => n5383, A3 => n5382, A4 => n5381
                           , ZN => n5385);
   U151 : AOI22_X1 port map( A1 => PC_FAIL(5), A2 => n5386, B1 => n5385, B2 => 
                           n5430, ZN => n5398);
   U152 : AOI22_X1 port map( A1 => n5428, A2 => CACHE_mem_17_0_port, B1 => 
                           n5433, B2 => CACHE_mem_18_0_port, ZN => n5390);
   U153 : AOI22_X1 port map( A1 => n5436, A2 => CACHE_mem_19_0_port, B1 => 
                           n5438, B2 => CACHE_mem_22_0_port, ZN => n5389);
   U154 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_23_0_port, B1 => 
                           n5437, B2 => CACHE_mem_21_0_port, ZN => n5388);
   U155 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_16_0_port, B1 => 
                           n5435, B2 => CACHE_mem_20_0_port, ZN => n5387);
   U156 : NAND4_X1 port map( A1 => n5390, A2 => n5389, A3 => n5388, A4 => n5387
                           , ZN => n5396);
   U157 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_24_0_port, B1 => 
                           n5428, B2 => CACHE_mem_25_0_port, ZN => n5394);
   U158 : AOI22_X1 port map( A1 => n5433, A2 => CACHE_mem_26_0_port, B1 => 
                           n5436, B2 => CACHE_mem_27_0_port, ZN => n5393);
   U159 : AOI22_X1 port map( A1 => n5435, A2 => CACHE_mem_28_0_port, B1 => 
                           n5438, B2 => CACHE_mem_30_0_port, ZN => n5392);
   U160 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_31_0_port, B1 => 
                           n5437, B2 => CACHE_mem_29_0_port, ZN => n5391);
   U161 : NAND4_X1 port map( A1 => n5394, A2 => n5393, A3 => n5392, A4 => n5391
                           , ZN => n5395);
   U162 : OAI221_X1 port map( B1 => PC_FAIL(5), B2 => n5396, C1 => n5430, C2 =>
                           n5395, A => PC_FAIL(6), ZN => n5397);
   U163 : OAI21_X1 port map( B1 => PC_FAIL(6), B2 => n5398, A => n5397, ZN => 
                           n5451);
   U164 : NAND2_X1 port map( A1 => RST, A2 => WRONG_PRE, ZN => n5465);
   U165 : NOR2_X1 port map( A1 => n5400, A2 => n5430, ZN => n5402);
   U166 : NAND2_X1 port map( A1 => PC_FAIL(6), A2 => n5402, ZN => n5399);
   U167 : OAI21_X1 port map( B1 => n5405, B2 => n5399, A => RST, ZN => N612);
   U168 : OAI21_X1 port map( B1 => n5406, B2 => n5399, A => RST, ZN => N613);
   U169 : OAI21_X1 port map( B1 => n5407, B2 => n5399, A => RST, ZN => N614);
   U170 : OAI21_X1 port map( B1 => n5408, B2 => n5399, A => RST, ZN => N615);
   U171 : INV_X1 port map( A => n5436, ZN => n5409);
   U172 : OAI21_X1 port map( B1 => n5409, B2 => n5399, A => RST, ZN => N616);
   U173 : OAI21_X1 port map( B1 => n5410, B2 => n5399, A => RST, ZN => N617);
   U174 : OAI21_X1 port map( B1 => n5411, B2 => n5399, A => RST, ZN => N618);
   U175 : OAI21_X1 port map( B1 => n5413, B2 => n5399, A => RST, ZN => N619);
   U176 : NOR2_X1 port map( A1 => PC_FAIL(5), A2 => n5400, ZN => n5404);
   U177 : NAND2_X1 port map( A1 => PC_FAIL(6), A2 => n5404, ZN => n5401);
   U178 : OAI21_X1 port map( B1 => n5405, B2 => n5401, A => RST, ZN => N620);
   U179 : OAI21_X1 port map( B1 => n5406, B2 => n5401, A => RST, ZN => N621);
   U180 : OAI21_X1 port map( B1 => n5407, B2 => n5401, A => RST, ZN => N622);
   U181 : OAI21_X1 port map( B1 => n5408, B2 => n5401, A => RST, ZN => N623);
   U182 : OAI21_X1 port map( B1 => n5409, B2 => n5401, A => RST, ZN => N624);
   U183 : OAI21_X1 port map( B1 => n5410, B2 => n5401, A => RST, ZN => N625);
   U184 : OAI21_X1 port map( B1 => n5411, B2 => n5401, A => RST, ZN => N626);
   U185 : OAI21_X1 port map( B1 => n5413, B2 => n5401, A => RST, ZN => N627);
   U186 : NAND2_X1 port map( A1 => n5402, A2 => n5431, ZN => n5403);
   U187 : OAI21_X1 port map( B1 => n5405, B2 => n5403, A => RST, ZN => N628);
   U188 : OAI21_X1 port map( B1 => n5406, B2 => n5403, A => RST, ZN => N629);
   U189 : OAI21_X1 port map( B1 => n5407, B2 => n5403, A => RST, ZN => N630);
   U190 : OAI21_X1 port map( B1 => n5408, B2 => n5403, A => RST, ZN => N631);
   U191 : OAI21_X1 port map( B1 => n5409, B2 => n5403, A => RST, ZN => N632);
   U192 : OAI21_X1 port map( B1 => n5410, B2 => n5403, A => RST, ZN => N633);
   U193 : OAI21_X1 port map( B1 => n5411, B2 => n5403, A => RST, ZN => N634);
   U194 : OAI21_X1 port map( B1 => n5413, B2 => n5403, A => RST, ZN => N635);
   U195 : NAND2_X1 port map( A1 => n5404, A2 => n5431, ZN => n5412);
   U196 : OAI21_X1 port map( B1 => n5405, B2 => n5412, A => RST, ZN => N636);
   U197 : OAI21_X1 port map( B1 => n5406, B2 => n5412, A => RST, ZN => N637);
   U198 : OAI21_X1 port map( B1 => n5407, B2 => n5412, A => RST, ZN => N638);
   U199 : OAI21_X1 port map( B1 => n5408, B2 => n5412, A => RST, ZN => N639);
   U200 : OAI21_X1 port map( B1 => n5409, B2 => n5412, A => RST, ZN => N640);
   U201 : OAI21_X1 port map( B1 => n5410, B2 => n5412, A => RST, ZN => N641);
   U202 : OAI21_X1 port map( B1 => n5411, B2 => n5412, A => RST, ZN => N642);
   U203 : OAI21_X1 port map( B1 => n5413, B2 => n5412, A => RST, ZN => N643);
   U204 : AOI22_X1 port map( A1 => n5428, A2 => CACHE_mem_9_1_port, B1 => n5436
                           , B2 => CACHE_mem_11_1_port, ZN => n5449);
   U205 : NOR2_X1 port map( A1 => PC_FAIL(6), A2 => n5430, ZN => n5417);
   U206 : AOI22_X1 port map( A1 => n5438, A2 => CACHE_mem_14_1_port, B1 => 
                           n5437, B2 => CACHE_mem_13_1_port, ZN => n5416);
   U207 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_15_1_port, B1 => 
                           n5434, B2 => CACHE_mem_8_1_port, ZN => n5415);
   U208 : AOI22_X1 port map( A1 => n5433, A2 => CACHE_mem_10_1_port, B1 => 
                           n5435, B2 => CACHE_mem_12_1_port, ZN => n5414);
   U209 : AND4_X1 port map( A1 => n5417, A2 => n5416, A3 => n5415, A4 => n5414,
                           ZN => n5448);
   U210 : AOI211_X1 port map( C1 => n5438, C2 => CACHE_mem_30_1_port, A => 
                           n5430, B => n5431, ZN => n5418);
   U211 : INV_X1 port map( A => n5418, ZN => n5423);
   U212 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_24_1_port, B1 => 
                           n5435, B2 => CACHE_mem_28_1_port, ZN => n5421);
   U213 : AOI22_X1 port map( A1 => n5428, A2 => CACHE_mem_25_1_port, B1 => 
                           n5437, B2 => CACHE_mem_29_1_port, ZN => n5420);
   U214 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_31_1_port, B1 => 
                           n5436, B2 => CACHE_mem_27_1_port, ZN => n5419);
   U215 : NAND3_X1 port map( A1 => n5421, A2 => n5420, A3 => n5419, ZN => n5422
                           );
   U216 : AOI211_X1 port map( C1 => n5433, C2 => CACHE_mem_26_1_port, A => 
                           n5423, B => n5422, ZN => n5447);
   U217 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_16_1_port, B1 => 
                           n5436, B2 => CACHE_mem_19_1_port, ZN => n5424);
   U218 : NAND3_X1 port map( A1 => PC_FAIL(6), A2 => n5424, A3 => n5430, ZN => 
                           n5445);
   U219 : AOI22_X1 port map( A1 => n5428, A2 => CACHE_mem_17_1_port, B1 => 
                           n5433, B2 => CACHE_mem_18_1_port, ZN => n5427);
   U220 : AOI22_X1 port map( A1 => n5435, A2 => CACHE_mem_20_1_port, B1 => 
                           n5438, B2 => CACHE_mem_22_1_port, ZN => n5426);
   U221 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_23_1_port, B1 => 
                           n5437, B2 => CACHE_mem_21_1_port, ZN => n5425);
   U222 : NAND3_X1 port map( A1 => n5427, A2 => n5426, A3 => n5425, ZN => n5444
                           );
   U223 : AOI22_X1 port map( A1 => n5429, A2 => CACHE_mem_7_1_port, B1 => n5428
                           , B2 => CACHE_mem_1_1_port, ZN => n5432);
   U224 : NAND3_X1 port map( A1 => n5432, A2 => n5431, A3 => n5430, ZN => n5443
                           );
   U225 : AOI22_X1 port map( A1 => n5434, A2 => CACHE_mem_0_1_port, B1 => n5433
                           , B2 => CACHE_mem_2_1_port, ZN => n5441);
   U226 : AOI22_X1 port map( A1 => n5436, A2 => CACHE_mem_3_1_port, B1 => n5435
                           , B2 => CACHE_mem_4_1_port, ZN => n5440);
   U227 : AOI22_X1 port map( A1 => n5438, A2 => CACHE_mem_6_1_port, B1 => n5437
                           , B2 => CACHE_mem_5_1_port, ZN => n5439);
   U228 : NAND3_X1 port map( A1 => n5441, A2 => n5440, A3 => n5439, ZN => n5442
                           );
   U229 : OAI22_X1 port map( A1 => n5445, A2 => n5444, B1 => n5443, B2 => n5442
                           , ZN => n5446);
   U230 : NOR2_X1 port map( A1 => n5467, A2 => n5453, ZN => n5450);
   U231 : XNOR2_X1 port map( A => n5451, B => n5450, ZN => n5452);
   U232 : AOI21_X1 port map( B1 => n5467, B2 => n5453, A => n5452, ZN => n5454)
                           ;
   U233 : NOR2_X1 port map( A1 => n5455, A2 => n5321, ZN => TAKEN);
   U234 : AND3_X1 port map( A1 => n5467, A2 => IR_FAIL(0), A3 => PC_FAIL(0), ZN
                           => add_53_aco_n2);
   U235 : AND2_X1 port map( A1 => PC_IN(0), A2 => IR_IN(0), ZN => add_59_n1);
   U236 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(4), ZN => n10);
   U237 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(6), ZN => n11);
   U238 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(7), ZN => n12);
   U239 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(8), ZN => n13);
   U240 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(9), ZN => n14);
   U241 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(10), ZN => n15);
   U242 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(11), ZN => n16);
   U243 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(12), ZN => n17);
   U244 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(13), ZN => n18);
   U245 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(14), ZN => n19);
   U246 : AOI221_X1 port map( B1 => n5461, B2 => PC_IN(4), C1 => n5457, C2 => 
                           n5456, A => n5325, ZN => n286);
   U247 : AOI211_X1 port map( C1 => n5460, C2 => n5459, A => n5458, B => n5324,
                           ZN => n291);
   U248 : AOI211_X1 port map( C1 => n5463, C2 => n5462, A => n5461, B => n5324,
                           ZN => n59_port);
   U249 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(1), ZN => n6);
   U250 : NOR2_X1 port map( A1 => PC_IN(0), A2 => IR_IN(0), ZN => n5466);
   U251 : AOI21_X1 port map( B1 => IR_FAIL(0), B2 => n5467, A => PC_FAIL(0), ZN
                           => n5464);
   U252 : OAI33_X1 port map( A1 => n5516, A2 => add_59_n1, A3 => n5466, B1 => 
                           n5465, B2 => n5464, B3 => add_53_aco_n2, ZN => 
                           n60_port);
   U253 : NOR2_X1 port map( A1 => PC_IN(2), A2 => n5324, ZN => n62_port);
   U254 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(5), ZN => n7);
   U255 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(2), ZN => n8);
   U256 : AND2_X1 port map( A1 => n5467, A2 => IR_FAIL(3), ZN => n9);
   U257 : OAI211_X1 port map( C1 => n5491, C2 => PC_IN(22), A => n5490, B => 
                           RST, ZN => n5468);
   U258 : INV_X1 port map( A => n5468, ZN => n292);
   U259 : OAI211_X1 port map( C1 => n5494, C2 => PC_IN(20), A => n5493, B => 
                           RST, ZN => n5469);
   U260 : INV_X1 port map( A => n5469, ZN => n290);
   U261 : OAI211_X1 port map( C1 => n5500, C2 => PC_IN(16), A => n5499, B => 
                           RST, ZN => n5470);
   U262 : INV_X1 port map( A => n5470, ZN => n289);
   U263 : OAI211_X1 port map( C1 => n5485, C2 => PC_IN(26), A => n5484, B => 
                           RST, ZN => n5471);
   U264 : INV_X1 port map( A => n5471, ZN => n288);
   U265 : OAI211_X1 port map( C1 => n5488, C2 => PC_IN(24), A => n5487, B => 
                           RST, ZN => n5472);
   U266 : INV_X1 port map( A => n5472, ZN => n287);
   U267 : OAI211_X1 port map( C1 => n5509, C2 => PC_IN(10), A => n5508, B => 
                           RST, ZN => n5473);
   U268 : INV_X1 port map( A => n5473, ZN => n285);
   U269 : OAI211_X1 port map( C1 => n5506, C2 => PC_IN(12), A => n5505, B => 
                           RST, ZN => n5474);
   U270 : INV_X1 port map( A => n5474, ZN => n284);
   U271 : OAI211_X1 port map( C1 => n5497, C2 => PC_IN(18), A => n5496, B => 
                           RST, ZN => n5475);
   U272 : INV_X1 port map( A => n5475, ZN => n283);
   U273 : OAI211_X1 port map( C1 => n5482, C2 => PC_IN(28), A => n5481, B => 
                           RST, ZN => n5476);
   U274 : INV_X1 port map( A => n5476, ZN => n282);
   U275 : OAI211_X1 port map( C1 => n5503, C2 => PC_IN(14), A => n5502, B => 
                           RST, ZN => n5477);
   U276 : INV_X1 port map( A => n5477, ZN => n281);
   U277 : OAI211_X1 port map( C1 => n5512, C2 => PC_IN(8), A => n5511, B => RST
                           , ZN => n5478);
   U278 : INV_X1 port map( A => n5478, ZN => n280);
   U279 : AOI211_X1 port map( C1 => n5481, C2 => n5480, A => n5479, B => n5324,
                           ZN => n58_port);
   U280 : AOI211_X1 port map( C1 => n5484, C2 => n5483, A => n5482, B => n5324,
                           ZN => n57_port);
   U281 : AOI211_X1 port map( C1 => n5487, C2 => n5486, A => n5485, B => n5324,
                           ZN => n56_port);
   U282 : AOI211_X1 port map( C1 => n5490, C2 => n5489, A => n5488, B => n5324,
                           ZN => n55_port);
   U283 : AOI211_X1 port map( C1 => n5493, C2 => n5492, A => n5491, B => n5324,
                           ZN => n54_port);
   U284 : AOI211_X1 port map( C1 => n5496, C2 => n5495, A => n5494, B => n5325,
                           ZN => n53_port);
   U285 : AOI211_X1 port map( C1 => n5499, C2 => n5498, A => n5497, B => n5325,
                           ZN => n52_port);
   U286 : AOI211_X1 port map( C1 => n5502, C2 => n5501, A => n5500, B => n5325,
                           ZN => n51_port);
   U287 : AOI211_X1 port map( C1 => n5505, C2 => n5504, A => n5503, B => n5325,
                           ZN => n50_port);
   U288 : AOI211_X1 port map( C1 => n5508, C2 => n5507, A => n5506, B => n5325,
                           ZN => n49_port);
   U289 : AOI211_X1 port map( C1 => n5511, C2 => n5510, A => n5509, B => n5325,
                           ZN => n48_port);
   U290 : AOI211_X1 port map( C1 => n5514, C2 => n5513, A => n5512, B => n5324,
                           ZN => n47_port);
   U291 : AOI222_X1 port map( A1 => n5548, A2 => N47, B1 => n5320, B2 => N220, 
                           C1 => n5547, C2 => N82, ZN => n5517);
   U292 : INV_X1 port map( A => n5517, ZN => n46);
   U293 : AOI222_X1 port map( A1 => n5548, A2 => N48, B1 => n5320, B2 => N221, 
                           C1 => n5322, C2 => N83, ZN => n5518);
   U294 : INV_X1 port map( A => n5518, ZN => n45);
   U295 : AOI222_X1 port map( A1 => n5548, A2 => N49, B1 => n5320, B2 => N222, 
                           C1 => n5547, C2 => N84, ZN => n5519);
   U296 : INV_X1 port map( A => n5519, ZN => n44);
   U297 : AOI222_X1 port map( A1 => n5548, A2 => N50, B1 => n5320, B2 => N223, 
                           C1 => n5322, C2 => N85, ZN => n5520);
   U298 : INV_X1 port map( A => n5520, ZN => n43);
   U299 : AOI222_X1 port map( A1 => n5548, A2 => N51, B1 => n5320, B2 => N224, 
                           C1 => n5547, C2 => N86, ZN => n5521);
   U300 : INV_X1 port map( A => n5521, ZN => n42);
   U301 : AOI222_X1 port map( A1 => n5548, A2 => N52, B1 => n5320, B2 => N225, 
                           C1 => n5322, C2 => N87, ZN => n5522);
   U302 : INV_X1 port map( A => n5522, ZN => n41);
   U303 : AOI222_X1 port map( A1 => n5548, A2 => N53, B1 => n5320, B2 => N226, 
                           C1 => n5547, C2 => N88, ZN => n5523);
   U304 : INV_X1 port map( A => n5523, ZN => n40);
   U305 : AOI222_X1 port map( A1 => n5548, A2 => N54, B1 => n5320, B2 => N227, 
                           C1 => n5547, C2 => N89, ZN => n5524);
   U306 : INV_X1 port map( A => n5524, ZN => n39);
   U307 : AOI222_X1 port map( A1 => n5548, A2 => N55, B1 => n5320, B2 => N228, 
                           C1 => n5547, C2 => N90, ZN => n5525);
   U308 : INV_X1 port map( A => n5525, ZN => n38);
   U309 : AOI222_X1 port map( A1 => n5548, A2 => N56, B1 => n5320, B2 => N229, 
                           C1 => n5547, C2 => N91, ZN => n5526);
   U310 : INV_X1 port map( A => n5526, ZN => n37);
   U311 : AOI222_X1 port map( A1 => n5548, A2 => N57, B1 => n5320, B2 => N230, 
                           C1 => n5547, C2 => N92, ZN => n5527);
   U312 : INV_X1 port map( A => n5527, ZN => n36);
   U313 : AOI222_X1 port map( A1 => n5548, A2 => N58, B1 => n5320, B2 => N231, 
                           C1 => n5547, C2 => N93, ZN => n5528);
   U314 : INV_X1 port map( A => n5528, ZN => n35);
   U315 : AOI222_X1 port map( A1 => n5548, A2 => N59, B1 => n5320, B2 => N232, 
                           C1 => n5322, C2 => N94, ZN => n5529);
   U316 : INV_X1 port map( A => n5529, ZN => n34);
   U317 : AOI222_X1 port map( A1 => n5548, A2 => N60, B1 => n5320, B2 => N233, 
                           C1 => n5322, C2 => N95, ZN => n5530);
   U318 : INV_X1 port map( A => n5530, ZN => n33);
   U319 : AOI222_X1 port map( A1 => n5548, A2 => N61, B1 => n5320, B2 => N234, 
                           C1 => n5322, C2 => N96, ZN => n5531);
   U320 : INV_X1 port map( A => n5531, ZN => n32);
   U321 : AOI222_X1 port map( A1 => n5548, A2 => N62, B1 => n5320, B2 => N235, 
                           C1 => n5322, C2 => N97, ZN => n5532);
   U322 : INV_X1 port map( A => n5532, ZN => n31);
   U323 : AOI222_X1 port map( A1 => n5548, A2 => N63, B1 => n5320, B2 => N236, 
                           C1 => n5322, C2 => N98, ZN => n5533);
   U324 : INV_X1 port map( A => n5533, ZN => n30);
   U325 : AOI222_X1 port map( A1 => n5548, A2 => N64, B1 => n5320, B2 => N237, 
                           C1 => n5322, C2 => N99, ZN => n5534);
   U326 : INV_X1 port map( A => n5534, ZN => n29);
   U327 : AOI222_X1 port map( A1 => n5548, A2 => N65, B1 => n5320, B2 => N238, 
                           C1 => n5322, C2 => N100, ZN => n5535);
   U328 : INV_X1 port map( A => n5535, ZN => n28);
   U329 : AOI222_X1 port map( A1 => n5548, A2 => N66, B1 => n5320, B2 => N239, 
                           C1 => n5547, C2 => N101, ZN => n5536);
   U330 : INV_X1 port map( A => n5536, ZN => n27);
   U331 : AOI222_X1 port map( A1 => n5548, A2 => N67, B1 => n5320, B2 => N240, 
                           C1 => n5322, C2 => N102, ZN => n5537);
   U332 : INV_X1 port map( A => n5537, ZN => n26);
   U333 : AOI222_X1 port map( A1 => n5548, A2 => N68, B1 => n5320, B2 => N241, 
                           C1 => n5547, C2 => N103, ZN => n5538);
   U334 : INV_X1 port map( A => n5538, ZN => n25);
   U335 : AOI222_X1 port map( A1 => n5548, A2 => N69, B1 => n5320, B2 => N242, 
                           C1 => n5322, C2 => N104, ZN => n5539);
   U336 : INV_X1 port map( A => n5539, ZN => n24);
   U337 : AOI222_X1 port map( A1 => n5548, A2 => N70, B1 => n5320, B2 => N243, 
                           C1 => n5547, C2 => N105, ZN => n5540);
   U338 : INV_X1 port map( A => n5540, ZN => n23);
   U339 : AOI222_X1 port map( A1 => n5548, A2 => N71, B1 => n5320, B2 => N244, 
                           C1 => n5322, C2 => N106, ZN => n5541);
   U340 : INV_X1 port map( A => n5541, ZN => n22);
   U341 : AOI222_X1 port map( A1 => n5548, A2 => N72, B1 => n5320, B2 => N245, 
                           C1 => n5322, C2 => N107, ZN => n5542);
   U342 : INV_X1 port map( A => n5542, ZN => n21);
   U343 : AOI222_X1 port map( A1 => n5548, A2 => N73, B1 => n5320, B2 => N246, 
                           C1 => n5322, C2 => N108, ZN => n5543);
   U344 : INV_X1 port map( A => n5543, ZN => n20);
   U345 : AOI222_X1 port map( A1 => n5548, A2 => N74, B1 => n5320, B2 => N247, 
                           C1 => n5322, C2 => N109, ZN => n5544);
   U346 : INV_X1 port map( A => n5544, ZN => n4);
   U347 : AOI222_X1 port map( A1 => n5548, A2 => N75, B1 => n5320, B2 => N248, 
                           C1 => n5322, C2 => N110, ZN => n5545);
   U348 : INV_X1 port map( A => n5545, ZN => n3);
   U349 : AOI222_X1 port map( A1 => n5548, A2 => N76, B1 => n5320, B2 => N249, 
                           C1 => n5322, C2 => N111, ZN => n5546);
   U350 : INV_X1 port map( A => n5546, ZN => n2);
   U351 : AOI222_X1 port map( A1 => n5548, A2 => N77, B1 => n5320, B2 => N250, 
                           C1 => n5322, C2 => N112, ZN => n5549);
   U352 : INV_X1 port map( A => n5549, ZN => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity register_file_N32_addBit5 is

   port( RESET, RE, WE : in std_logic;  ADD_WR, ADD_RDA, ADD_RDB : in 
         std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUTA, OUTB : out std_logic_vector (31 downto 0));

end register_file_N32_addBit5;

architecture SYN_A of register_file_N32_addBit5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N243, N244, N245, N246, N247, 
      N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, 
      N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, n36859, 
      n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, 
      n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, 
      n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, 
      n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, 
      n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, 
      n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, 
      n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, 
      n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, 
      n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, 
      n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, 
      n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, 
      n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, 
      n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, 
      n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, 
      n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, 
      n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, 
      n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, 
      n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, 
      n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, 
      n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, 
      n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, 
      n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, 
      n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, 
      n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, 
      n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, 
      n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, 
      n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, 
      n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, 
      n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, 
      n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, 
      n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, 
      n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, 
      n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, 
      n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, 
      n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, 
      n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, 
      n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, 
      n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, 
      n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, 
      n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, 
      n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, 
      n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, 
      n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, 
      n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, 
      n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, 
      n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, 
      n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, 
      n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, 
      n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, 
      n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, 
      n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, 
      n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, 
      n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, 
      n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, 
      n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, 
      n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, 
      n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, 
      n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, 
      n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, 
      n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, 
      n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, 
      n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, 
      n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, 
      n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, 
      n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, 
      n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, 
      n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, 
      n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, 
      n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, 
      n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, 
      n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, 
      n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, 
      n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, 
      n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, 
      n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, 
      n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, 
      n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, 
      n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, 
      n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, 
      n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, 
      n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, 
      n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, 
      n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, 
      n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, 
      n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, 
      n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, 
      n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, 
      n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, 
      n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, 
      n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, 
      n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, 
      n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, 
      n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, 
      n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, 
      n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, 
      n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, 
      n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, 
      n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, 
      n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, 
      n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, 
      n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, 
      n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, 
      n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, 
      n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, 
      n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, 
      n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, 
      n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, 
      n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, 
      n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, 
      n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, 
      n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, 
      n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, 
      n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, 
      n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, 
      n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, 
      n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, 
      n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, 
      n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, 
      n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, 
      n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, 
      n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, 
      n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, 
      n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, 
      n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, 
      n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, 
      n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, 
      n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, 
      n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, 
      n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, 
      n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, 
      n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, 
      n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, 
      n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, 
      n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, 
      n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, 
      n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, 
      n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, 
      n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, 
      n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, 
      n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, 
      n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, 
      n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, 
      n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, 
      n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, 
      n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, 
      n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, 
      n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, 
      n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, 
      n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, 
      n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, 
      n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, 
      n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, 
      n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, 
      n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, 
      n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, 
      n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, 
      n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, 
      n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, 
      n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, 
      n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, 
      n38300, n38301, n38302, n38303, n38304, n38305 : std_logic;

begin
   
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => n37757, D => N275, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => n37757, D => N274, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => n37757, D => N273, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => N305, D => N272, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => n37757, D => N271, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N305, D => N270, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => n37757, D => N269, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => n37757, D => N268, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => n37757, D => N267, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => n37757, D => N266, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => N305, D => N265, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => n37757, D => N264, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => n37757, D => N263, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => N305, D => N262, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => N305, D => N261, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => n37757, D => N260, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N305, D => N259, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => N305, D => N258, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N305, D => N257, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N305, D => N256, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => n37757, D => N255, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => N305, D => N254, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => N305, D => N253, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => N305, D => N252, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => n37757, D => N251, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => n37757, D => N250, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => n37757, D => N249, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => N305, D => N248, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => N305, D => N247, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => N305, D => N246, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => n37757, D => N245, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => n37757, D => N244, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => n37758, D => N275, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => n37758, D => N274, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => n37758, D => N273, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => n37758, D => N272, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => n37758, D => N271, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => n37758, D => N270, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => N304, D => N269, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => N304, D => N268, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => n37758, D => N267, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => n37758, D => N266, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => n37758, D => N265, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => n37758, D => N264, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => n37758, D => N263, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => N304, D => N262, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => n37758, D => N261, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N304, D => N260, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => n37758, D => N259, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N304, D => N258, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N304, D => N257, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N304, D => N256, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => N304, D => N255, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => n37758, D => N254, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => N304, D => N253, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => N304, D => N252, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => n37758, D => N251, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => n37758, D => N250, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => N304, D => N249, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => N304, D => N248, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => N304, D => N247, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => N304, D => N246, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => n37758, D => N245, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => N304, D => N244, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => n37759, D => N275, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => n37759, D => N274, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => n37759, D => N273, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => n37759, D => N272, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => n37759, D => N271, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => n37759, D => N270, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => N303, D => N269, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => N303, D => N268, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => n37759, D => N267, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => n37759, D => N266, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => n37759, D => N265, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => n37759, D => N264, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => n37759, D => N263, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => N303, D => N262, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => n37759, D => N261, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N303, D => N260, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => n37759, D => N259, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N303, D => N258, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N303, D => N257, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N303, D => N256, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => N303, D => N255, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => n37759, D => N254, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => N303, D => N253, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => N303, D => N252, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => n37759, D => N251, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => n37759, D => N250, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => N303, D => N249, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => N303, D => N248, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => N303, D => N247, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => N303, D => N246, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => n37759, D => N245, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => N303, D => N244, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => n37760, D => N275, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => n37760, D => N274, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => n37760, D => N273, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => n37760, D => N272, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => n37760, D => N271, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => n37760, D => N270, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => N302, D => N269, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => N302, D => N268, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => n37760, D => N267, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => n37760, D => N266, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => n37760, D => N265, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => n37760, D => N264, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => n37760, D => N263, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => N302, D => N262, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => n37760, D => N261, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N302, D => N260, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => n37760, D => N259, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N302, D => N258, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N302, D => N257, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N302, D => N256, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => N302, D => N255, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => n37760, D => N254, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => N302, D => N253, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => N302, D => N252, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => N302, D => N251, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => n37760, D => N250, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => N302, D => N249, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => N302, D => N248, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => N302, D => N247, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => N302, D => N246, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => n37760, D => N245, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => n37760, D => N244, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => n37761, D => N275, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => n37761, D => N274, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => n37761, D => N273, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => n37761, D => N272, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => n37761, D => N271, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => n37761, D => N270, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => N301, D => N269, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => N301, D => N268, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => n37761, D => N267, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => n37761, D => N266, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => n37761, D => N265, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => n37761, D => N264, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => n37761, D => N263, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => N301, D => N262, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => n37761, D => N261, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N301, D => N260, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => n37761, D => N259, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N301, D => N258, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N301, D => N257, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N301, D => N256, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => N301, D => N255, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => n37761, D => N254, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => N301, D => N253, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => N301, D => N252, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => n37761, D => N251, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => n37761, D => N250, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => N301, D => N249, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => N301, D => N248, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => N301, D => N247, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => N301, D => N246, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => n37761, D => N245, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => N301, D => N244, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => n37762, D => N275, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => n37762, D => N274, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => n37762, D => N273, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => n37762, D => N272, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => n37762, D => N271, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => n37762, D => N270, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => N300, D => N269, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => N300, D => N268, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => n37762, D => N267, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => n37762, D => N266, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => n37762, D => N265, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => n37762, D => N264, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => n37762, D => N263, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => N300, D => N262, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => n37762, D => N261, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N300, D => N260, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => n37762, D => N259, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N300, D => N258, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N300, D => N257, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N300, D => N256, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => N300, D => N255, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => n37762, D => N254, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => N300, D => N253, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => N300, D => N252, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => N300, D => N251, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => n37762, D => N250, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => N300, D => N249, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => N300, D => N248, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => N300, D => N247, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => N300, D => N246, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => n37762, D => N245, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => n37762, D => N244, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => n37763, D => N275, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => n37763, D => N274, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => n37763, D => N273, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => n37763, D => N272, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => n37763, D => N271, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => n37763, D => N270, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => N299, D => N269, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => N299, D => N268, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => n37763, D => N267, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => n37763, D => N266, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => n37763, D => N265, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => n37763, D => N264, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => n37763, D => N263, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => N299, D => N262, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => n37763, D => N261, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N299, D => N260, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => n37763, D => N259, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N299, D => N258, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N299, D => N257, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N299, D => N256, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => N299, D => N255, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => n37763, D => N254, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => N299, D => N253, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => N299, D => N252, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => n37763, D => N251, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => n37763, D => N250, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => N299, D => N249, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => N299, D => N248, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => N299, D => N247, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => N299, D => N246, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => n37763, D => N245, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => N299, D => N244, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => n37764, D => N275, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => n37764, D => N274, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => n37764, D => N273, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => n37764, D => N272, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => n37764, D => N271, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => n37764, D => N270, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => N298, D => N269, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => N298, D => N268, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => n37764, D => N267, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => n37764, D => N266, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => n37764, D => N265, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => n37764, D => N264, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => n37764, D => N263, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => N298, D => N262, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => n37764, D => N261, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => N298, D => N260, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => n37764, D => N259, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N298, D => N258, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N298, D => N257, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N298, D => N256, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => N298, D => N255, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => n37764, D => N254, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => N298, D => N253, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => N298, D => N252, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => n37764, D => N251, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => n37764, D => N250, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => N298, D => N249, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => N298, D => N248, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => N298, D => N247, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => N298, D => N246, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => n37764, D => N245, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N298, D => N244, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => n37765, D => N275, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => n37765, D => N274, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => n37765, D => N273, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => n37765, D => N272, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => n37765, D => N271, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => n37765, D => N270, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => N297, D => N269, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => N297, D => N268, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => n37765, D => N267, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => n37765, D => N266, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => n37765, D => N265, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => n37765, D => N264, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => n37765, D => N263, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => N297, D => N262, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => n37765, D => N261, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N297, D => N260, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => n37765, D => N259, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N297, D => N258, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N297, D => N257, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N297, D => N256, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => N297, D => N255, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => n37765, D => N254, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => N297, D => N253, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => N297, D => N252, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => n37765, D => N251, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => n37765, D => N250, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => N297, D => N249, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => N297, D => N248, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => N297, D => N247, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => N297, D => N246, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => n37765, D => N245, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => N297, D => N244, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => n37766, D => N275, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => n37766, D => N274, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => n37766, D => N273, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => n37766, D => N272, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => n37766, D => N271, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => n37766, D => N270, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => N296, D => N269, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => N296, D => N268, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => n37766, D => N267, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => N296, D => N266, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => n37766, D => N265, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => n37766, D => N264, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => n37766, D => N263, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => N296, D => N262, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N296, D => N261, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => n37766, D => N260, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N296, D => N259, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => n37766, D => N258, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => n37766, D => N257, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N296, D => N256, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => n37766, D => N255, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => n37766, D => N254, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => N296, D => N253, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => N296, D => N252, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => N296, D => N251, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => n37766, D => N250, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => N296, D => N249, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => N296, D => N248, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => N296, D => N247, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => N296, D => N246, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => n37766, D => N245, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N296, D => N244, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => n37767, D => N275, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => n37767, D => N274, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => n37767, D => N273, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => n37767, D => N272, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => n37767, D => N271, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => n37767, D => N270, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => N295, D => N269, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => N295, D => N268, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => n37767, D => N267, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => n37767, D => N266, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => n37767, D => N265, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => n37767, D => N264, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => n37767, D => N263, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => N295, D => N262, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => n37767, D => N261, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N295, D => N260, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => n37767, D => N259, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N295, D => N258, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N295, D => N257, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N295, D => N256, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => N295, D => N255, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => n37767, D => N254, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => N295, D => N253, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => N295, D => N252, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => n37767, D => N251, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => n37767, D => N250, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => N295, D => N249, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => N295, D => N248, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => N295, D => N247, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => N295, D => N246, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => n37767, D => N245, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => N295, D => N244, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => n37768, D => N275, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => n37768, D => N274, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => n37768, D => N273, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => n37768, D => N272, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => n37768, D => N271, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => n37768, D => N270, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => N294, D => N269, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => N294, D => N268, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => n37768, D => N267, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => n37768, D => N266, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => n37768, D => N265, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => n37768, D => N264, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => n37768, D => N263, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => N294, D => N262, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => n37768, D => N261, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N294, D => N260, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => n37768, D => N259, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N294, D => N258, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N294, D => N257, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N294, D => N256, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => n37768, D => N255, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => n37768, D => N254, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => N294, D => N253, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => N294, D => N252, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => N294, D => N251, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => n37768, D => N250, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => N294, D => N249, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => N294, D => N248, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => N294, D => N247, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => N294, D => N246, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => n37768, D => N245, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => N294, D => N244, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => n37769, D => N275, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => n37769, D => N274, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => n37769, D => N273, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => n37769, D => N272, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => n37769, D => N271, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => n37769, D => N270, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => N293, D => N269, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => N293, D => N268, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => n37769, D => N267, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => n37769, D => N266, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => n37769, D => N265, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => n37769, D => N264, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => n37769, D => N263, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => N293, D => N262, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => n37769, D => N261, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N293, D => N260, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => n37769, D => N259, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N293, D => N258, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N293, D => N257, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N293, D => N256, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => N293, D => N255, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => n37769, D => N254, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => N293, D => N253, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => N293, D => N252, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => n37769, D => N251, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => n37769, D => N250, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => N293, D => N249, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => N293, D => N248, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => N293, D => N247, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => N293, D => N246, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => n37769, D => N245, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => N293, D => N244, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => n37770, D => N275, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => n37770, D => N274, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => n37770, D => N273, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => n37770, D => N272, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => n37770, D => N271, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => n37770, D => N270, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => N292, D => N269, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => N292, D => N268, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => n37770, D => N267, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => n37770, D => N266, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => n37770, D => N265, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => n37770, D => N264, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => n37770, D => N263, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => N292, D => N262, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => n37770, D => N261, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N292, D => N260, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => n37770, D => N259, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N292, D => N258, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N292, D => N257, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N292, D => N256, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => N292, D => N255, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => n37770, D => N254, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => N292, D => N253, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => N292, D => N252, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => n37770, D => N251, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => n37770, D => N250, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => N292, D => N249, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => N292, D => N248, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => N292, D => N247, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => N292, D => N246, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => n37770, D => N245, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => N292, D => N244, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => n37771, D => N275, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => n37771, D => N274, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => n37771, D => N273, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => n37771, D => N272, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => n37771, D => N271, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => n37771, D => N270, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => N291, D => N269, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => N291, D => N268, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => n37771, D => N267, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => n37771, D => N266, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => n37771, D => N265, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => n37771, D => N264, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => n37771, D => N263, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => N291, D => N262, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => n37771, D => N261, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N291, D => N260, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => n37771, D => N259, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N291, D => N258, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N291, D => N257, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N291, D => N256, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => N291, D => N255, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => n37771, D => N254, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => N291, D => N253, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => N291, D => N252, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => n37771, D => N251, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => n37771, D => N250, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => N291, D => N249, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => N291, D => N248, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => N291, D => N247, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => N291, D => N246, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => n37771, D => N245, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => N291, D => N244, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => n37772, D => N275, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => n37772, D => N274, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => n37772, D => N273, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => n37772, D => N272, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => n37772, D => N271, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => n37772, D => N270, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => N290, D => N269, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => N290, D => N268, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => n37772, D => N267, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => n37772, D => N266, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => n37772, D => N265, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => n37772, D => N264, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => n37772, D => N263, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => N290, D => N262, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => n37772, D => N261, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N290, D => N260, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => n37772, D => N259, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N290, D => N258, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N290, D => N257, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N290, D => N256, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => N290, D => N255, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => n37772, D => N254, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => N290, D => N253, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => N290, D => N252, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => n37772, D => N251, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => n37772, D => N250, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => N290, D => N249, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => N290, D => N248, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => N290, D => N247, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => N290, D => N246, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => n37772, D => N245, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => N290, D => N244, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => n37773, D => N275, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => n37773, D => N274, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => n37773, D => N273, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => n37773, D => N272, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => n37773, D => N271, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => n37773, D => N270, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => N289, D => N269, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => N289, D => N268, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => n37773, D => N267, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => n37773, D => N266, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => n37773, D => N265, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => n37773, D => N264, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => n37773, D => N263, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => N289, D => N262, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => n37773, D => N261, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N289, D => N260, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => n37773, D => N259, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N289, D => N258, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N289, D => N257, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N289, D => N256, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => N289, D => N255, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => n37773, D => N254, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => N289, D => N253, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => N289, D => N252, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => n37773, D => N251, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => n37773, D => N250, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => N289, D => N249, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => N289, D => N248, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => N289, D => N247, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => N289, D => N246, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => n37773, D => N245, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => N289, D => N244, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => n37774, D => N275, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => n37774, D => N274, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => n37774, D => N273, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => n37774, D => N272, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => n37774, D => N271, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => n37774, D => N270, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => N288, D => N269, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => N288, D => N268, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => n37774, D => N267, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => n37774, D => N266, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => n37774, D => N265, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => n37774, D => N264, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => n37774, D => N263, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => N288, D => N262, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => n37774, D => N261, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N288, D => N260, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => n37774, D => N259, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N288, D => N258, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N288, D => N257, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N288, D => N256, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => N288, D => N255, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => n37774, D => N254, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => N288, D => N253, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => N288, D => N252, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => n37774, D => N251, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => n37774, D => N250, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => N288, D => N249, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => N288, D => N248, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => N288, D => N247, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => N288, D => N246, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => n37774, D => N245, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => N288, D => N244, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => n37775, D => N275, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => n37775, D => N274, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => n37775, D => N273, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => n37775, D => N272, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => n37775, D => N271, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => n37775, D => N270, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => N287, D => N269, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => N287, D => N268, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => n37775, D => N267, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => n37775, D => N266, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => n37775, D => N265, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => n37775, D => N264, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => n37775, D => N263, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => N287, D => N262, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => n37775, D => N261, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N287, D => N260, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => n37775, D => N259, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N287, D => N258, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N287, D => N257, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N287, D => N256, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => N287, D => N255, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => n37775, D => N254, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => N287, D => N253, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => N287, D => N252, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => n37775, D => N251, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => n37775, D => N250, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => N287, D => N249, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => N287, D => N248, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => N287, D => N247, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => N287, D => N246, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => n37775, D => N245, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => N287, D => N244, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => n37776, D => N275, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => n37776, D => N274, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => n37776, D => N273, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => n37776, D => N272, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => n37776, D => N271, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => n37776, D => N270, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => N286, D => N269, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => N286, D => N268, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => n37776, D => N267, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => n37776, D => N266, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => n37776, D => N265, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => n37776, D => N264, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => n37776, D => N263, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => N286, D => N262, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => n37776, D => N261, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N286, D => N260, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => n37776, D => N259, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N286, D => N258, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N286, D => N257, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N286, D => N256, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => N286, D => N255, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => n37776, D => N254, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => N286, D => N253, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => N286, D => N252, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => n37776, D => N251, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => n37776, D => N250, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => N286, D => N249, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => N286, D => N248, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => N286, D => N247, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => N286, D => N246, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => n37776, D => N245, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => N286, D => N244, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => n37777, D => N275, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => n37777, D => N274, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => n37777, D => N273, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => n37777, D => N272, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => n37777, D => N271, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => n37777, D => N270, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => N285, D => N269, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => N285, D => N268, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => n37777, D => N267, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => n37777, D => N266, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => n37777, D => N265, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => n37777, D => N264, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => n37777, D => N263, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => N285, D => N262, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => n37777, D => N261, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N285, D => N260, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => n37777, D => N259, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N285, D => N258, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N285, D => N257, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N285, D => N256, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => N285, D => N255, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => n37777, D => N254, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => N285, D => N253, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => N285, D => N252, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => n37777, D => N251, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => n37777, D => N250, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => N285, D => N249, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => N285, D => N248, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => N285, D => N247, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => N285, D => N246, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => n37777, D => N245, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => N285, D => N244, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => n37778, D => N275, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => n37778, D => N274, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => n37778, D => N273, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => n37778, D => N272, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => n37778, D => N271, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => n37778, D => N270, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => N284, D => N269, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => N284, D => N268, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => n37778, D => N267, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => n37778, D => N266, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => n37778, D => N265, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => n37778, D => N264, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => n37778, D => N263, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => N284, D => N262, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => n37778, D => N261, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N284, D => N260, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => n37778, D => N259, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N284, D => N258, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N284, D => N257, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N284, D => N256, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => N284, D => N255, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => n37778, D => N254, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => N284, D => N253, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => N284, D => N252, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => n37778, D => N251, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => n37778, D => N250, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => N284, D => N249, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => N284, D => N248, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => N284, D => N247, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => N284, D => N246, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => n37778, D => N245, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => N284, D => N244, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => n37779, D => N275, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => n37779, D => N274, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => n37779, D => N273, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => n37779, D => N272, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => n37779, D => N271, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => n37779, D => N270, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => N283, D => N269, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => N283, D => N268, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => n37779, D => N267, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => n37779, D => N266, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => n37779, D => N265, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => n37779, D => N264, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => n37779, D => N263, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => N283, D => N262, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => n37779, D => N261, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N283, D => N260, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => n37779, D => N259, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N283, D => N258, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N283, D => N257, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N283, D => N256, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => N283, D => N255, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => n37779, D => N254, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => N283, D => N253, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => N283, D => N252, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => n37779, D => N251, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => n37779, D => N250, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => N283, D => N249, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => N283, D => N248, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => N283, D => N247, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => N283, D => N246, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => n37779, D => N245, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => N283, D => N244, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => n37780, D => N275, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => n37780, D => N274, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => n37780, D => N273, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => n37780, D => N272, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => n37780, D => N271, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => n37780, D => N270, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => n37780, D => N269, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => n37780, D => N268, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => n37780, D => N267, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => N282, D => N266, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => n37780, D => N265, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => n37780, D => N264, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => n37780, D => N263, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => N282, D => N262, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N282, D => N261, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N282, D => N260, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => n37780, D => N259, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N282, D => N258, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N282, D => N257, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => N282, D => N256, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => n37780, D => N255, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => n37780, D => N254, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => N282, D => N253, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => N282, D => N252, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => n37780, D => N251, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => n37780, D => N250, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => N282, D => N249, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => N282, D => N248, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => N282, D => N247, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => N282, D => N246, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => N282, D => N245, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => N282, D => N244, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => n37781, D => N275, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => n37781, D => N274, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => n37781, D => N273, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => n37781, D => N272, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => n37781, D => N271, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => n37781, D => N270, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => N281, D => N269, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => N281, D => N268, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => n37781, D => N267, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => n37781, D => N266, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => n37781, D => N265, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => n37781, D => N264, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => n37781, D => N263, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => N281, D => N262, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => n37781, D => N261, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N281, D => N260, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => n37781, D => N259, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N281, D => N258, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N281, D => N257, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N281, D => N256, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => N281, D => N255, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => n37781, D => N254, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => N281, D => N253, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => N281, D => N252, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => n37781, D => N251, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => n37781, D => N250, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => N281, D => N249, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => N281, D => N248, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => N281, D => N247, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => N281, D => N246, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => n37781, D => N245, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => N281, D => N244, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => n37782, D => N275, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => n37782, D => N274, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => n37782, D => N273, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => n37782, D => N272, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => n37782, D => N271, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => n37782, D => N270, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => N280, D => N269, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => N280, D => N268, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => n37782, D => N267, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => n37782, D => N266, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => n37782, D => N265, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => n37782, D => N264, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => n37782, D => N263, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => N280, D => N262, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => n37782, D => N261, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N280, D => N260, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => n37782, D => N259, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N280, D => N258, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N280, D => N257, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N280, D => N256, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => N280, D => N255, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => n37782, D => N254, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => N280, D => N253, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => N280, D => N252, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => n37782, D => N251, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => n37782, D => N250, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => N280, D => N249, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => N280, D => N248, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => N280, D => N247, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => N280, D => N246, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => n37782, D => N245, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => N280, D => N244, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => n37783, D => N275, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => n37783, D => N274, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => n37783, D => N273, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => n37783, D => N272, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => n37783, D => N271, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => n37783, D => N270, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => N279, D => N269, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => N279, D => N268, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => n37783, D => N267, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => n37783, D => N266, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => n37783, D => N265, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => n37783, D => N264, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => n37783, D => N263, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => N279, D => N262, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => n37783, D => N261, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N279, D => N260, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => n37783, D => N259, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N279, D => N258, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N279, D => N257, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N279, D => N256, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => N279, D => N255, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => n37783, D => N254, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => N279, D => N253, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => N279, D => N252, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => n37783, D => N251, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => n37783, D => N250, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => N279, D => N249, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => N279, D => N248, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => N279, D => N247, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => N279, D => N246, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => n37783, D => N245, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => N279, D => N244, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => n37784, D => N275, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => n37784, D => N274, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => n37784, D => N273, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => n37784, D => N272, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => n37784, D => N271, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => n37784, D => N270, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => N278, D => N269, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => N278, D => N268, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => n37784, D => N267, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => n37784, D => N266, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => n37784, D => N265, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => n37784, D => N264, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => n37784, D => N263, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => N278, D => N262, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => n37784, D => N261, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N278, D => N260, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => n37784, D => N259, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N278, D => N258, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N278, D => N257, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N278, D => N256, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => N278, D => N255, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => n37784, D => N254, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => N278, D => N253, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => N278, D => N252, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => n37784, D => N251, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => n37784, D => N250, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => N278, D => N249, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => N278, D => N248, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => N278, D => N247, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => N278, D => N246, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => n37784, D => N245, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => N278, D => N244, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => n37785, D => N275, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => n37785, D => N274, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => n37785, D => N273, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => n37785, D => N272, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => n37785, D => N271, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => n37785, D => N270, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => N277, D => N269, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => N277, D => N268, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => n37785, D => N267, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => n37785, D => N266, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => n37785, D => N265, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => n37785, D => N264, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => n37785, D => N263, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => N277, D => N262, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => n37785, D => N261, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N277, D => N260, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => n37785, D => N259, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N277, D => N258, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N277, D => N257, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N277, D => N256, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => N277, D => N255, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => n37785, D => N254, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => N277, D => N253, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => N277, D => N252, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => n37785, D => N251, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => n37785, D => N250, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => N277, D => N249, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => N277, D => N248, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => N277, D => N247, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => N277, D => N246, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => n37785, D => N245, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => N277, D => N244, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => n37786, D => N275, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => n37786, D => N274, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => n37786, D => N273, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => n37786, D => N272, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => n37786, D => N271, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => n37786, D => N270, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => N276, D => N269, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => N276, D => N268, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => n37786, D => N267, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => n37786, D => N266, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => n37786, D => N265, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => n37786, D => N264, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => n37786, D => N263, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => N276, D => N262, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => n37786, D => N261, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N276, D => N260, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => n37786, D => N259, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N276, D => N258, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N276, D => N257, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N276, D => N256, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => N276, D => N255, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => n37786, D => N254, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => N276, D => N253, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => N276, D => N252, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => n37786, D => N251, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => n37786, D => N250, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => N276, D => N249, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => N276, D => N248, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => N276, D => N247, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => N276, D => N246, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => n37786, D => N245, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => N276, D => N244, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => n37787, D => N275, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => n37787, D => N274, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => n37787, D => N273, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => n37787, D => N272, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => n37787, D => N271, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => n37787, D => N270, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => n37787, D => N269, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => n37787, D => N268, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => n37787, D => N267, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => n37787, D => N266, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => n37787, D => N265, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => N243, D => N264, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => n37787, D => N263, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => N243, D => N262, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => n37787, D => N261, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N243, D => N260, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => n37787, D => N259, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N243, D => N258, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N243, D => N257, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N243, D => N256, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => n37787, D => N255, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => n37787, D => N254, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => N243, D => N253, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => N243, D => N252, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => N243, D => N251, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => N243, D => N250, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => N243, D => N249, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => N243, D => N248, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => N243, D => N247, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => N243, D => N246, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => N243, D => N245, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => n37787, D => N244, Q => 
                           REGISTERS_31_0_port);
   U3 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n37741, B1 => 
                           REGISTERS_30_17_port, B2 => n37742, ZN => n36859);
   U4 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n37743, B1 => 
                           REGISTERS_27_17_port, B2 => n37744, ZN => n36860);
   U5 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n37745, B1 => 
                           REGISTERS_10_17_port, B2 => n37746, ZN => n36861);
   U6 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n37747, B1 => 
                           REGISTERS_6_17_port, B2 => n37748, ZN => n36862);
   U7 : NAND4_X1 port map( A1 => n36859, A2 => n36860, A3 => n36861, A4 => 
                           n36862, ZN => n36863);
   U8 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n37749, B1 => 
                           REGISTERS_26_17_port, B2 => n37750, ZN => n36864);
   U9 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n37751, B1 => 
                           REGISTERS_21_17_port, B2 => n37752, ZN => n36865);
   U10 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n37753, B1 => 
                           REGISTERS_23_17_port, B2 => n37754, ZN => n36866);
   U11 : AOI22_X1 port map( A1 => REGISTERS_19_17_port, A2 => n37755, B1 => 
                           REGISTERS_14_17_port, B2 => n37756, ZN => n36867);
   U12 : NAND4_X1 port map( A1 => n36864, A2 => n36865, A3 => n36866, A4 => 
                           n36867, ZN => n36868);
   U13 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n37726, B1 => 
                           REGISTERS_11_17_port, B2 => n37727, ZN => n36869);
   U14 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n37728, B1 => 
                           REGISTERS_1_17_port, B2 => n37729, ZN => n36870);
   U15 : AOI222_X1 port map( A1 => REGISTERS_15_17_port, A2 => n37730, B1 => 
                           REGISTERS_12_17_port, B2 => n37731, C1 => 
                           REGISTERS_13_17_port, C2 => n37732, ZN => n36871);
   U16 : NAND3_X1 port map( A1 => n36869, A2 => n36870, A3 => n36871, ZN => 
                           n36872);
   U17 : AOI22_X1 port map( A1 => REGISTERS_22_17_port, A2 => n37733, B1 => 
                           REGISTERS_20_17_port, B2 => n37734, ZN => n36873);
   U18 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n37735, B1 => 
                           REGISTERS_18_17_port, B2 => n37736, ZN => n36874);
   U19 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n37737, B1 => 
                           REGISTERS_2_17_port, B2 => n37738, ZN => n36875);
   U20 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n37739, B1 => 
                           REGISTERS_3_17_port, B2 => n37740, ZN => n36876);
   U21 : NAND4_X1 port map( A1 => n36873, A2 => n36874, A3 => n36875, A4 => 
                           n36876, ZN => n36877);
   U22 : OR4_X1 port map( A1 => n36863, A2 => n36868, A3 => n36872, A4 => 
                           n36877, ZN => OUTA(17));
   U23 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n37741, B1 => 
                           REGISTERS_30_16_port, B2 => n37742, ZN => n36878);
   U24 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n37743, B1 => 
                           REGISTERS_27_16_port, B2 => n37744, ZN => n36879);
   U25 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n37745, B1 => 
                           REGISTERS_10_16_port, B2 => n37746, ZN => n36880);
   U26 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n37747, B1 => 
                           REGISTERS_6_16_port, B2 => n37748, ZN => n36881);
   U27 : NAND4_X1 port map( A1 => n36878, A2 => n36879, A3 => n36880, A4 => 
                           n36881, ZN => n36882);
   U28 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n37749, B1 => 
                           REGISTERS_26_16_port, B2 => n37750, ZN => n36883);
   U29 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n37751, B1 => 
                           REGISTERS_21_16_port, B2 => n37752, ZN => n36884);
   U30 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n37753, B1 => 
                           REGISTERS_23_16_port, B2 => n37754, ZN => n36885);
   U31 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n37755, B1 => 
                           REGISTERS_14_16_port, B2 => n37756, ZN => n36886);
   U32 : NAND4_X1 port map( A1 => n36883, A2 => n36884, A3 => n36885, A4 => 
                           n36886, ZN => n36887);
   U33 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n37726, B1 => 
                           REGISTERS_11_16_port, B2 => n37727, ZN => n36888);
   U34 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n37728, B1 => 
                           REGISTERS_1_16_port, B2 => n37729, ZN => n36889);
   U35 : AOI222_X1 port map( A1 => REGISTERS_15_16_port, A2 => n37730, B1 => 
                           REGISTERS_12_16_port, B2 => n37731, C1 => 
                           REGISTERS_13_16_port, C2 => n37732, ZN => n36890);
   U36 : NAND3_X1 port map( A1 => n36888, A2 => n36889, A3 => n36890, ZN => 
                           n36891);
   U37 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n37733, B1 => 
                           REGISTERS_20_16_port, B2 => n37734, ZN => n36892);
   U38 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n37735, B1 => 
                           REGISTERS_18_16_port, B2 => n37736, ZN => n36893);
   U39 : AOI22_X1 port map( A1 => REGISTERS_31_16_port, A2 => n37737, B1 => 
                           REGISTERS_2_16_port, B2 => n37738, ZN => n36894);
   U40 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n37739, B1 => 
                           REGISTERS_3_16_port, B2 => n37740, ZN => n36895);
   U41 : NAND4_X1 port map( A1 => n36892, A2 => n36893, A3 => n36894, A4 => 
                           n36895, ZN => n36896);
   U42 : OR4_X1 port map( A1 => n36882, A2 => n36887, A3 => n36891, A4 => 
                           n36896, ZN => OUTA(16));
   U43 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n37741, B1 => 
                           REGISTERS_30_15_port, B2 => n37742, ZN => n36897);
   U44 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n37743, B1 => 
                           REGISTERS_27_15_port, B2 => n37744, ZN => n36898);
   U45 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n37745, B1 => 
                           REGISTERS_10_15_port, B2 => n37746, ZN => n36899);
   U46 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n37747, B1 => 
                           REGISTERS_6_15_port, B2 => n37748, ZN => n36900);
   U47 : NAND4_X1 port map( A1 => n36897, A2 => n36898, A3 => n36899, A4 => 
                           n36900, ZN => n36901);
   U48 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n37749, B1 => 
                           REGISTERS_26_15_port, B2 => n37750, ZN => n36902);
   U49 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n37751, B1 => 
                           REGISTERS_21_15_port, B2 => n37752, ZN => n36903);
   U50 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n37753, B1 => 
                           REGISTERS_23_15_port, B2 => n37754, ZN => n36904);
   U51 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n37755, B1 => 
                           REGISTERS_14_15_port, B2 => n37756, ZN => n36905);
   U52 : NAND4_X1 port map( A1 => n36902, A2 => n36903, A3 => n36904, A4 => 
                           n36905, ZN => n36906);
   U53 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n37726, B1 => 
                           REGISTERS_11_15_port, B2 => n37727, ZN => n36907);
   U54 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n37728, B1 => 
                           REGISTERS_1_15_port, B2 => n37729, ZN => n36908);
   U55 : AOI222_X1 port map( A1 => REGISTERS_15_15_port, A2 => n37730, B1 => 
                           REGISTERS_12_15_port, B2 => n37731, C1 => 
                           REGISTERS_13_15_port, C2 => n37732, ZN => n36909);
   U56 : NAND3_X1 port map( A1 => n36907, A2 => n36908, A3 => n36909, ZN => 
                           n36910);
   U57 : AOI22_X1 port map( A1 => REGISTERS_22_15_port, A2 => n37733, B1 => 
                           REGISTERS_20_15_port, B2 => n37734, ZN => n36911);
   U58 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n37735, B1 => 
                           REGISTERS_18_15_port, B2 => n37736, ZN => n36912);
   U59 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n37737, B1 => 
                           REGISTERS_2_15_port, B2 => n37738, ZN => n36913);
   U60 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n37739, B1 => 
                           REGISTERS_3_15_port, B2 => n37740, ZN => n36914);
   U61 : NAND4_X1 port map( A1 => n36911, A2 => n36912, A3 => n36913, A4 => 
                           n36914, ZN => n36915);
   U62 : OR4_X1 port map( A1 => n36901, A2 => n36906, A3 => n36910, A4 => 
                           n36915, ZN => OUTA(15));
   U63 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n37741, B1 => 
                           REGISTERS_30_14_port, B2 => n37742, ZN => n36916);
   U64 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n37743, B1 => 
                           REGISTERS_27_14_port, B2 => n37744, ZN => n36917);
   U65 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n37745, B1 => 
                           REGISTERS_10_14_port, B2 => n37746, ZN => n36918);
   U66 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n37747, B1 => 
                           REGISTERS_6_14_port, B2 => n37748, ZN => n36919);
   U67 : NAND4_X1 port map( A1 => n36916, A2 => n36917, A3 => n36918, A4 => 
                           n36919, ZN => n36920);
   U68 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n37749, B1 => 
                           REGISTERS_26_14_port, B2 => n37750, ZN => n36921);
   U69 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n37751, B1 => 
                           REGISTERS_21_14_port, B2 => n37752, ZN => n36922);
   U70 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n37753, B1 => 
                           REGISTERS_23_14_port, B2 => n37754, ZN => n36923);
   U71 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n37755, B1 => 
                           REGISTERS_14_14_port, B2 => n37756, ZN => n36924);
   U72 : NAND4_X1 port map( A1 => n36921, A2 => n36922, A3 => n36923, A4 => 
                           n36924, ZN => n36925);
   U73 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n37726, B1 => 
                           REGISTERS_11_14_port, B2 => n37727, ZN => n36926);
   U74 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n37728, B1 => 
                           REGISTERS_1_14_port, B2 => n37729, ZN => n36927);
   U75 : AOI222_X1 port map( A1 => REGISTERS_15_14_port, A2 => n37730, B1 => 
                           REGISTERS_12_14_port, B2 => n37731, C1 => 
                           REGISTERS_13_14_port, C2 => n37732, ZN => n36928);
   U76 : NAND3_X1 port map( A1 => n36926, A2 => n36927, A3 => n36928, ZN => 
                           n36929);
   U77 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n37733, B1 => 
                           REGISTERS_20_14_port, B2 => n37734, ZN => n36930);
   U78 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n37735, B1 => 
                           REGISTERS_18_14_port, B2 => n37736, ZN => n36931);
   U79 : AOI22_X1 port map( A1 => REGISTERS_31_14_port, A2 => n37737, B1 => 
                           REGISTERS_2_14_port, B2 => n37738, ZN => n36932);
   U80 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n37739, B1 => 
                           REGISTERS_3_14_port, B2 => n37740, ZN => n36933);
   U81 : NAND4_X1 port map( A1 => n36930, A2 => n36931, A3 => n36932, A4 => 
                           n36933, ZN => n36934);
   U82 : OR4_X1 port map( A1 => n36920, A2 => n36925, A3 => n36929, A4 => 
                           n36934, ZN => OUTA(14));
   U83 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n37741, B1 => 
                           REGISTERS_30_13_port, B2 => n37742, ZN => n36935);
   U84 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n37743, B1 => 
                           REGISTERS_27_13_port, B2 => n37744, ZN => n36936);
   U85 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n37745, B1 => 
                           REGISTERS_10_13_port, B2 => n37746, ZN => n36937);
   U86 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n37747, B1 => 
                           REGISTERS_6_13_port, B2 => n37748, ZN => n36938);
   U87 : NAND4_X1 port map( A1 => n36935, A2 => n36936, A3 => n36937, A4 => 
                           n36938, ZN => n36939);
   U88 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n37749, B1 => 
                           REGISTERS_26_13_port, B2 => n37750, ZN => n36940);
   U89 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n37751, B1 => 
                           REGISTERS_21_13_port, B2 => n37752, ZN => n36941);
   U90 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n37753, B1 => 
                           REGISTERS_23_13_port, B2 => n37754, ZN => n36942);
   U91 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n37755, B1 => 
                           REGISTERS_14_13_port, B2 => n37756, ZN => n36943);
   U92 : NAND4_X1 port map( A1 => n36940, A2 => n36941, A3 => n36942, A4 => 
                           n36943, ZN => n36944);
   U93 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n37726, B1 => 
                           REGISTERS_11_13_port, B2 => n37727, ZN => n36945);
   U94 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n37728, B1 => 
                           REGISTERS_1_13_port, B2 => n37729, ZN => n36946);
   U95 : AOI222_X1 port map( A1 => REGISTERS_15_13_port, A2 => n37730, B1 => 
                           REGISTERS_12_13_port, B2 => n37731, C1 => 
                           REGISTERS_13_13_port, C2 => n37732, ZN => n36947);
   U96 : NAND3_X1 port map( A1 => n36945, A2 => n36946, A3 => n36947, ZN => 
                           n36948);
   U97 : AOI22_X1 port map( A1 => REGISTERS_22_13_port, A2 => n37733, B1 => 
                           REGISTERS_20_13_port, B2 => n37734, ZN => n36949);
   U98 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n37735, B1 => 
                           REGISTERS_18_13_port, B2 => n37736, ZN => n36950);
   U99 : AOI22_X1 port map( A1 => REGISTERS_31_13_port, A2 => n37737, B1 => 
                           REGISTERS_2_13_port, B2 => n37738, ZN => n36951);
   U100 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n37739, B1 => 
                           REGISTERS_3_13_port, B2 => n37740, ZN => n36952);
   U101 : NAND4_X1 port map( A1 => n36949, A2 => n36950, A3 => n36951, A4 => 
                           n36952, ZN => n36953);
   U102 : OR4_X1 port map( A1 => n36939, A2 => n36944, A3 => n36948, A4 => 
                           n36953, ZN => OUTA(13));
   U103 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n37741, B1 => 
                           REGISTERS_30_12_port, B2 => n37742, ZN => n36954);
   U104 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n37743, B1 => 
                           REGISTERS_27_12_port, B2 => n37744, ZN => n36955);
   U105 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n37745, B1 => 
                           REGISTERS_10_12_port, B2 => n37746, ZN => n36956);
   U106 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n37747, B1 => 
                           REGISTERS_6_12_port, B2 => n37748, ZN => n36957);
   U107 : NAND4_X1 port map( A1 => n36954, A2 => n36955, A3 => n36956, A4 => 
                           n36957, ZN => n36958);
   U108 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n37749, B1 => 
                           REGISTERS_26_12_port, B2 => n37750, ZN => n36959);
   U109 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n37751, B1 => 
                           REGISTERS_21_12_port, B2 => n37752, ZN => n36960);
   U110 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n37753, B1 => 
                           REGISTERS_23_12_port, B2 => n37754, ZN => n36961);
   U111 : AOI22_X1 port map( A1 => REGISTERS_19_12_port, A2 => n37755, B1 => 
                           REGISTERS_14_12_port, B2 => n37756, ZN => n36962);
   U112 : NAND4_X1 port map( A1 => n36959, A2 => n36960, A3 => n36961, A4 => 
                           n36962, ZN => n36963);
   U113 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n37726, B1 => 
                           REGISTERS_11_12_port, B2 => n37727, ZN => n36964);
   U114 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n37728, B1 => 
                           REGISTERS_1_12_port, B2 => n37729, ZN => n36965);
   U115 : AOI222_X1 port map( A1 => REGISTERS_15_12_port, A2 => n37730, B1 => 
                           REGISTERS_12_12_port, B2 => n37731, C1 => 
                           REGISTERS_13_12_port, C2 => n37732, ZN => n36966);
   U116 : NAND3_X1 port map( A1 => n36964, A2 => n36965, A3 => n36966, ZN => 
                           n36967);
   U117 : AOI22_X1 port map( A1 => REGISTERS_22_12_port, A2 => n37733, B1 => 
                           REGISTERS_20_12_port, B2 => n37734, ZN => n36968);
   U118 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n37735, B1 => 
                           REGISTERS_18_12_port, B2 => n37736, ZN => n36969);
   U119 : AOI22_X1 port map( A1 => REGISTERS_31_12_port, A2 => n37737, B1 => 
                           REGISTERS_2_12_port, B2 => n37738, ZN => n36970);
   U120 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n37739, B1 => 
                           REGISTERS_3_12_port, B2 => n37740, ZN => n36971);
   U121 : NAND4_X1 port map( A1 => n36968, A2 => n36969, A3 => n36970, A4 => 
                           n36971, ZN => n36972);
   U122 : OR4_X1 port map( A1 => n36958, A2 => n36963, A3 => n36967, A4 => 
                           n36972, ZN => OUTA(12));
   U123 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n37741, B1 => 
                           REGISTERS_30_11_port, B2 => n37742, ZN => n36973);
   U124 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n37743, B1 => 
                           REGISTERS_27_11_port, B2 => n37744, ZN => n36974);
   U125 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n37745, B1 => 
                           REGISTERS_10_11_port, B2 => n37746, ZN => n36975);
   U126 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n37747, B1 => 
                           REGISTERS_6_11_port, B2 => n37748, ZN => n36976);
   U127 : NAND4_X1 port map( A1 => n36973, A2 => n36974, A3 => n36975, A4 => 
                           n36976, ZN => n36977);
   U128 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n37749, B1 => 
                           REGISTERS_26_11_port, B2 => n37750, ZN => n36978);
   U129 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n37751, B1 => 
                           REGISTERS_21_11_port, B2 => n37752, ZN => n36979);
   U130 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n37753, B1 => 
                           REGISTERS_23_11_port, B2 => n37754, ZN => n36980);
   U131 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n37755, B1 => 
                           REGISTERS_14_11_port, B2 => n37756, ZN => n36981);
   U132 : NAND4_X1 port map( A1 => n36978, A2 => n36979, A3 => n36980, A4 => 
                           n36981, ZN => n36982);
   U133 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n37726, B1 => 
                           REGISTERS_11_11_port, B2 => n37727, ZN => n36983);
   U134 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n37728, B1 => 
                           REGISTERS_1_11_port, B2 => n37729, ZN => n36984);
   U135 : AOI222_X1 port map( A1 => REGISTERS_15_11_port, A2 => n37730, B1 => 
                           REGISTERS_12_11_port, B2 => n37731, C1 => 
                           REGISTERS_13_11_port, C2 => n37732, ZN => n36985);
   U136 : NAND3_X1 port map( A1 => n36983, A2 => n36984, A3 => n36985, ZN => 
                           n36986);
   U137 : AOI22_X1 port map( A1 => REGISTERS_22_11_port, A2 => n37733, B1 => 
                           REGISTERS_20_11_port, B2 => n37734, ZN => n36987);
   U138 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n37735, B1 => 
                           REGISTERS_18_11_port, B2 => n37736, ZN => n36988);
   U139 : AOI22_X1 port map( A1 => REGISTERS_31_11_port, A2 => n37737, B1 => 
                           REGISTERS_2_11_port, B2 => n37738, ZN => n36989);
   U140 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n37739, B1 => 
                           REGISTERS_3_11_port, B2 => n37740, ZN => n36990);
   U141 : NAND4_X1 port map( A1 => n36987, A2 => n36988, A3 => n36989, A4 => 
                           n36990, ZN => n36991);
   U142 : OR4_X1 port map( A1 => n36977, A2 => n36982, A3 => n36986, A4 => 
                           n36991, ZN => OUTA(11));
   U143 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n37741, B1 => 
                           REGISTERS_30_10_port, B2 => n37742, ZN => n36992);
   U144 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n37743, B1 => 
                           REGISTERS_27_10_port, B2 => n37744, ZN => n36993);
   U145 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n37745, B1 => 
                           REGISTERS_10_10_port, B2 => n37746, ZN => n36994);
   U146 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n37747, B1 => 
                           REGISTERS_6_10_port, B2 => n37748, ZN => n36995);
   U147 : NAND4_X1 port map( A1 => n36992, A2 => n36993, A3 => n36994, A4 => 
                           n36995, ZN => n36996);
   U148 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n37749, B1 => 
                           REGISTERS_26_10_port, B2 => n37750, ZN => n36997);
   U149 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n37751, B1 => 
                           REGISTERS_21_10_port, B2 => n37752, ZN => n36998);
   U150 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n37753, B1 => 
                           REGISTERS_23_10_port, B2 => n37754, ZN => n36999);
   U151 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n37755, B1 => 
                           REGISTERS_14_10_port, B2 => n37756, ZN => n37000);
   U152 : NAND4_X1 port map( A1 => n36997, A2 => n36998, A3 => n36999, A4 => 
                           n37000, ZN => n37001);
   U153 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n37726, B1 => 
                           REGISTERS_11_10_port, B2 => n37727, ZN => n37002);
   U154 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n37728, B1 => 
                           REGISTERS_1_10_port, B2 => n37729, ZN => n37003);
   U155 : AOI222_X1 port map( A1 => REGISTERS_15_10_port, A2 => n37730, B1 => 
                           REGISTERS_12_10_port, B2 => n37731, C1 => 
                           REGISTERS_13_10_port, C2 => n37732, ZN => n37004);
   U156 : NAND3_X1 port map( A1 => n37002, A2 => n37003, A3 => n37004, ZN => 
                           n37005);
   U157 : AOI22_X1 port map( A1 => REGISTERS_22_10_port, A2 => n37733, B1 => 
                           REGISTERS_20_10_port, B2 => n37734, ZN => n37006);
   U158 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n37735, B1 => 
                           REGISTERS_18_10_port, B2 => n37736, ZN => n37007);
   U159 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n37737, B1 => 
                           REGISTERS_2_10_port, B2 => n37738, ZN => n37008);
   U160 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n37739, B1 => 
                           REGISTERS_3_10_port, B2 => n37740, ZN => n37009);
   U161 : NAND4_X1 port map( A1 => n37006, A2 => n37007, A3 => n37008, A4 => 
                           n37009, ZN => n37010);
   U162 : OR4_X1 port map( A1 => n36996, A2 => n37001, A3 => n37005, A4 => 
                           n37010, ZN => OUTA(10));
   U163 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_7_port, B1 => 
                           n37701, B2 => REGISTERS_16_7_port, ZN => n37011);
   U164 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_7_port, B1 => 
                           n37710, B2 => REGISTERS_6_7_port, ZN => n37012);
   U165 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_7_port, B1 => 
                           n37707, B2 => REGISTERS_24_7_port, ZN => n37013);
   U166 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_7_port, B1 => 
                           n37705, B2 => REGISTERS_12_7_port, ZN => n37014);
   U167 : NAND4_X1 port map( A1 => n37011, A2 => n37012, A3 => n37013, A4 => 
                           n37014, ZN => n37015);
   U168 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_7_port, B1 => 
                           n37703, B2 => REGISTERS_1_7_port, ZN => n37016);
   U169 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_7_port, B1 => 
                           n37699, B2 => REGISTERS_20_7_port, ZN => n37017);
   U170 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_7_port, B1 => 
                           n37700, B2 => REGISTERS_18_7_port, ZN => n37018);
   U171 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_7_port, B1 => 
                           n37718, B2 => REGISTERS_28_7_port, ZN => n37019);
   U172 : NAND4_X1 port map( A1 => n37016, A2 => n37017, A3 => n37018, A4 => 
                           n37019, ZN => n37020);
   U173 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_7_port, B1 => 
                           n37720, B2 => REGISTERS_11_7_port, ZN => n37021);
   U174 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_7_port, B1 => 
                           n38278, B2 => REGISTERS_2_7_port, ZN => n37022);
   U175 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_7_port, B1 => 
                           n37697, B2 => REGISTERS_13_7_port, C1 => n37722, C2 
                           => REGISTERS_19_7_port, ZN => n37023);
   U176 : NAND3_X1 port map( A1 => n37021, A2 => n37022, A3 => n37023, ZN => 
                           n37024);
   U177 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_7_port, B1 => 
                           n37715, B2 => REGISTERS_8_7_port, ZN => n37025);
   U178 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_7_port, B1 => 
                           n37711, B2 => REGISTERS_3_7_port, ZN => n37026);
   U179 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_7_port, B1 => 
                           n37717, B2 => REGISTERS_4_7_port, ZN => n37027);
   U180 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_7_port, B1 => 
                           n37724, B2 => REGISTERS_15_7_port, ZN => n37028);
   U181 : NAND4_X1 port map( A1 => n37025, A2 => n37026, A3 => n37027, A4 => 
                           n37028, ZN => n37029);
   U182 : OR4_X1 port map( A1 => n37015, A2 => n37020, A3 => n37024, A4 => 
                           n37029, ZN => OUTB(7));
   U183 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n37741, B1 => 
                           REGISTERS_30_7_port, B2 => n37742, ZN => n37030);
   U184 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n37743, B1 => 
                           REGISTERS_27_7_port, B2 => n37744, ZN => n37031);
   U185 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n37745, B1 => 
                           REGISTERS_10_7_port, B2 => n37746, ZN => n37032);
   U186 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n37747, B1 => 
                           REGISTERS_6_7_port, B2 => n37748, ZN => n37033);
   U187 : NAND4_X1 port map( A1 => n37030, A2 => n37031, A3 => n37032, A4 => 
                           n37033, ZN => n37034);
   U188 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n37749, B1 => 
                           REGISTERS_26_7_port, B2 => n37750, ZN => n37035);
   U189 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n37751, B1 => 
                           REGISTERS_21_7_port, B2 => n37752, ZN => n37036);
   U190 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n37753, B1 => 
                           REGISTERS_23_7_port, B2 => n37754, ZN => n37037);
   U191 : AOI22_X1 port map( A1 => REGISTERS_19_7_port, A2 => n37755, B1 => 
                           REGISTERS_14_7_port, B2 => n37756, ZN => n37038);
   U192 : NAND4_X1 port map( A1 => n37035, A2 => n37036, A3 => n37037, A4 => 
                           n37038, ZN => n37039);
   U193 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n37726, B1 => 
                           REGISTERS_11_7_port, B2 => n37727, ZN => n37040);
   U194 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n37728, B1 => 
                           REGISTERS_1_7_port, B2 => n37729, ZN => n37041);
   U195 : AOI222_X1 port map( A1 => REGISTERS_15_7_port, A2 => n37730, B1 => 
                           REGISTERS_12_7_port, B2 => n37731, C1 => 
                           REGISTERS_13_7_port, C2 => n38211, ZN => n37042);
   U196 : NAND3_X1 port map( A1 => n37040, A2 => n37041, A3 => n37042, ZN => 
                           n37043);
   U197 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n37733, B1 => 
                           REGISTERS_20_7_port, B2 => n37734, ZN => n37044);
   U198 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n37735, B1 => 
                           REGISTERS_18_7_port, B2 => n37736, ZN => n37045);
   U199 : AOI22_X1 port map( A1 => REGISTERS_31_7_port, A2 => n37737, B1 => 
                           REGISTERS_2_7_port, B2 => n37738, ZN => n37046);
   U200 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n37739, B1 => 
                           REGISTERS_3_7_port, B2 => n37740, ZN => n37047);
   U201 : NAND4_X1 port map( A1 => n37044, A2 => n37045, A3 => n37046, A4 => 
                           n37047, ZN => n37048);
   U202 : OR4_X1 port map( A1 => n37034, A2 => n37039, A3 => n37043, A4 => 
                           n37048, ZN => OUTA(7));
   U203 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_6_port, B1 => 
                           n37701, B2 => REGISTERS_16_6_port, ZN => n37049);
   U204 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_6_port, B1 => 
                           n37710, B2 => REGISTERS_6_6_port, ZN => n37050);
   U205 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_6_port, B1 => 
                           n37707, B2 => REGISTERS_24_6_port, ZN => n37051);
   U206 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_6_port, B1 => 
                           n37705, B2 => REGISTERS_12_6_port, ZN => n37052);
   U207 : NAND4_X1 port map( A1 => n37049, A2 => n37050, A3 => n37051, A4 => 
                           n37052, ZN => n37053);
   U208 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_6_port, B1 => 
                           n37703, B2 => REGISTERS_1_6_port, ZN => n37054);
   U209 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_6_port, B1 => 
                           n37699, B2 => REGISTERS_20_6_port, ZN => n37055);
   U210 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_6_port, B1 => 
                           n37700, B2 => REGISTERS_18_6_port, ZN => n37056);
   U211 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_6_port, B1 => 
                           n37718, B2 => REGISTERS_28_6_port, ZN => n37057);
   U212 : NAND4_X1 port map( A1 => n37054, A2 => n37055, A3 => n37056, A4 => 
                           n37057, ZN => n37058);
   U213 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_6_port, B1 => 
                           n37720, B2 => REGISTERS_11_6_port, ZN => n37059);
   U214 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_6_port, B1 => 
                           n38278, B2 => REGISTERS_2_6_port, ZN => n37060);
   U215 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_6_port, B1 => 
                           n37697, B2 => REGISTERS_13_6_port, C1 => n37722, C2 
                           => REGISTERS_19_6_port, ZN => n37061);
   U216 : NAND3_X1 port map( A1 => n37059, A2 => n37060, A3 => n37061, ZN => 
                           n37062);
   U217 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_6_port, B1 => 
                           n37715, B2 => REGISTERS_8_6_port, ZN => n37063);
   U218 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_6_port, B1 => 
                           n37711, B2 => REGISTERS_3_6_port, ZN => n37064);
   U219 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_6_port, B1 => 
                           n37717, B2 => REGISTERS_4_6_port, ZN => n37065);
   U220 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_6_port, B1 => 
                           n37724, B2 => REGISTERS_15_6_port, ZN => n37066);
   U221 : NAND4_X1 port map( A1 => n37063, A2 => n37064, A3 => n37065, A4 => 
                           n37066, ZN => n37067);
   U222 : OR4_X1 port map( A1 => n37053, A2 => n37058, A3 => n37062, A4 => 
                           n37067, ZN => OUTB(6));
   U223 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n37741, B1 => 
                           REGISTERS_30_1_port, B2 => n37742, ZN => n37068);
   U224 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n37743, B1 => 
                           REGISTERS_27_1_port, B2 => n37744, ZN => n37069);
   U225 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n37745, B1 => 
                           REGISTERS_10_1_port, B2 => n37746, ZN => n37070);
   U226 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n37747, B1 => 
                           REGISTERS_6_1_port, B2 => n37748, ZN => n37071);
   U227 : NAND4_X1 port map( A1 => n37068, A2 => n37069, A3 => n37070, A4 => 
                           n37071, ZN => n37072);
   U228 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n37749, B1 => 
                           REGISTERS_26_1_port, B2 => n37750, ZN => n37073);
   U229 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n37751, B1 => 
                           REGISTERS_21_1_port, B2 => n37752, ZN => n37074);
   U230 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n37753, B1 => 
                           REGISTERS_23_1_port, B2 => n37754, ZN => n37075);
   U231 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n37755, B1 => 
                           REGISTERS_14_1_port, B2 => n37756, ZN => n37076);
   U232 : NAND4_X1 port map( A1 => n37073, A2 => n37074, A3 => n37075, A4 => 
                           n37076, ZN => n37077);
   U233 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n37726, B1 => 
                           REGISTERS_11_1_port, B2 => n37727, ZN => n37078);
   U234 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n37728, B1 => 
                           REGISTERS_1_1_port, B2 => n37729, ZN => n37079);
   U235 : AOI222_X1 port map( A1 => REGISTERS_15_1_port, A2 => n37730, B1 => 
                           REGISTERS_12_1_port, B2 => n37731, C1 => 
                           REGISTERS_13_1_port, C2 => n37732, ZN => n37080);
   U236 : NAND3_X1 port map( A1 => n37078, A2 => n37079, A3 => n37080, ZN => 
                           n37081);
   U237 : AOI22_X1 port map( A1 => REGISTERS_22_1_port, A2 => n37733, B1 => 
                           REGISTERS_20_1_port, B2 => n37734, ZN => n37082);
   U238 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n37735, B1 => 
                           REGISTERS_18_1_port, B2 => n37736, ZN => n37083);
   U239 : AOI22_X1 port map( A1 => REGISTERS_31_1_port, A2 => n37737, B1 => 
                           REGISTERS_2_1_port, B2 => n37738, ZN => n37084);
   U240 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n37739, B1 => 
                           REGISTERS_3_1_port, B2 => n37740, ZN => n37085);
   U241 : NAND4_X1 port map( A1 => n37082, A2 => n37083, A3 => n37084, A4 => 
                           n37085, ZN => n37086);
   U242 : OR4_X1 port map( A1 => n37072, A2 => n37077, A3 => n37081, A4 => 
                           n37086, ZN => OUTA(1));
   U243 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_5_port, B1 => 
                           n37701, B2 => REGISTERS_16_5_port, ZN => n37087);
   U244 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_5_port, B1 => 
                           n37710, B2 => REGISTERS_6_5_port, ZN => n37088);
   U245 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_5_port, B1 => 
                           n37707, B2 => REGISTERS_24_5_port, ZN => n37089);
   U246 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_5_port, B1 => 
                           n37705, B2 => REGISTERS_12_5_port, ZN => n37090);
   U247 : NAND4_X1 port map( A1 => n37087, A2 => n37088, A3 => n37089, A4 => 
                           n37090, ZN => n37091);
   U248 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_5_port, B1 => 
                           n37703, B2 => REGISTERS_1_5_port, ZN => n37092);
   U249 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_5_port, B1 => 
                           n37699, B2 => REGISTERS_20_5_port, ZN => n37093);
   U250 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_5_port, B1 => 
                           n37700, B2 => REGISTERS_18_5_port, ZN => n37094);
   U251 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_5_port, B1 => 
                           n37718, B2 => REGISTERS_28_5_port, ZN => n37095);
   U252 : NAND4_X1 port map( A1 => n37092, A2 => n37093, A3 => n37094, A4 => 
                           n37095, ZN => n37096);
   U253 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_5_port, B1 => 
                           n37720, B2 => REGISTERS_11_5_port, ZN => n37097);
   U254 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_5_port, B1 => 
                           n38278, B2 => REGISTERS_2_5_port, ZN => n37098);
   U255 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_5_port, B1 => 
                           n37697, B2 => REGISTERS_13_5_port, C1 => n37722, C2 
                           => REGISTERS_19_5_port, ZN => n37099);
   U256 : NAND3_X1 port map( A1 => n37097, A2 => n37098, A3 => n37099, ZN => 
                           n37100);
   U257 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_5_port, B1 => 
                           n37715, B2 => REGISTERS_8_5_port, ZN => n37101);
   U258 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_5_port, B1 => 
                           n37711, B2 => REGISTERS_3_5_port, ZN => n37102);
   U259 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_5_port, B1 => 
                           n37717, B2 => REGISTERS_4_5_port, ZN => n37103);
   U260 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_5_port, B1 => 
                           n37724, B2 => REGISTERS_15_5_port, ZN => n37104);
   U261 : NAND4_X1 port map( A1 => n37101, A2 => n37102, A3 => n37103, A4 => 
                           n37104, ZN => n37105);
   U262 : OR4_X1 port map( A1 => n37091, A2 => n37096, A3 => n37100, A4 => 
                           n37105, ZN => OUTB(5));
   U263 : AOI22_X1 port map( A1 => n37741, A2 => REGISTERS_29_0_port, B1 => 
                           n37742, B2 => REGISTERS_30_0_port, ZN => n37106);
   U264 : AOI22_X1 port map( A1 => n37743, A2 => REGISTERS_4_0_port, B1 => 
                           n37744, B2 => REGISTERS_27_0_port, ZN => n37107);
   U265 : AOI22_X1 port map( A1 => n37745, A2 => REGISTERS_28_0_port, B1 => 
                           n37746, B2 => REGISTERS_10_0_port, ZN => n37108);
   U266 : AOI22_X1 port map( A1 => n37747, A2 => REGISTERS_7_0_port, B1 => 
                           n37748, B2 => REGISTERS_6_0_port, ZN => n37109);
   U267 : NAND4_X1 port map( A1 => n37106, A2 => n37107, A3 => n37108, A4 => 
                           n37109, ZN => n37110);
   U268 : AOI22_X1 port map( A1 => n37749, A2 => REGISTERS_5_0_port, B1 => 
                           n37750, B2 => REGISTERS_26_0_port, ZN => n37111);
   U269 : AOI22_X1 port map( A1 => n37751, A2 => REGISTERS_25_0_port, B1 => 
                           n37752, B2 => REGISTERS_21_0_port, ZN => n37112);
   U270 : AOI22_X1 port map( A1 => n37753, A2 => REGISTERS_17_0_port, B1 => 
                           n37754, B2 => REGISTERS_23_0_port, ZN => n37113);
   U271 : AOI22_X1 port map( A1 => n37755, A2 => REGISTERS_19_0_port, B1 => 
                           n37756, B2 => REGISTERS_14_0_port, ZN => n37114);
   U272 : NAND4_X1 port map( A1 => n37111, A2 => n37112, A3 => n37113, A4 => 
                           n37114, ZN => n37115);
   U273 : AOI22_X1 port map( A1 => n37726, A2 => REGISTERS_16_0_port, B1 => 
                           n37727, B2 => REGISTERS_11_0_port, ZN => n37116);
   U274 : AOI22_X1 port map( A1 => n37728, A2 => REGISTERS_24_0_port, B1 => 
                           n37729, B2 => REGISTERS_1_0_port, ZN => n37117);
   U275 : AOI222_X1 port map( A1 => n37730, A2 => REGISTERS_15_0_port, B1 => 
                           n37731, B2 => REGISTERS_12_0_port, C1 => n37732, C2 
                           => REGISTERS_13_0_port, ZN => n37118);
   U276 : NAND3_X1 port map( A1 => n37116, A2 => n37117, A3 => n37118, ZN => 
                           n37119);
   U277 : AOI22_X1 port map( A1 => n37733, A2 => REGISTERS_22_0_port, B1 => 
                           n37734, B2 => REGISTERS_20_0_port, ZN => n37120);
   U278 : AOI22_X1 port map( A1 => n37735, A2 => REGISTERS_9_0_port, B1 => 
                           n37736, B2 => REGISTERS_18_0_port, ZN => n37121);
   U279 : AOI22_X1 port map( A1 => n37737, A2 => REGISTERS_31_0_port, B1 => 
                           n37738, B2 => REGISTERS_2_0_port, ZN => n37122);
   U280 : AOI22_X1 port map( A1 => n37739, A2 => REGISTERS_8_0_port, B1 => 
                           n37740, B2 => REGISTERS_3_0_port, ZN => n37123);
   U281 : NAND4_X1 port map( A1 => n37120, A2 => n37121, A3 => n37122, A4 => 
                           n37123, ZN => n37124);
   U282 : OR4_X1 port map( A1 => n37110, A2 => n37115, A3 => n37119, A4 => 
                           n37124, ZN => OUTA(0));
   U283 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_31_port, B1 => 
                           n37701, B2 => REGISTERS_16_31_port, ZN => n37125);
   U284 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_31_port, B1 => 
                           n37710, B2 => REGISTERS_6_31_port, ZN => n37126);
   U285 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_31_port, B1 => 
                           n37707, B2 => REGISTERS_24_31_port, ZN => n37127);
   U286 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_31_port, B1 => 
                           n37705, B2 => REGISTERS_12_31_port, ZN => n37128);
   U287 : NAND4_X1 port map( A1 => n37125, A2 => n37126, A3 => n37127, A4 => 
                           n37128, ZN => n37129);
   U288 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_31_port, B1 => 
                           n37703, B2 => REGISTERS_1_31_port, ZN => n37130);
   U289 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_31_port, B1 => 
                           n37699, B2 => REGISTERS_20_31_port, ZN => n37131);
   U290 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_31_port, B1 => 
                           n37700, B2 => REGISTERS_18_31_port, ZN => n37132);
   U291 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_31_port, B1 => 
                           n37718, B2 => REGISTERS_28_31_port, ZN => n37133);
   U292 : NAND4_X1 port map( A1 => n37130, A2 => n37131, A3 => n37132, A4 => 
                           n37133, ZN => n37134);
   U293 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_31_port, B1 => 
                           n37720, B2 => REGISTERS_11_31_port, ZN => n37135);
   U294 : AOI22_X1 port map( A1 => n38277, A2 => REGISTERS_31_31_port, B1 => 
                           n37721, B2 => REGISTERS_2_31_port, ZN => n37136);
   U295 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_31_port, B1 => 
                           n37697, B2 => REGISTERS_13_31_port, C1 => n37722, C2
                           => REGISTERS_19_31_port, ZN => n37137);
   U296 : NAND3_X1 port map( A1 => n37135, A2 => n37136, A3 => n37137, ZN => 
                           n37138);
   U297 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_31_port, B1 => 
                           n37715, B2 => REGISTERS_8_31_port, ZN => n37139);
   U298 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_31_port, B1 => 
                           n37711, B2 => REGISTERS_3_31_port, ZN => n37140);
   U299 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_31_port, B1 => 
                           n37717, B2 => REGISTERS_4_31_port, ZN => n37141);
   U300 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_31_port, B1 => 
                           n38289, B2 => REGISTERS_15_31_port, ZN => n37142);
   U301 : NAND4_X1 port map( A1 => n37139, A2 => n37140, A3 => n37141, A4 => 
                           n37142, ZN => n37143);
   U302 : OR4_X1 port map( A1 => n37129, A2 => n37134, A3 => n37138, A4 => 
                           n37143, ZN => OUTB(31));
   U303 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_4_port, B1 => 
                           n37701, B2 => REGISTERS_16_4_port, ZN => n37144);
   U304 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_4_port, B1 => 
                           n37710, B2 => REGISTERS_6_4_port, ZN => n37145);
   U305 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_4_port, B1 => 
                           n37707, B2 => REGISTERS_24_4_port, ZN => n37146);
   U306 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_4_port, B1 => 
                           n37705, B2 => REGISTERS_12_4_port, ZN => n37147);
   U307 : NAND4_X1 port map( A1 => n37144, A2 => n37145, A3 => n37146, A4 => 
                           n37147, ZN => n37148);
   U308 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_4_port, B1 => 
                           n37703, B2 => REGISTERS_1_4_port, ZN => n37149);
   U309 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_4_port, B1 => 
                           n37699, B2 => REGISTERS_20_4_port, ZN => n37150);
   U310 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_4_port, B1 => 
                           n37700, B2 => REGISTERS_18_4_port, ZN => n37151);
   U311 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_4_port, B1 => 
                           n37718, B2 => REGISTERS_28_4_port, ZN => n37152);
   U312 : NAND4_X1 port map( A1 => n37149, A2 => n37150, A3 => n37151, A4 => 
                           n37152, ZN => n37153);
   U313 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_4_port, B1 => 
                           n37720, B2 => REGISTERS_11_4_port, ZN => n37154);
   U314 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_4_port, B1 => 
                           n38278, B2 => REGISTERS_2_4_port, ZN => n37155);
   U315 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_4_port, B1 => 
                           n37697, B2 => REGISTERS_13_4_port, C1 => n37722, C2 
                           => REGISTERS_19_4_port, ZN => n37156);
   U316 : NAND3_X1 port map( A1 => n37154, A2 => n37155, A3 => n37156, ZN => 
                           n37157);
   U317 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_4_port, B1 => 
                           n37715, B2 => REGISTERS_8_4_port, ZN => n37158);
   U318 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_4_port, B1 => 
                           n37711, B2 => REGISTERS_3_4_port, ZN => n37159);
   U319 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_4_port, B1 => 
                           n37717, B2 => REGISTERS_4_4_port, ZN => n37160);
   U320 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_4_port, B1 => 
                           n37724, B2 => REGISTERS_15_4_port, ZN => n37161);
   U321 : NAND4_X1 port map( A1 => n37158, A2 => n37159, A3 => n37160, A4 => 
                           n37161, ZN => n37162);
   U322 : OR4_X1 port map( A1 => n37148, A2 => n37153, A3 => n37157, A4 => 
                           n37162, ZN => OUTB(4));
   U323 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n38228, B1 => 
                           REGISTERS_30_4_port, B2 => n38229, ZN => n37163);
   U324 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n38230, B1 => 
                           REGISTERS_27_4_port, B2 => n38231, ZN => n37164);
   U325 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n38232, B1 => 
                           REGISTERS_10_4_port, B2 => n38233, ZN => n37165);
   U326 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n38234, B1 => 
                           REGISTERS_6_4_port, B2 => n38235, ZN => n37166);
   U327 : NAND4_X1 port map( A1 => n37163, A2 => n37164, A3 => n37165, A4 => 
                           n37166, ZN => n37167);
   U328 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n38240, B1 => 
                           REGISTERS_26_4_port, B2 => n38241, ZN => n37168);
   U329 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n38242, B1 => 
                           REGISTERS_21_4_port, B2 => n38243, ZN => n37169);
   U330 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n38244, B1 => 
                           REGISTERS_23_4_port, B2 => n38245, ZN => n37170);
   U331 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n38246, B1 => 
                           REGISTERS_14_4_port, B2 => n38247, ZN => n37171);
   U332 : NAND4_X1 port map( A1 => n37168, A2 => n37169, A3 => n37170, A4 => 
                           n37171, ZN => n37172);
   U333 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n38205, B1 => 
                           REGISTERS_11_4_port, B2 => n38206, ZN => n37173);
   U334 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n38207, B1 => 
                           REGISTERS_1_4_port, B2 => n38208, ZN => n37174);
   U335 : AOI222_X1 port map( A1 => REGISTERS_15_4_port, A2 => n38209, B1 => 
                           REGISTERS_12_4_port, B2 => n38210, C1 => 
                           REGISTERS_13_4_port, C2 => n38211, ZN => n37175);
   U336 : NAND3_X1 port map( A1 => n37173, A2 => n37174, A3 => n37175, ZN => 
                           n37176);
   U337 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n38216, B1 => 
                           REGISTERS_20_4_port, B2 => n38217, ZN => n37177);
   U338 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n38218, B1 => 
                           REGISTERS_18_4_port, B2 => n38219, ZN => n37178);
   U339 : AOI22_X1 port map( A1 => REGISTERS_31_4_port, A2 => n38220, B1 => 
                           REGISTERS_2_4_port, B2 => n38221, ZN => n37179);
   U340 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n38222, B1 => 
                           REGISTERS_3_4_port, B2 => n38223, ZN => n37180);
   U341 : NAND4_X1 port map( A1 => n37177, A2 => n37178, A3 => n37179, A4 => 
                           n37180, ZN => n37181);
   U342 : OR4_X1 port map( A1 => n37167, A2 => n37172, A3 => n37176, A4 => 
                           n37181, ZN => OUTA(4));
   U343 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_30_port, B1 => 
                           n37701, B2 => REGISTERS_16_30_port, ZN => n37182);
   U344 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_30_port, B1 => 
                           n37710, B2 => REGISTERS_6_30_port, ZN => n37183);
   U345 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_30_port, B1 => 
                           n37707, B2 => REGISTERS_24_30_port, ZN => n37184);
   U346 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_30_port, B1 => 
                           n37705, B2 => REGISTERS_12_30_port, ZN => n37185);
   U347 : NAND4_X1 port map( A1 => n37182, A2 => n37183, A3 => n37184, A4 => 
                           n37185, ZN => n37186);
   U348 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_30_port, B1 => 
                           n37703, B2 => REGISTERS_1_30_port, ZN => n37187);
   U349 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_30_port, B1 => 
                           n37699, B2 => REGISTERS_20_30_port, ZN => n37188);
   U350 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_30_port, B1 => 
                           n37700, B2 => REGISTERS_18_30_port, ZN => n37189);
   U351 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_30_port, B1 => 
                           n37718, B2 => REGISTERS_28_30_port, ZN => n37190);
   U352 : NAND4_X1 port map( A1 => n37187, A2 => n37188, A3 => n37189, A4 => 
                           n37190, ZN => n37191);
   U353 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_30_port, B1 => 
                           n37720, B2 => REGISTERS_11_30_port, ZN => n37192);
   U354 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_30_port, B1 => 
                           n37721, B2 => REGISTERS_2_30_port, ZN => n37193);
   U355 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_30_port, B1 => 
                           n37697, B2 => REGISTERS_13_30_port, C1 => n37722, C2
                           => REGISTERS_19_30_port, ZN => n37194);
   U356 : NAND3_X1 port map( A1 => n37192, A2 => n37193, A3 => n37194, ZN => 
                           n37195);
   U357 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_30_port, B1 => 
                           n37715, B2 => REGISTERS_8_30_port, ZN => n37196);
   U358 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_30_port, B1 => 
                           n37711, B2 => REGISTERS_3_30_port, ZN => n37197);
   U359 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_30_port, B1 => 
                           n37717, B2 => REGISTERS_4_30_port, ZN => n37198);
   U360 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_30_port, B1 => 
                           n37724, B2 => REGISTERS_15_30_port, ZN => n37199);
   U361 : NAND4_X1 port map( A1 => n37196, A2 => n37197, A3 => n37198, A4 => 
                           n37199, ZN => n37200);
   U362 : OR4_X1 port map( A1 => n37186, A2 => n37191, A3 => n37195, A4 => 
                           n37200, ZN => OUTB(30));
   U363 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_29_port, B1 => 
                           n37701, B2 => REGISTERS_16_29_port, ZN => n37201);
   U364 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_29_port, B1 => 
                           n37710, B2 => REGISTERS_6_29_port, ZN => n37202);
   U365 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_29_port, B1 => 
                           n37707, B2 => REGISTERS_24_29_port, ZN => n37203);
   U366 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_29_port, B1 => 
                           n37705, B2 => REGISTERS_12_29_port, ZN => n37204);
   U367 : NAND4_X1 port map( A1 => n37201, A2 => n37202, A3 => n37203, A4 => 
                           n37204, ZN => n37205);
   U368 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_29_port, B1 => 
                           n37703, B2 => REGISTERS_1_29_port, ZN => n37206);
   U369 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_29_port, B1 => 
                           n37699, B2 => REGISTERS_20_29_port, ZN => n37207);
   U370 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_29_port, B1 => 
                           n37700, B2 => REGISTERS_18_29_port, ZN => n37208);
   U371 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_29_port, B1 => 
                           n37718, B2 => REGISTERS_28_29_port, ZN => n37209);
   U372 : NAND4_X1 port map( A1 => n37206, A2 => n37207, A3 => n37208, A4 => 
                           n37209, ZN => n37210);
   U373 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_29_port, B1 => 
                           n37720, B2 => REGISTERS_11_29_port, ZN => n37211);
   U374 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_29_port, B1 => 
                           n37721, B2 => REGISTERS_2_29_port, ZN => n37212);
   U375 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_29_port, B1 => 
                           n37697, B2 => REGISTERS_13_29_port, C1 => n37722, C2
                           => REGISTERS_19_29_port, ZN => n37213);
   U376 : NAND3_X1 port map( A1 => n37211, A2 => n37212, A3 => n37213, ZN => 
                           n37214);
   U377 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_29_port, B1 => 
                           n37715, B2 => REGISTERS_8_29_port, ZN => n37215);
   U378 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_29_port, B1 => 
                           n37711, B2 => REGISTERS_3_29_port, ZN => n37216);
   U379 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_29_port, B1 => 
                           n37717, B2 => REGISTERS_4_29_port, ZN => n37217);
   U380 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_29_port, B1 => 
                           n37724, B2 => REGISTERS_15_29_port, ZN => n37218);
   U381 : NAND4_X1 port map( A1 => n37215, A2 => n37216, A3 => n37217, A4 => 
                           n37218, ZN => n37219);
   U382 : OR4_X1 port map( A1 => n37205, A2 => n37210, A3 => n37214, A4 => 
                           n37219, ZN => OUTB(29));
   U383 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_28_port, B1 => 
                           n37701, B2 => REGISTERS_16_28_port, ZN => n37220);
   U384 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_28_port, B1 => 
                           n37710, B2 => REGISTERS_6_28_port, ZN => n37221);
   U385 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_28_port, B1 => 
                           n37707, B2 => REGISTERS_24_28_port, ZN => n37222);
   U386 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_28_port, B1 => 
                           n37705, B2 => REGISTERS_12_28_port, ZN => n37223);
   U387 : NAND4_X1 port map( A1 => n37220, A2 => n37221, A3 => n37222, A4 => 
                           n37223, ZN => n37224);
   U388 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_28_port, B1 => 
                           n37703, B2 => REGISTERS_1_28_port, ZN => n37225);
   U389 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_28_port, B1 => 
                           n37699, B2 => REGISTERS_20_28_port, ZN => n37226);
   U390 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_28_port, B1 => 
                           n37700, B2 => REGISTERS_18_28_port, ZN => n37227);
   U391 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_28_port, B1 => 
                           n37718, B2 => REGISTERS_28_28_port, ZN => n37228);
   U392 : NAND4_X1 port map( A1 => n37225, A2 => n37226, A3 => n37227, A4 => 
                           n37228, ZN => n37229);
   U393 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_28_port, B1 => 
                           n37720, B2 => REGISTERS_11_28_port, ZN => n37230);
   U394 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_28_port, B1 => 
                           n37721, B2 => REGISTERS_2_28_port, ZN => n37231);
   U395 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_28_port, B1 => 
                           n37697, B2 => REGISTERS_13_28_port, C1 => n37722, C2
                           => REGISTERS_19_28_port, ZN => n37232);
   U396 : NAND3_X1 port map( A1 => n37230, A2 => n37231, A3 => n37232, ZN => 
                           n37233);
   U397 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_28_port, B1 => 
                           n37715, B2 => REGISTERS_8_28_port, ZN => n37234);
   U398 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_28_port, B1 => 
                           n37711, B2 => REGISTERS_3_28_port, ZN => n37235);
   U399 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_28_port, B1 => 
                           n37717, B2 => REGISTERS_4_28_port, ZN => n37236);
   U400 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_28_port, B1 => 
                           n37724, B2 => REGISTERS_15_28_port, ZN => n37237);
   U401 : NAND4_X1 port map( A1 => n37234, A2 => n37235, A3 => n37236, A4 => 
                           n37237, ZN => n37238);
   U402 : OR4_X1 port map( A1 => n37224, A2 => n37229, A3 => n37233, A4 => 
                           n37238, ZN => OUTB(28));
   U403 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_27_port, B1 => 
                           n37701, B2 => REGISTERS_16_27_port, ZN => n37239);
   U404 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_27_port, B1 => 
                           n37710, B2 => REGISTERS_6_27_port, ZN => n37240);
   U405 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_27_port, B1 => 
                           n37707, B2 => REGISTERS_24_27_port, ZN => n37241);
   U406 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_27_port, B1 => 
                           n37705, B2 => REGISTERS_12_27_port, ZN => n37242);
   U407 : NAND4_X1 port map( A1 => n37239, A2 => n37240, A3 => n37241, A4 => 
                           n37242, ZN => n37243);
   U408 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_27_port, B1 => 
                           n37703, B2 => REGISTERS_1_27_port, ZN => n37244);
   U409 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_27_port, B1 => 
                           n37699, B2 => REGISTERS_20_27_port, ZN => n37245);
   U410 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_27_port, B1 => 
                           n37700, B2 => REGISTERS_18_27_port, ZN => n37246);
   U411 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_27_port, B1 => 
                           n37718, B2 => REGISTERS_28_27_port, ZN => n37247);
   U412 : NAND4_X1 port map( A1 => n37244, A2 => n37245, A3 => n37246, A4 => 
                           n37247, ZN => n37248);
   U413 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_27_port, B1 => 
                           n37720, B2 => REGISTERS_11_27_port, ZN => n37249);
   U414 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_27_port, B1 => 
                           n37721, B2 => REGISTERS_2_27_port, ZN => n37250);
   U415 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_27_port, B1 => 
                           n37697, B2 => REGISTERS_13_27_port, C1 => n37722, C2
                           => REGISTERS_19_27_port, ZN => n37251);
   U416 : NAND3_X1 port map( A1 => n37249, A2 => n37250, A3 => n37251, ZN => 
                           n37252);
   U417 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_27_port, B1 => 
                           n37715, B2 => REGISTERS_8_27_port, ZN => n37253);
   U418 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_27_port, B1 => 
                           n37711, B2 => REGISTERS_3_27_port, ZN => n37254);
   U419 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_27_port, B1 => 
                           n37717, B2 => REGISTERS_4_27_port, ZN => n37255);
   U420 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_27_port, B1 => 
                           n37724, B2 => REGISTERS_15_27_port, ZN => n37256);
   U421 : NAND4_X1 port map( A1 => n37253, A2 => n37254, A3 => n37255, A4 => 
                           n37256, ZN => n37257);
   U422 : OR4_X1 port map( A1 => n37243, A2 => n37248, A3 => n37252, A4 => 
                           n37257, ZN => OUTB(27));
   U423 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_26_port, B1 => 
                           n37701, B2 => REGISTERS_16_26_port, ZN => n37258);
   U424 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_26_port, B1 => 
                           n37710, B2 => REGISTERS_6_26_port, ZN => n37259);
   U425 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_26_port, B1 => 
                           n37707, B2 => REGISTERS_24_26_port, ZN => n37260);
   U426 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_26_port, B1 => 
                           n37705, B2 => REGISTERS_12_26_port, ZN => n37261);
   U427 : NAND4_X1 port map( A1 => n37258, A2 => n37259, A3 => n37260, A4 => 
                           n37261, ZN => n37262);
   U428 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_26_port, B1 => 
                           n37703, B2 => REGISTERS_1_26_port, ZN => n37263);
   U429 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_26_port, B1 => 
                           n37699, B2 => REGISTERS_20_26_port, ZN => n37264);
   U430 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_26_port, B1 => 
                           n37700, B2 => REGISTERS_18_26_port, ZN => n37265);
   U431 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_26_port, B1 => 
                           n37718, B2 => REGISTERS_28_26_port, ZN => n37266);
   U432 : NAND4_X1 port map( A1 => n37263, A2 => n37264, A3 => n37265, A4 => 
                           n37266, ZN => n37267);
   U433 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_26_port, B1 => 
                           n37720, B2 => REGISTERS_11_26_port, ZN => n37268);
   U434 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_26_port, B1 => 
                           n37721, B2 => REGISTERS_2_26_port, ZN => n37269);
   U435 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_26_port, B1 => 
                           n37697, B2 => REGISTERS_13_26_port, C1 => n37722, C2
                           => REGISTERS_19_26_port, ZN => n37270);
   U436 : NAND3_X1 port map( A1 => n37268, A2 => n37269, A3 => n37270, ZN => 
                           n37271);
   U437 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_26_port, B1 => 
                           n37715, B2 => REGISTERS_8_26_port, ZN => n37272);
   U438 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_26_port, B1 => 
                           n37711, B2 => REGISTERS_3_26_port, ZN => n37273);
   U439 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_26_port, B1 => 
                           n37717, B2 => REGISTERS_4_26_port, ZN => n37274);
   U440 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_26_port, B1 => 
                           n37724, B2 => REGISTERS_15_26_port, ZN => n37275);
   U441 : NAND4_X1 port map( A1 => n37272, A2 => n37273, A3 => n37274, A4 => 
                           n37275, ZN => n37276);
   U442 : OR4_X1 port map( A1 => n37262, A2 => n37267, A3 => n37271, A4 => 
                           n37276, ZN => OUTB(26));
   U443 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_25_port, B1 => 
                           n37701, B2 => REGISTERS_16_25_port, ZN => n37277);
   U444 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_25_port, B1 => 
                           n37710, B2 => REGISTERS_6_25_port, ZN => n37278);
   U445 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_25_port, B1 => 
                           n37707, B2 => REGISTERS_24_25_port, ZN => n37279);
   U446 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_25_port, B1 => 
                           n37705, B2 => REGISTERS_12_25_port, ZN => n37280);
   U447 : NAND4_X1 port map( A1 => n37277, A2 => n37278, A3 => n37279, A4 => 
                           n37280, ZN => n37281);
   U448 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_25_port, B1 => 
                           n37703, B2 => REGISTERS_1_25_port, ZN => n37282);
   U449 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_25_port, B1 => 
                           n37699, B2 => REGISTERS_20_25_port, ZN => n37283);
   U450 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_25_port, B1 => 
                           n37700, B2 => REGISTERS_18_25_port, ZN => n37284);
   U451 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_25_port, B1 => 
                           n37718, B2 => REGISTERS_28_25_port, ZN => n37285);
   U452 : NAND4_X1 port map( A1 => n37282, A2 => n37283, A3 => n37284, A4 => 
                           n37285, ZN => n37286);
   U453 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_25_port, B1 => 
                           n37720, B2 => REGISTERS_11_25_port, ZN => n37287);
   U454 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_25_port, B1 => 
                           n37721, B2 => REGISTERS_2_25_port, ZN => n37288);
   U455 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_25_port, B1 => 
                           n37697, B2 => REGISTERS_13_25_port, C1 => n37722, C2
                           => REGISTERS_19_25_port, ZN => n37289);
   U456 : NAND3_X1 port map( A1 => n37287, A2 => n37288, A3 => n37289, ZN => 
                           n37290);
   U457 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_25_port, B1 => 
                           n37715, B2 => REGISTERS_8_25_port, ZN => n37291);
   U458 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_25_port, B1 => 
                           n37711, B2 => REGISTERS_3_25_port, ZN => n37292);
   U459 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_25_port, B1 => 
                           n37717, B2 => REGISTERS_4_25_port, ZN => n37293);
   U460 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_25_port, B1 => 
                           n37724, B2 => REGISTERS_15_25_port, ZN => n37294);
   U461 : NAND4_X1 port map( A1 => n37291, A2 => n37292, A3 => n37293, A4 => 
                           n37294, ZN => n37295);
   U462 : OR4_X1 port map( A1 => n37281, A2 => n37286, A3 => n37290, A4 => 
                           n37295, ZN => OUTB(25));
   U463 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_24_port, B1 => 
                           n37701, B2 => REGISTERS_16_24_port, ZN => n37296);
   U464 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_24_port, B1 => 
                           n37710, B2 => REGISTERS_6_24_port, ZN => n37297);
   U465 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_24_port, B1 => 
                           n37707, B2 => REGISTERS_24_24_port, ZN => n37298);
   U466 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_24_port, B1 => 
                           n37705, B2 => REGISTERS_12_24_port, ZN => n37299);
   U467 : NAND4_X1 port map( A1 => n37296, A2 => n37297, A3 => n37298, A4 => 
                           n37299, ZN => n37300);
   U468 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_24_port, B1 => 
                           n37703, B2 => REGISTERS_1_24_port, ZN => n37301);
   U469 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_24_port, B1 => 
                           n37699, B2 => REGISTERS_20_24_port, ZN => n37302);
   U470 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_24_port, B1 => 
                           n37700, B2 => REGISTERS_18_24_port, ZN => n37303);
   U471 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_24_port, B1 => 
                           n37718, B2 => REGISTERS_28_24_port, ZN => n37304);
   U472 : NAND4_X1 port map( A1 => n37301, A2 => n37302, A3 => n37303, A4 => 
                           n37304, ZN => n37305);
   U473 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_24_port, B1 => 
                           n37720, B2 => REGISTERS_11_24_port, ZN => n37306);
   U474 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_24_port, B1 => 
                           n37721, B2 => REGISTERS_2_24_port, ZN => n37307);
   U475 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_24_port, B1 => 
                           n37697, B2 => REGISTERS_13_24_port, C1 => n37722, C2
                           => REGISTERS_19_24_port, ZN => n37308);
   U476 : NAND3_X1 port map( A1 => n37306, A2 => n37307, A3 => n37308, ZN => 
                           n37309);
   U477 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_24_port, B1 => 
                           n37715, B2 => REGISTERS_8_24_port, ZN => n37310);
   U478 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_24_port, B1 => 
                           n37711, B2 => REGISTERS_3_24_port, ZN => n37311);
   U479 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_24_port, B1 => 
                           n37717, B2 => REGISTERS_4_24_port, ZN => n37312);
   U480 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_24_port, B1 => 
                           n37724, B2 => REGISTERS_15_24_port, ZN => n37313);
   U481 : NAND4_X1 port map( A1 => n37310, A2 => n37311, A3 => n37312, A4 => 
                           n37313, ZN => n37314);
   U482 : OR4_X1 port map( A1 => n37300, A2 => n37305, A3 => n37309, A4 => 
                           n37314, ZN => OUTB(24));
   U483 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_23_port, B1 => 
                           n37701, B2 => REGISTERS_16_23_port, ZN => n37315);
   U484 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_23_port, B1 => 
                           n37710, B2 => REGISTERS_6_23_port, ZN => n37316);
   U485 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_23_port, B1 => 
                           n37707, B2 => REGISTERS_24_23_port, ZN => n37317);
   U486 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_23_port, B1 => 
                           n37705, B2 => REGISTERS_12_23_port, ZN => n37318);
   U487 : NAND4_X1 port map( A1 => n37315, A2 => n37316, A3 => n37317, A4 => 
                           n37318, ZN => n37319);
   U488 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_23_port, B1 => 
                           n37703, B2 => REGISTERS_1_23_port, ZN => n37320);
   U489 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_23_port, B1 => 
                           n37699, B2 => REGISTERS_20_23_port, ZN => n37321);
   U490 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_23_port, B1 => 
                           n37700, B2 => REGISTERS_18_23_port, ZN => n37322);
   U491 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_23_port, B1 => 
                           n37718, B2 => REGISTERS_28_23_port, ZN => n37323);
   U492 : NAND4_X1 port map( A1 => n37320, A2 => n37321, A3 => n37322, A4 => 
                           n37323, ZN => n37324);
   U493 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_23_port, B1 => 
                           n37720, B2 => REGISTERS_11_23_port, ZN => n37325);
   U494 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_23_port, B1 => 
                           n37721, B2 => REGISTERS_2_23_port, ZN => n37326);
   U495 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_23_port, B1 => 
                           n37697, B2 => REGISTERS_13_23_port, C1 => n37722, C2
                           => REGISTERS_19_23_port, ZN => n37327);
   U496 : NAND3_X1 port map( A1 => n37325, A2 => n37326, A3 => n37327, ZN => 
                           n37328);
   U497 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_23_port, B1 => 
                           n37715, B2 => REGISTERS_8_23_port, ZN => n37329);
   U498 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_23_port, B1 => 
                           n37711, B2 => REGISTERS_3_23_port, ZN => n37330);
   U499 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_23_port, B1 => 
                           n37717, B2 => REGISTERS_4_23_port, ZN => n37331);
   U500 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_23_port, B1 => 
                           n37724, B2 => REGISTERS_15_23_port, ZN => n37332);
   U501 : NAND4_X1 port map( A1 => n37329, A2 => n37330, A3 => n37331, A4 => 
                           n37332, ZN => n37333);
   U502 : OR4_X1 port map( A1 => n37319, A2 => n37324, A3 => n37328, A4 => 
                           n37333, ZN => OUTB(23));
   U503 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_22_port, B1 => 
                           n37701, B2 => REGISTERS_16_22_port, ZN => n37334);
   U504 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_22_port, B1 => 
                           n37710, B2 => REGISTERS_6_22_port, ZN => n37335);
   U505 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_22_port, B1 => 
                           n37707, B2 => REGISTERS_24_22_port, ZN => n37336);
   U506 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_22_port, B1 => 
                           n37705, B2 => REGISTERS_12_22_port, ZN => n37337);
   U507 : NAND4_X1 port map( A1 => n37334, A2 => n37335, A3 => n37336, A4 => 
                           n37337, ZN => n37338);
   U508 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_22_port, B1 => 
                           n37703, B2 => REGISTERS_1_22_port, ZN => n37339);
   U509 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_22_port, B1 => 
                           n37699, B2 => REGISTERS_20_22_port, ZN => n37340);
   U510 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_22_port, B1 => 
                           n37700, B2 => REGISTERS_18_22_port, ZN => n37341);
   U511 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_22_port, B1 => 
                           n37718, B2 => REGISTERS_28_22_port, ZN => n37342);
   U512 : NAND4_X1 port map( A1 => n37339, A2 => n37340, A3 => n37341, A4 => 
                           n37342, ZN => n37343);
   U513 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_22_port, B1 => 
                           n37720, B2 => REGISTERS_11_22_port, ZN => n37344);
   U514 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_22_port, B1 => 
                           n37721, B2 => REGISTERS_2_22_port, ZN => n37345);
   U515 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_22_port, B1 => 
                           n37697, B2 => REGISTERS_13_22_port, C1 => n37722, C2
                           => REGISTERS_19_22_port, ZN => n37346);
   U516 : NAND3_X1 port map( A1 => n37344, A2 => n37345, A3 => n37346, ZN => 
                           n37347);
   U517 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_22_port, B1 => 
                           n37715, B2 => REGISTERS_8_22_port, ZN => n37348);
   U518 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_22_port, B1 => 
                           n37711, B2 => REGISTERS_3_22_port, ZN => n37349);
   U519 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_22_port, B1 => 
                           n37717, B2 => REGISTERS_4_22_port, ZN => n37350);
   U520 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_22_port, B1 => 
                           n37724, B2 => REGISTERS_15_22_port, ZN => n37351);
   U521 : NAND4_X1 port map( A1 => n37348, A2 => n37349, A3 => n37350, A4 => 
                           n37351, ZN => n37352);
   U522 : OR4_X1 port map( A1 => n37338, A2 => n37343, A3 => n37347, A4 => 
                           n37352, ZN => OUTB(22));
   U523 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_21_port, B1 => 
                           n37701, B2 => REGISTERS_16_21_port, ZN => n37353);
   U524 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_21_port, B1 => 
                           n37710, B2 => REGISTERS_6_21_port, ZN => n37354);
   U525 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_21_port, B1 => 
                           n37707, B2 => REGISTERS_24_21_port, ZN => n37355);
   U526 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_21_port, B1 => 
                           n37705, B2 => REGISTERS_12_21_port, ZN => n37356);
   U527 : NAND4_X1 port map( A1 => n37353, A2 => n37354, A3 => n37355, A4 => 
                           n37356, ZN => n37357);
   U528 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_21_port, B1 => 
                           n37703, B2 => REGISTERS_1_21_port, ZN => n37358);
   U529 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_21_port, B1 => 
                           n37699, B2 => REGISTERS_20_21_port, ZN => n37359);
   U530 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_21_port, B1 => 
                           n37700, B2 => REGISTERS_18_21_port, ZN => n37360);
   U531 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_21_port, B1 => 
                           n37718, B2 => REGISTERS_28_21_port, ZN => n37361);
   U532 : NAND4_X1 port map( A1 => n37358, A2 => n37359, A3 => n37360, A4 => 
                           n37361, ZN => n37362);
   U533 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_21_port, B1 => 
                           n37720, B2 => REGISTERS_11_21_port, ZN => n37363);
   U534 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_21_port, B1 => 
                           n37721, B2 => REGISTERS_2_21_port, ZN => n37364);
   U535 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_21_port, B1 => 
                           n37697, B2 => REGISTERS_13_21_port, C1 => n37722, C2
                           => REGISTERS_19_21_port, ZN => n37365);
   U536 : NAND3_X1 port map( A1 => n37363, A2 => n37364, A3 => n37365, ZN => 
                           n37366);
   U537 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_21_port, B1 => 
                           n37715, B2 => REGISTERS_8_21_port, ZN => n37367);
   U538 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_21_port, B1 => 
                           n37711, B2 => REGISTERS_3_21_port, ZN => n37368);
   U539 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_21_port, B1 => 
                           n37717, B2 => REGISTERS_4_21_port, ZN => n37369);
   U540 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_21_port, B1 => 
                           n37724, B2 => REGISTERS_15_21_port, ZN => n37370);
   U541 : NAND4_X1 port map( A1 => n37367, A2 => n37368, A3 => n37369, A4 => 
                           n37370, ZN => n37371);
   U542 : OR4_X1 port map( A1 => n37357, A2 => n37362, A3 => n37366, A4 => 
                           n37371, ZN => OUTB(21));
   U543 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_20_port, B1 => 
                           n37701, B2 => REGISTERS_16_20_port, ZN => n37372);
   U544 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_20_port, B1 => 
                           n37710, B2 => REGISTERS_6_20_port, ZN => n37373);
   U545 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_20_port, B1 => 
                           n37707, B2 => REGISTERS_24_20_port, ZN => n37374);
   U546 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_20_port, B1 => 
                           n37705, B2 => REGISTERS_12_20_port, ZN => n37375);
   U547 : NAND4_X1 port map( A1 => n37372, A2 => n37373, A3 => n37374, A4 => 
                           n37375, ZN => n37376);
   U548 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_20_port, B1 => 
                           n37703, B2 => REGISTERS_1_20_port, ZN => n37377);
   U549 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_20_port, B1 => 
                           n37699, B2 => REGISTERS_20_20_port, ZN => n37378);
   U550 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_20_port, B1 => 
                           n37700, B2 => REGISTERS_18_20_port, ZN => n37379);
   U551 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_20_port, B1 => 
                           n37718, B2 => REGISTERS_28_20_port, ZN => n37380);
   U552 : NAND4_X1 port map( A1 => n37377, A2 => n37378, A3 => n37379, A4 => 
                           n37380, ZN => n37381);
   U553 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_20_port, B1 => 
                           n37720, B2 => REGISTERS_11_20_port, ZN => n37382);
   U554 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_20_port, B1 => 
                           n37721, B2 => REGISTERS_2_20_port, ZN => n37383);
   U555 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_20_port, B1 => 
                           n37697, B2 => REGISTERS_13_20_port, C1 => n37722, C2
                           => REGISTERS_19_20_port, ZN => n37384);
   U556 : NAND3_X1 port map( A1 => n37382, A2 => n37383, A3 => n37384, ZN => 
                           n37385);
   U557 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_20_port, B1 => 
                           n37715, B2 => REGISTERS_8_20_port, ZN => n37386);
   U558 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_20_port, B1 => 
                           n37711, B2 => REGISTERS_3_20_port, ZN => n37387);
   U559 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_20_port, B1 => 
                           n37717, B2 => REGISTERS_4_20_port, ZN => n37388);
   U560 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_20_port, B1 => 
                           n37724, B2 => REGISTERS_15_20_port, ZN => n37389);
   U561 : NAND4_X1 port map( A1 => n37386, A2 => n37387, A3 => n37388, A4 => 
                           n37389, ZN => n37390);
   U562 : OR4_X1 port map( A1 => n37376, A2 => n37381, A3 => n37385, A4 => 
                           n37390, ZN => OUTB(20));
   U563 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_19_port, B1 => 
                           n37701, B2 => REGISTERS_16_19_port, ZN => n37391);
   U564 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_19_port, B1 => 
                           n37710, B2 => REGISTERS_6_19_port, ZN => n37392);
   U565 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_19_port, B1 => 
                           n37707, B2 => REGISTERS_24_19_port, ZN => n37393);
   U566 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_19_port, B1 => 
                           n37705, B2 => REGISTERS_12_19_port, ZN => n37394);
   U567 : NAND4_X1 port map( A1 => n37391, A2 => n37392, A3 => n37393, A4 => 
                           n37394, ZN => n37395);
   U568 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_19_port, B1 => 
                           n37703, B2 => REGISTERS_1_19_port, ZN => n37396);
   U569 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_19_port, B1 => 
                           n37699, B2 => REGISTERS_20_19_port, ZN => n37397);
   U570 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_19_port, B1 => 
                           n37700, B2 => REGISTERS_18_19_port, ZN => n37398);
   U571 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_19_port, B1 => 
                           n37718, B2 => REGISTERS_28_19_port, ZN => n37399);
   U572 : NAND4_X1 port map( A1 => n37396, A2 => n37397, A3 => n37398, A4 => 
                           n37399, ZN => n37400);
   U573 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_19_port, B1 => 
                           n37720, B2 => REGISTERS_11_19_port, ZN => n37401);
   U574 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_19_port, B1 => 
                           n37721, B2 => REGISTERS_2_19_port, ZN => n37402);
   U575 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_19_port, B1 => 
                           n37697, B2 => REGISTERS_13_19_port, C1 => n37722, C2
                           => REGISTERS_19_19_port, ZN => n37403);
   U576 : NAND3_X1 port map( A1 => n37401, A2 => n37402, A3 => n37403, ZN => 
                           n37404);
   U577 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_19_port, B1 => 
                           n37715, B2 => REGISTERS_8_19_port, ZN => n37405);
   U578 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_19_port, B1 => 
                           n37711, B2 => REGISTERS_3_19_port, ZN => n37406);
   U579 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_19_port, B1 => 
                           n37717, B2 => REGISTERS_4_19_port, ZN => n37407);
   U580 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_19_port, B1 => 
                           n37724, B2 => REGISTERS_15_19_port, ZN => n37408);
   U581 : NAND4_X1 port map( A1 => n37405, A2 => n37406, A3 => n37407, A4 => 
                           n37408, ZN => n37409);
   U582 : OR4_X1 port map( A1 => n37395, A2 => n37400, A3 => n37404, A4 => 
                           n37409, ZN => OUTB(19));
   U583 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_18_port, B1 => 
                           n37701, B2 => REGISTERS_16_18_port, ZN => n37410);
   U584 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_18_port, B1 => 
                           n37710, B2 => REGISTERS_6_18_port, ZN => n37411);
   U585 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_18_port, B1 => 
                           n37707, B2 => REGISTERS_24_18_port, ZN => n37412);
   U586 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_18_port, B1 => 
                           n37705, B2 => REGISTERS_12_18_port, ZN => n37413);
   U587 : NAND4_X1 port map( A1 => n37410, A2 => n37411, A3 => n37412, A4 => 
                           n37413, ZN => n37414);
   U588 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_18_port, B1 => 
                           n37703, B2 => REGISTERS_1_18_port, ZN => n37415);
   U589 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_18_port, B1 => 
                           n37699, B2 => REGISTERS_20_18_port, ZN => n37416);
   U590 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_18_port, B1 => 
                           n37700, B2 => REGISTERS_18_18_port, ZN => n37417);
   U591 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_18_port, B1 => 
                           n37718, B2 => REGISTERS_28_18_port, ZN => n37418);
   U592 : NAND4_X1 port map( A1 => n37415, A2 => n37416, A3 => n37417, A4 => 
                           n37418, ZN => n37419);
   U593 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_18_port, B1 => 
                           n37720, B2 => REGISTERS_11_18_port, ZN => n37420);
   U594 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_18_port, B1 => 
                           n37721, B2 => REGISTERS_2_18_port, ZN => n37421);
   U595 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_18_port, B1 => 
                           n37697, B2 => REGISTERS_13_18_port, C1 => n37722, C2
                           => REGISTERS_19_18_port, ZN => n37422);
   U596 : NAND3_X1 port map( A1 => n37420, A2 => n37421, A3 => n37422, ZN => 
                           n37423);
   U597 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_18_port, B1 => 
                           n37715, B2 => REGISTERS_8_18_port, ZN => n37424);
   U598 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_18_port, B1 => 
                           n37711, B2 => REGISTERS_3_18_port, ZN => n37425);
   U599 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_18_port, B1 => 
                           n37717, B2 => REGISTERS_4_18_port, ZN => n37426);
   U600 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_18_port, B1 => 
                           n37724, B2 => REGISTERS_15_18_port, ZN => n37427);
   U601 : NAND4_X1 port map( A1 => n37424, A2 => n37425, A3 => n37426, A4 => 
                           n37427, ZN => n37428);
   U602 : OR4_X1 port map( A1 => n37414, A2 => n37419, A3 => n37423, A4 => 
                           n37428, ZN => OUTB(18));
   U603 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_17_port, B1 => 
                           n37701, B2 => REGISTERS_16_17_port, ZN => n37429);
   U604 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_17_port, B1 => 
                           n37710, B2 => REGISTERS_6_17_port, ZN => n37430);
   U605 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_17_port, B1 => 
                           n37707, B2 => REGISTERS_24_17_port, ZN => n37431);
   U606 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_17_port, B1 => 
                           n37705, B2 => REGISTERS_12_17_port, ZN => n37432);
   U607 : NAND4_X1 port map( A1 => n37429, A2 => n37430, A3 => n37431, A4 => 
                           n37432, ZN => n37433);
   U608 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_17_port, B1 => 
                           n37703, B2 => REGISTERS_1_17_port, ZN => n37434);
   U609 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_17_port, B1 => 
                           n37699, B2 => REGISTERS_20_17_port, ZN => n37435);
   U610 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_17_port, B1 => 
                           n37700, B2 => REGISTERS_18_17_port, ZN => n37436);
   U611 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_17_port, B1 => 
                           n37718, B2 => REGISTERS_28_17_port, ZN => n37437);
   U612 : NAND4_X1 port map( A1 => n37434, A2 => n37435, A3 => n37436, A4 => 
                           n37437, ZN => n37438);
   U613 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_17_port, B1 => 
                           n37720, B2 => REGISTERS_11_17_port, ZN => n37439);
   U614 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_17_port, B1 => 
                           n37721, B2 => REGISTERS_2_17_port, ZN => n37440);
   U615 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_17_port, B1 => 
                           n37697, B2 => REGISTERS_13_17_port, C1 => n37722, C2
                           => REGISTERS_19_17_port, ZN => n37441);
   U616 : NAND3_X1 port map( A1 => n37439, A2 => n37440, A3 => n37441, ZN => 
                           n37442);
   U617 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_17_port, B1 => 
                           n37715, B2 => REGISTERS_8_17_port, ZN => n37443);
   U618 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_17_port, B1 => 
                           n37711, B2 => REGISTERS_3_17_port, ZN => n37444);
   U619 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_17_port, B1 => 
                           n37717, B2 => REGISTERS_4_17_port, ZN => n37445);
   U620 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_17_port, B1 => 
                           n37724, B2 => REGISTERS_15_17_port, ZN => n37446);
   U621 : NAND4_X1 port map( A1 => n37443, A2 => n37444, A3 => n37445, A4 => 
                           n37446, ZN => n37447);
   U622 : OR4_X1 port map( A1 => n37433, A2 => n37438, A3 => n37442, A4 => 
                           n37447, ZN => OUTB(17));
   U623 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_16_port, B1 => 
                           n37701, B2 => REGISTERS_16_16_port, ZN => n37448);
   U624 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_16_port, B1 => 
                           n37710, B2 => REGISTERS_6_16_port, ZN => n37449);
   U625 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_16_port, B1 => 
                           n37707, B2 => REGISTERS_24_16_port, ZN => n37450);
   U626 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_16_port, B1 => 
                           n37705, B2 => REGISTERS_12_16_port, ZN => n37451);
   U627 : NAND4_X1 port map( A1 => n37448, A2 => n37449, A3 => n37450, A4 => 
                           n37451, ZN => n37452);
   U628 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_16_port, B1 => 
                           n37703, B2 => REGISTERS_1_16_port, ZN => n37453);
   U629 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_16_port, B1 => 
                           n37699, B2 => REGISTERS_20_16_port, ZN => n37454);
   U630 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_16_port, B1 => 
                           n37700, B2 => REGISTERS_18_16_port, ZN => n37455);
   U631 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_16_port, B1 => 
                           n37718, B2 => REGISTERS_28_16_port, ZN => n37456);
   U632 : NAND4_X1 port map( A1 => n37453, A2 => n37454, A3 => n37455, A4 => 
                           n37456, ZN => n37457);
   U633 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_16_port, B1 => 
                           n37720, B2 => REGISTERS_11_16_port, ZN => n37458);
   U634 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_16_port, B1 => 
                           n37721, B2 => REGISTERS_2_16_port, ZN => n37459);
   U635 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_16_port, B1 => 
                           n37697, B2 => REGISTERS_13_16_port, C1 => n37722, C2
                           => REGISTERS_19_16_port, ZN => n37460);
   U636 : NAND3_X1 port map( A1 => n37458, A2 => n37459, A3 => n37460, ZN => 
                           n37461);
   U637 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_16_port, B1 => 
                           n37715, B2 => REGISTERS_8_16_port, ZN => n37462);
   U638 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_16_port, B1 => 
                           n37711, B2 => REGISTERS_3_16_port, ZN => n37463);
   U639 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_16_port, B1 => 
                           n37717, B2 => REGISTERS_4_16_port, ZN => n37464);
   U640 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_16_port, B1 => 
                           n37724, B2 => REGISTERS_15_16_port, ZN => n37465);
   U641 : NAND4_X1 port map( A1 => n37462, A2 => n37463, A3 => n37464, A4 => 
                           n37465, ZN => n37466);
   U642 : OR4_X1 port map( A1 => n37452, A2 => n37457, A3 => n37461, A4 => 
                           n37466, ZN => OUTB(16));
   U643 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_15_port, B1 => 
                           n37701, B2 => REGISTERS_16_15_port, ZN => n37467);
   U644 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_15_port, B1 => 
                           n37710, B2 => REGISTERS_6_15_port, ZN => n37468);
   U645 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_15_port, B1 => 
                           n37707, B2 => REGISTERS_24_15_port, ZN => n37469);
   U646 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_15_port, B1 => 
                           n37705, B2 => REGISTERS_12_15_port, ZN => n37470);
   U647 : NAND4_X1 port map( A1 => n37467, A2 => n37468, A3 => n37469, A4 => 
                           n37470, ZN => n37471);
   U648 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_15_port, B1 => 
                           n37703, B2 => REGISTERS_1_15_port, ZN => n37472);
   U649 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_15_port, B1 => 
                           n37699, B2 => REGISTERS_20_15_port, ZN => n37473);
   U650 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_15_port, B1 => 
                           n37700, B2 => REGISTERS_18_15_port, ZN => n37474);
   U651 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_15_port, B1 => 
                           n37718, B2 => REGISTERS_28_15_port, ZN => n37475);
   U652 : NAND4_X1 port map( A1 => n37472, A2 => n37473, A3 => n37474, A4 => 
                           n37475, ZN => n37476);
   U653 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_15_port, B1 => 
                           n37720, B2 => REGISTERS_11_15_port, ZN => n37477);
   U654 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_15_port, B1 => 
                           n37721, B2 => REGISTERS_2_15_port, ZN => n37478);
   U655 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_15_port, B1 => 
                           n37697, B2 => REGISTERS_13_15_port, C1 => n37722, C2
                           => REGISTERS_19_15_port, ZN => n37479);
   U656 : NAND3_X1 port map( A1 => n37477, A2 => n37478, A3 => n37479, ZN => 
                           n37480);
   U657 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_15_port, B1 => 
                           n37715, B2 => REGISTERS_8_15_port, ZN => n37481);
   U658 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_15_port, B1 => 
                           n37711, B2 => REGISTERS_3_15_port, ZN => n37482);
   U659 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_15_port, B1 => 
                           n37717, B2 => REGISTERS_4_15_port, ZN => n37483);
   U660 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_15_port, B1 => 
                           n37724, B2 => REGISTERS_15_15_port, ZN => n37484);
   U661 : NAND4_X1 port map( A1 => n37481, A2 => n37482, A3 => n37483, A4 => 
                           n37484, ZN => n37485);
   U662 : OR4_X1 port map( A1 => n37471, A2 => n37476, A3 => n37480, A4 => 
                           n37485, ZN => OUTB(15));
   U663 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_14_port, B1 => 
                           n37701, B2 => REGISTERS_16_14_port, ZN => n37486);
   U664 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_14_port, B1 => 
                           n37710, B2 => REGISTERS_6_14_port, ZN => n37487);
   U665 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_14_port, B1 => 
                           n37707, B2 => REGISTERS_24_14_port, ZN => n37488);
   U666 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_14_port, B1 => 
                           n37705, B2 => REGISTERS_12_14_port, ZN => n37489);
   U667 : NAND4_X1 port map( A1 => n37486, A2 => n37487, A3 => n37488, A4 => 
                           n37489, ZN => n37490);
   U668 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_14_port, B1 => 
                           n37703, B2 => REGISTERS_1_14_port, ZN => n37491);
   U669 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_14_port, B1 => 
                           n37699, B2 => REGISTERS_20_14_port, ZN => n37492);
   U670 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_14_port, B1 => 
                           n37700, B2 => REGISTERS_18_14_port, ZN => n37493);
   U671 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_14_port, B1 => 
                           n37718, B2 => REGISTERS_28_14_port, ZN => n37494);
   U672 : NAND4_X1 port map( A1 => n37491, A2 => n37492, A3 => n37493, A4 => 
                           n37494, ZN => n37495);
   U673 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_14_port, B1 => 
                           n37720, B2 => REGISTERS_11_14_port, ZN => n37496);
   U674 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_14_port, B1 => 
                           n37721, B2 => REGISTERS_2_14_port, ZN => n37497);
   U675 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_14_port, B1 => 
                           n37697, B2 => REGISTERS_13_14_port, C1 => n37722, C2
                           => REGISTERS_19_14_port, ZN => n37498);
   U676 : NAND3_X1 port map( A1 => n37496, A2 => n37497, A3 => n37498, ZN => 
                           n37499);
   U677 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_14_port, B1 => 
                           n37715, B2 => REGISTERS_8_14_port, ZN => n37500);
   U678 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_14_port, B1 => 
                           n37711, B2 => REGISTERS_3_14_port, ZN => n37501);
   U679 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_14_port, B1 => 
                           n37717, B2 => REGISTERS_4_14_port, ZN => n37502);
   U680 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_14_port, B1 => 
                           n37724, B2 => REGISTERS_15_14_port, ZN => n37503);
   U681 : NAND4_X1 port map( A1 => n37500, A2 => n37501, A3 => n37502, A4 => 
                           n37503, ZN => n37504);
   U682 : OR4_X1 port map( A1 => n37490, A2 => n37495, A3 => n37499, A4 => 
                           n37504, ZN => OUTB(14));
   U683 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_13_port, B1 => 
                           n37701, B2 => REGISTERS_16_13_port, ZN => n37505);
   U684 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_13_port, B1 => 
                           n37710, B2 => REGISTERS_6_13_port, ZN => n37506);
   U685 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_13_port, B1 => 
                           n37707, B2 => REGISTERS_24_13_port, ZN => n37507);
   U686 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_13_port, B1 => 
                           n37705, B2 => REGISTERS_12_13_port, ZN => n37508);
   U687 : NAND4_X1 port map( A1 => n37505, A2 => n37506, A3 => n37507, A4 => 
                           n37508, ZN => n37509);
   U688 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_13_port, B1 => 
                           n37703, B2 => REGISTERS_1_13_port, ZN => n37510);
   U689 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_13_port, B1 => 
                           n37699, B2 => REGISTERS_20_13_port, ZN => n37511);
   U690 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_13_port, B1 => 
                           n37700, B2 => REGISTERS_18_13_port, ZN => n37512);
   U691 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_13_port, B1 => 
                           n37718, B2 => REGISTERS_28_13_port, ZN => n37513);
   U692 : NAND4_X1 port map( A1 => n37510, A2 => n37511, A3 => n37512, A4 => 
                           n37513, ZN => n37514);
   U693 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_13_port, B1 => 
                           n37720, B2 => REGISTERS_11_13_port, ZN => n37515);
   U694 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_13_port, B1 => 
                           n37721, B2 => REGISTERS_2_13_port, ZN => n37516);
   U695 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_13_port, B1 => 
                           n37697, B2 => REGISTERS_13_13_port, C1 => n37722, C2
                           => REGISTERS_19_13_port, ZN => n37517);
   U696 : NAND3_X1 port map( A1 => n37515, A2 => n37516, A3 => n37517, ZN => 
                           n37518);
   U697 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_13_port, B1 => 
                           n37715, B2 => REGISTERS_8_13_port, ZN => n37519);
   U698 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_13_port, B1 => 
                           n37711, B2 => REGISTERS_3_13_port, ZN => n37520);
   U699 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_13_port, B1 => 
                           n37717, B2 => REGISTERS_4_13_port, ZN => n37521);
   U700 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_13_port, B1 => 
                           n37724, B2 => REGISTERS_15_13_port, ZN => n37522);
   U701 : NAND4_X1 port map( A1 => n37519, A2 => n37520, A3 => n37521, A4 => 
                           n37522, ZN => n37523);
   U702 : OR4_X1 port map( A1 => n37509, A2 => n37514, A3 => n37518, A4 => 
                           n37523, ZN => OUTB(13));
   U703 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_12_port, B1 => 
                           n37701, B2 => REGISTERS_16_12_port, ZN => n37524);
   U704 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_12_port, B1 => 
                           n37710, B2 => REGISTERS_6_12_port, ZN => n37525);
   U705 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_12_port, B1 => 
                           n37707, B2 => REGISTERS_24_12_port, ZN => n37526);
   U706 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_12_port, B1 => 
                           n37705, B2 => REGISTERS_12_12_port, ZN => n37527);
   U707 : NAND4_X1 port map( A1 => n37524, A2 => n37525, A3 => n37526, A4 => 
                           n37527, ZN => n37528);
   U708 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_12_port, B1 => 
                           n37703, B2 => REGISTERS_1_12_port, ZN => n37529);
   U709 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_12_port, B1 => 
                           n37699, B2 => REGISTERS_20_12_port, ZN => n37530);
   U710 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_12_port, B1 => 
                           n37700, B2 => REGISTERS_18_12_port, ZN => n37531);
   U711 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_12_port, B1 => 
                           n37718, B2 => REGISTERS_28_12_port, ZN => n37532);
   U712 : NAND4_X1 port map( A1 => n37529, A2 => n37530, A3 => n37531, A4 => 
                           n37532, ZN => n37533);
   U713 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_12_port, B1 => 
                           n37720, B2 => REGISTERS_11_12_port, ZN => n37534);
   U714 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_12_port, B1 => 
                           n37721, B2 => REGISTERS_2_12_port, ZN => n37535);
   U715 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_12_port, B1 => 
                           n37697, B2 => REGISTERS_13_12_port, C1 => n37722, C2
                           => REGISTERS_19_12_port, ZN => n37536);
   U716 : NAND3_X1 port map( A1 => n37534, A2 => n37535, A3 => n37536, ZN => 
                           n37537);
   U717 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_12_port, B1 => 
                           n37715, B2 => REGISTERS_8_12_port, ZN => n37538);
   U718 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_12_port, B1 => 
                           n37711, B2 => REGISTERS_3_12_port, ZN => n37539);
   U719 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_12_port, B1 => 
                           n37717, B2 => REGISTERS_4_12_port, ZN => n37540);
   U720 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_12_port, B1 => 
                           n37724, B2 => REGISTERS_15_12_port, ZN => n37541);
   U721 : NAND4_X1 port map( A1 => n37538, A2 => n37539, A3 => n37540, A4 => 
                           n37541, ZN => n37542);
   U722 : OR4_X1 port map( A1 => n37528, A2 => n37533, A3 => n37537, A4 => 
                           n37542, ZN => OUTB(12));
   U723 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_11_port, B1 => 
                           n37701, B2 => REGISTERS_16_11_port, ZN => n37543);
   U724 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_11_port, B1 => 
                           n37710, B2 => REGISTERS_6_11_port, ZN => n37544);
   U725 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_11_port, B1 => 
                           n37707, B2 => REGISTERS_24_11_port, ZN => n37545);
   U726 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_11_port, B1 => 
                           n37705, B2 => REGISTERS_12_11_port, ZN => n37546);
   U727 : NAND4_X1 port map( A1 => n37543, A2 => n37544, A3 => n37545, A4 => 
                           n37546, ZN => n37547);
   U728 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_11_port, B1 => 
                           n37703, B2 => REGISTERS_1_11_port, ZN => n37548);
   U729 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_11_port, B1 => 
                           n37699, B2 => REGISTERS_20_11_port, ZN => n37549);
   U730 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_11_port, B1 => 
                           n37700, B2 => REGISTERS_18_11_port, ZN => n37550);
   U731 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_11_port, B1 => 
                           n37718, B2 => REGISTERS_28_11_port, ZN => n37551);
   U732 : NAND4_X1 port map( A1 => n37548, A2 => n37549, A3 => n37550, A4 => 
                           n37551, ZN => n37552);
   U733 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_11_port, B1 => 
                           n37720, B2 => REGISTERS_11_11_port, ZN => n37553);
   U734 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_11_port, B1 => 
                           n37721, B2 => REGISTERS_2_11_port, ZN => n37554);
   U735 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_11_port, B1 => 
                           n37697, B2 => REGISTERS_13_11_port, C1 => n37722, C2
                           => REGISTERS_19_11_port, ZN => n37555);
   U736 : NAND3_X1 port map( A1 => n37553, A2 => n37554, A3 => n37555, ZN => 
                           n37556);
   U737 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_11_port, B1 => 
                           n37715, B2 => REGISTERS_8_11_port, ZN => n37557);
   U738 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_11_port, B1 => 
                           n37711, B2 => REGISTERS_3_11_port, ZN => n37558);
   U739 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_11_port, B1 => 
                           n37717, B2 => REGISTERS_4_11_port, ZN => n37559);
   U740 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_11_port, B1 => 
                           n37724, B2 => REGISTERS_15_11_port, ZN => n37560);
   U741 : NAND4_X1 port map( A1 => n37557, A2 => n37558, A3 => n37559, A4 => 
                           n37560, ZN => n37561);
   U742 : OR4_X1 port map( A1 => n37547, A2 => n37552, A3 => n37556, A4 => 
                           n37561, ZN => OUTB(11));
   U743 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_10_port, B1 => 
                           n37701, B2 => REGISTERS_16_10_port, ZN => n37562);
   U744 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_10_port, B1 => 
                           n37710, B2 => REGISTERS_6_10_port, ZN => n37563);
   U745 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_10_port, B1 => 
                           n37707, B2 => REGISTERS_24_10_port, ZN => n37564);
   U746 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_10_port, B1 => 
                           n37705, B2 => REGISTERS_12_10_port, ZN => n37565);
   U747 : NAND4_X1 port map( A1 => n37562, A2 => n37563, A3 => n37564, A4 => 
                           n37565, ZN => n37566);
   U748 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_10_port, B1 => 
                           n37703, B2 => REGISTERS_1_10_port, ZN => n37567);
   U749 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_10_port, B1 => 
                           n37699, B2 => REGISTERS_20_10_port, ZN => n37568);
   U750 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_10_port, B1 => 
                           n37700, B2 => REGISTERS_18_10_port, ZN => n37569);
   U751 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_10_port, B1 => 
                           n37718, B2 => REGISTERS_28_10_port, ZN => n37570);
   U752 : NAND4_X1 port map( A1 => n37567, A2 => n37568, A3 => n37569, A4 => 
                           n37570, ZN => n37571);
   U753 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_10_port, B1 => 
                           n37720, B2 => REGISTERS_11_10_port, ZN => n37572);
   U754 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_10_port, B1 => 
                           n37721, B2 => REGISTERS_2_10_port, ZN => n37573);
   U755 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_10_port, B1 => 
                           n37697, B2 => REGISTERS_13_10_port, C1 => n37722, C2
                           => REGISTERS_19_10_port, ZN => n37574);
   U756 : NAND3_X1 port map( A1 => n37572, A2 => n37573, A3 => n37574, ZN => 
                           n37575);
   U757 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_10_port, B1 => 
                           n37715, B2 => REGISTERS_8_10_port, ZN => n37576);
   U758 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_10_port, B1 => 
                           n37711, B2 => REGISTERS_3_10_port, ZN => n37577);
   U759 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_10_port, B1 => 
                           n37717, B2 => REGISTERS_4_10_port, ZN => n37578);
   U760 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_10_port, B1 => 
                           n37724, B2 => REGISTERS_15_10_port, ZN => n37579);
   U761 : NAND4_X1 port map( A1 => n37576, A2 => n37577, A3 => n37578, A4 => 
                           n37579, ZN => n37580);
   U762 : OR4_X1 port map( A1 => n37566, A2 => n37571, A3 => n37575, A4 => 
                           n37580, ZN => OUTB(10));
   U763 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_9_port, B1 => 
                           n37701, B2 => REGISTERS_16_9_port, ZN => n37581);
   U764 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_9_port, B1 => 
                           n37710, B2 => REGISTERS_6_9_port, ZN => n37582);
   U765 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_9_port, B1 => 
                           n37707, B2 => REGISTERS_24_9_port, ZN => n37583);
   U766 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_9_port, B1 => 
                           n37705, B2 => REGISTERS_12_9_port, ZN => n37584);
   U767 : NAND4_X1 port map( A1 => n37581, A2 => n37582, A3 => n37583, A4 => 
                           n37584, ZN => n37585);
   U768 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_9_port, B1 => 
                           n37703, B2 => REGISTERS_1_9_port, ZN => n37586);
   U769 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_9_port, B1 => 
                           n37699, B2 => REGISTERS_20_9_port, ZN => n37587);
   U770 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_9_port, B1 => 
                           n37700, B2 => REGISTERS_18_9_port, ZN => n37588);
   U771 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_9_port, B1 => 
                           n37718, B2 => REGISTERS_28_9_port, ZN => n37589);
   U772 : NAND4_X1 port map( A1 => n37586, A2 => n37587, A3 => n37588, A4 => 
                           n37589, ZN => n37590);
   U773 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_9_port, B1 => 
                           n37720, B2 => REGISTERS_11_9_port, ZN => n37591);
   U774 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_9_port, B1 => 
                           n37721, B2 => REGISTERS_2_9_port, ZN => n37592);
   U775 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_9_port, B1 => 
                           n37697, B2 => REGISTERS_13_9_port, C1 => n37722, C2 
                           => REGISTERS_19_9_port, ZN => n37593);
   U776 : NAND3_X1 port map( A1 => n37591, A2 => n37592, A3 => n37593, ZN => 
                           n37594);
   U777 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_9_port, B1 => 
                           n37715, B2 => REGISTERS_8_9_port, ZN => n37595);
   U778 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_9_port, B1 => 
                           n37711, B2 => REGISTERS_3_9_port, ZN => n37596);
   U779 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_9_port, B1 => 
                           n37717, B2 => REGISTERS_4_9_port, ZN => n37597);
   U780 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_9_port, B1 => 
                           n37724, B2 => REGISTERS_15_9_port, ZN => n37598);
   U781 : NAND4_X1 port map( A1 => n37595, A2 => n37596, A3 => n37597, A4 => 
                           n37598, ZN => n37599);
   U782 : OR4_X1 port map( A1 => n37585, A2 => n37590, A3 => n37594, A4 => 
                           n37599, ZN => OUTB(9));
   U783 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_8_port, B1 => 
                           n37701, B2 => REGISTERS_16_8_port, ZN => n37600);
   U784 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_8_port, B1 => 
                           n37710, B2 => REGISTERS_6_8_port, ZN => n37601);
   U785 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_8_port, B1 => 
                           n37707, B2 => REGISTERS_24_8_port, ZN => n37602);
   U786 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_8_port, B1 => 
                           n37705, B2 => REGISTERS_12_8_port, ZN => n37603);
   U787 : NAND4_X1 port map( A1 => n37600, A2 => n37601, A3 => n37602, A4 => 
                           n37603, ZN => n37604);
   U788 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_8_port, B1 => 
                           n37703, B2 => REGISTERS_1_8_port, ZN => n37605);
   U789 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_8_port, B1 => 
                           n37699, B2 => REGISTERS_20_8_port, ZN => n37606);
   U790 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_8_port, B1 => 
                           n37700, B2 => REGISTERS_18_8_port, ZN => n37607);
   U791 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_8_port, B1 => 
                           n37718, B2 => REGISTERS_28_8_port, ZN => n37608);
   U792 : NAND4_X1 port map( A1 => n37605, A2 => n37606, A3 => n37607, A4 => 
                           n37608, ZN => n37609);
   U793 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_8_port, B1 => 
                           n37720, B2 => REGISTERS_11_8_port, ZN => n37610);
   U794 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_8_port, B1 => 
                           n37721, B2 => REGISTERS_2_8_port, ZN => n37611);
   U795 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_8_port, B1 => 
                           n37697, B2 => REGISTERS_13_8_port, C1 => n37722, C2 
                           => REGISTERS_19_8_port, ZN => n37612);
   U796 : NAND3_X1 port map( A1 => n37610, A2 => n37611, A3 => n37612, ZN => 
                           n37613);
   U797 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_8_port, B1 => 
                           n37715, B2 => REGISTERS_8_8_port, ZN => n37614);
   U798 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_8_port, B1 => 
                           n37711, B2 => REGISTERS_3_8_port, ZN => n37615);
   U799 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_8_port, B1 => 
                           n37717, B2 => REGISTERS_4_8_port, ZN => n37616);
   U800 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_8_port, B1 => 
                           n37724, B2 => REGISTERS_15_8_port, ZN => n37617);
   U801 : NAND4_X1 port map( A1 => n37614, A2 => n37615, A3 => n37616, A4 => 
                           n37617, ZN => n37618);
   U802 : OR4_X1 port map( A1 => n37604, A2 => n37609, A3 => n37613, A4 => 
                           n37618, ZN => OUTB(8));
   U803 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_3_port, B1 => 
                           n37701, B2 => REGISTERS_16_3_port, ZN => n37619);
   U804 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_3_port, B1 => 
                           n37710, B2 => REGISTERS_6_3_port, ZN => n37620);
   U805 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_3_port, B1 => 
                           n37707, B2 => REGISTERS_24_3_port, ZN => n37621);
   U806 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_3_port, B1 => 
                           n37705, B2 => REGISTERS_12_3_port, ZN => n37622);
   U807 : NAND4_X1 port map( A1 => n37619, A2 => n37620, A3 => n37621, A4 => 
                           n37622, ZN => n37623);
   U808 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_3_port, B1 => 
                           n37703, B2 => REGISTERS_1_3_port, ZN => n37624);
   U809 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_3_port, B1 => 
                           n37699, B2 => REGISTERS_20_3_port, ZN => n37625);
   U810 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_3_port, B1 => 
                           n37700, B2 => REGISTERS_18_3_port, ZN => n37626);
   U811 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_3_port, B1 => 
                           n37718, B2 => REGISTERS_28_3_port, ZN => n37627);
   U812 : NAND4_X1 port map( A1 => n37624, A2 => n37625, A3 => n37626, A4 => 
                           n37627, ZN => n37628);
   U813 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_3_port, B1 => 
                           n37720, B2 => REGISTERS_11_3_port, ZN => n37629);
   U814 : AOI22_X1 port map( A1 => n38277, A2 => REGISTERS_31_3_port, B1 => 
                           n38278, B2 => REGISTERS_2_3_port, ZN => n37630);
   U815 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_3_port, B1 => 
                           n37697, B2 => REGISTERS_13_3_port, C1 => n37722, C2 
                           => REGISTERS_19_3_port, ZN => n37631);
   U816 : NAND3_X1 port map( A1 => n37629, A2 => n37630, A3 => n37631, ZN => 
                           n37632);
   U817 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_3_port, B1 => 
                           n37715, B2 => REGISTERS_8_3_port, ZN => n37633);
   U818 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_3_port, B1 => 
                           n37711, B2 => REGISTERS_3_3_port, ZN => n37634);
   U819 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_3_port, B1 => 
                           n37717, B2 => REGISTERS_4_3_port, ZN => n37635);
   U820 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_3_port, B1 => 
                           n38289, B2 => REGISTERS_15_3_port, ZN => n37636);
   U821 : NAND4_X1 port map( A1 => n37633, A2 => n37634, A3 => n37635, A4 => 
                           n37636, ZN => n37637);
   U822 : OR4_X1 port map( A1 => n37623, A2 => n37628, A3 => n37632, A4 => 
                           n37637, ZN => OUTB(3));
   U823 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_2_port, B1 => 
                           n37701, B2 => REGISTERS_16_2_port, ZN => n37638);
   U824 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_2_port, B1 => 
                           n37710, B2 => REGISTERS_6_2_port, ZN => n37639);
   U825 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_2_port, B1 => 
                           n37707, B2 => REGISTERS_24_2_port, ZN => n37640);
   U826 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_2_port, B1 => 
                           n37705, B2 => REGISTERS_12_2_port, ZN => n37641);
   U827 : NAND4_X1 port map( A1 => n37638, A2 => n37639, A3 => n37640, A4 => 
                           n37641, ZN => n37642);
   U828 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_2_port, B1 => 
                           n37703, B2 => REGISTERS_1_2_port, ZN => n37643);
   U829 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_2_port, B1 => 
                           n37699, B2 => REGISTERS_20_2_port, ZN => n37644);
   U830 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_2_port, B1 => 
                           n37700, B2 => REGISTERS_18_2_port, ZN => n37645);
   U831 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_2_port, B1 => 
                           n37718, B2 => REGISTERS_28_2_port, ZN => n37646);
   U832 : NAND4_X1 port map( A1 => n37643, A2 => n37644, A3 => n37645, A4 => 
                           n37646, ZN => n37647);
   U833 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_2_port, B1 => 
                           n37720, B2 => REGISTERS_11_2_port, ZN => n37648);
   U834 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_2_port, B1 => 
                           n37721, B2 => REGISTERS_2_2_port, ZN => n37649);
   U835 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_2_port, B1 => 
                           n37697, B2 => REGISTERS_13_2_port, C1 => n37722, C2 
                           => REGISTERS_19_2_port, ZN => n37650);
   U836 : NAND3_X1 port map( A1 => n37648, A2 => n37649, A3 => n37650, ZN => 
                           n37651);
   U837 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_2_port, B1 => 
                           n37715, B2 => REGISTERS_8_2_port, ZN => n37652);
   U838 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_2_port, B1 => 
                           n37711, B2 => REGISTERS_3_2_port, ZN => n37653);
   U839 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_2_port, B1 => 
                           n37717, B2 => REGISTERS_4_2_port, ZN => n37654);
   U840 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_2_port, B1 => 
                           n37724, B2 => REGISTERS_15_2_port, ZN => n37655);
   U841 : NAND4_X1 port map( A1 => n37652, A2 => n37653, A3 => n37654, A4 => 
                           n37655, ZN => n37656);
   U842 : OR4_X1 port map( A1 => n37642, A2 => n37647, A3 => n37651, A4 => 
                           n37656, ZN => OUTB(2));
   U843 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_1_port, B1 => 
                           n37701, B2 => REGISTERS_16_1_port, ZN => n37657);
   U844 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_1_port, B1 => 
                           n37710, B2 => REGISTERS_6_1_port, ZN => n37658);
   U845 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_1_port, B1 => 
                           n37707, B2 => REGISTERS_24_1_port, ZN => n37659);
   U846 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_1_port, B1 => 
                           n37705, B2 => REGISTERS_12_1_port, ZN => n37660);
   U847 : NAND4_X1 port map( A1 => n37657, A2 => n37658, A3 => n37659, A4 => 
                           n37660, ZN => n37661);
   U848 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_1_port, B1 => 
                           n37703, B2 => REGISTERS_1_1_port, ZN => n37662);
   U849 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_1_port, B1 => 
                           n37699, B2 => REGISTERS_20_1_port, ZN => n37663);
   U850 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_1_port, B1 => 
                           n37700, B2 => REGISTERS_18_1_port, ZN => n37664);
   U851 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_1_port, B1 => 
                           n37718, B2 => REGISTERS_28_1_port, ZN => n37665);
   U852 : NAND4_X1 port map( A1 => n37662, A2 => n37663, A3 => n37664, A4 => 
                           n37665, ZN => n37666);
   U853 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_1_port, B1 => 
                           n37720, B2 => REGISTERS_11_1_port, ZN => n37667);
   U854 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_1_port, B1 => 
                           n37721, B2 => REGISTERS_2_1_port, ZN => n37668);
   U855 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_1_port, B1 => 
                           n37697, B2 => REGISTERS_13_1_port, C1 => n37722, C2 
                           => REGISTERS_19_1_port, ZN => n37669);
   U856 : NAND3_X1 port map( A1 => n37667, A2 => n37668, A3 => n37669, ZN => 
                           n37670);
   U857 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_1_port, B1 => 
                           n37715, B2 => REGISTERS_8_1_port, ZN => n37671);
   U858 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_1_port, B1 => 
                           n37711, B2 => REGISTERS_3_1_port, ZN => n37672);
   U859 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_1_port, B1 => 
                           n37717, B2 => REGISTERS_4_1_port, ZN => n37673);
   U860 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_1_port, B1 => 
                           n37724, B2 => REGISTERS_15_1_port, ZN => n37674);
   U861 : NAND4_X1 port map( A1 => n37671, A2 => n37672, A3 => n37673, A4 => 
                           n37674, ZN => n37675);
   U862 : OR4_X1 port map( A1 => n37661, A2 => n37666, A3 => n37670, A4 => 
                           n37675, ZN => OUTB(1));
   U863 : AOI22_X1 port map( A1 => n37702, A2 => REGISTERS_9_0_port, B1 => 
                           n37701, B2 => REGISTERS_16_0_port, ZN => n37676);
   U864 : AOI22_X1 port map( A1 => n37708, A2 => REGISTERS_23_0_port, B1 => 
                           n37710, B2 => REGISTERS_6_0_port, ZN => n37677);
   U865 : AOI22_X1 port map( A1 => n37706, A2 => REGISTERS_14_0_port, B1 => 
                           n37707, B2 => REGISTERS_24_0_port, ZN => n37678);
   U866 : AOI22_X1 port map( A1 => n37704, A2 => REGISTERS_10_0_port, B1 => 
                           n37705, B2 => REGISTERS_12_0_port, ZN => n37679);
   U867 : NAND4_X1 port map( A1 => n37676, A2 => n37677, A3 => n37678, A4 => 
                           n37679, ZN => n37680);
   U868 : AOI22_X1 port map( A1 => n37723, A2 => REGISTERS_27_0_port, B1 => 
                           n37703, B2 => REGISTERS_1_0_port, ZN => n37681);
   U869 : AOI22_X1 port map( A1 => n37695, A2 => REGISTERS_21_0_port, B1 => 
                           n37699, B2 => REGISTERS_20_0_port, ZN => n37682);
   U870 : AOI22_X1 port map( A1 => n37698, A2 => REGISTERS_7_0_port, B1 => 
                           n37700, B2 => REGISTERS_18_0_port, ZN => n37683);
   U871 : AOI22_X1 port map( A1 => n37716, A2 => REGISTERS_5_0_port, B1 => 
                           n37718, B2 => REGISTERS_28_0_port, ZN => n37684);
   U872 : NAND4_X1 port map( A1 => n37681, A2 => n37682, A3 => n37683, A4 => 
                           n37684, ZN => n37685);
   U873 : AOI22_X1 port map( A1 => n37709, A2 => REGISTERS_25_0_port, B1 => 
                           n37720, B2 => REGISTERS_11_0_port, ZN => n37686);
   U874 : AOI22_X1 port map( A1 => n37725, A2 => REGISTERS_31_0_port, B1 => 
                           n37721, B2 => REGISTERS_2_0_port, ZN => n37687);
   U875 : AOI222_X1 port map( A1 => n37696, A2 => REGISTERS_29_0_port, B1 => 
                           n37697, B2 => REGISTERS_13_0_port, C1 => n37722, C2 
                           => REGISTERS_19_0_port, ZN => n37688);
   U876 : NAND3_X1 port map( A1 => n37686, A2 => n37687, A3 => n37688, ZN => 
                           n37689);
   U877 : AOI22_X1 port map( A1 => n37712, A2 => REGISTERS_26_0_port, B1 => 
                           n37715, B2 => REGISTERS_8_0_port, ZN => n37690);
   U878 : AOI22_X1 port map( A1 => n37714, A2 => REGISTERS_30_0_port, B1 => 
                           n37711, B2 => REGISTERS_3_0_port, ZN => n37691);
   U879 : AOI22_X1 port map( A1 => n37719, A2 => REGISTERS_17_0_port, B1 => 
                           n37717, B2 => REGISTERS_4_0_port, ZN => n37692);
   U880 : AOI22_X1 port map( A1 => n37713, A2 => REGISTERS_22_0_port, B1 => 
                           n37724, B2 => REGISTERS_15_0_port, ZN => n37693);
   U881 : NAND4_X1 port map( A1 => n37690, A2 => n37691, A3 => n37692, A4 => 
                           n37693, ZN => n37694);
   U882 : OR4_X1 port map( A1 => n37680, A2 => n37685, A3 => n37689, A4 => 
                           n37694, ZN => OUTB(0));
   U883 : BUF_X2 port map( A => n38300, Z => n37695);
   U884 : BUF_X2 port map( A => n38279, Z => n37696);
   U885 : BUF_X2 port map( A => n38280, Z => n37697);
   U886 : BUF_X2 port map( A => n38302, Z => n37698);
   U887 : BUF_X2 port map( A => n38301, Z => n37699);
   U888 : BUF_X2 port map( A => n38303, Z => n37700);
   U889 : BUF_X2 port map( A => n38291, Z => n37701);
   U890 : BUF_X2 port map( A => n38290, Z => n37702);
   U891 : BUF_X2 port map( A => n38299, Z => n37703);
   U892 : BUF_X2 port map( A => n38296, Z => n37704);
   U893 : BUF_X2 port map( A => n38297, Z => n37705);
   U894 : BUF_X2 port map( A => n38294, Z => n37706);
   U895 : BUF_X2 port map( A => n38295, Z => n37707);
   U896 : BUF_X2 port map( A => n38292, Z => n37708);
   U897 : BUF_X2 port map( A => n38275, Z => n37709);
   U898 : BUF_X2 port map( A => n38293, Z => n37710);
   U899 : BUF_X2 port map( A => n38285, Z => n37711);
   U900 : BUF_X2 port map( A => n38282, Z => n37712);
   U901 : BUF_X2 port map( A => n38288, Z => n37713);
   U902 : BUF_X2 port map( A => n38284, Z => n37714);
   U903 : BUF_X2 port map( A => n38283, Z => n37715);
   U904 : BUF_X2 port map( A => n38304, Z => n37716);
   U905 : BUF_X2 port map( A => n38287, Z => n37717);
   U906 : BUF_X2 port map( A => n38305, Z => n37718);
   U907 : BUF_X2 port map( A => n38286, Z => n37719);
   U908 : BUF_X2 port map( A => n38276, Z => n37720);
   U909 : BUF_X2 port map( A => n38278, Z => n37721);
   U910 : BUF_X2 port map( A => n38281, Z => n37722);
   U911 : BUF_X2 port map( A => n38298, Z => n37723);
   U912 : BUF_X2 port map( A => n38289, Z => n37724);
   U913 : BUF_X2 port map( A => n38277, Z => n37725);
   U914 : NOR3_X2 port map( A1 => ADD_RDA(2), A2 => n37811, A3 => n37813, ZN =>
                           n38221);
   U915 : BUF_X1 port map( A => n38230, Z => n37743);
   U916 : BUF_X1 port map( A => n38221, Z => n37738);
   U917 : BUF_X1 port map( A => n38231, Z => n37744);
   U918 : BUF_X1 port map( A => n38218, Z => n37735);
   U919 : BUF_X1 port map( A => n38246, Z => n37755);
   U920 : BUF_X1 port map( A => n38243, Z => n37752);
   U921 : BUF_X1 port map( A => n38241, Z => n37750);
   U922 : BUF_X1 port map( A => n38210, Z => n37731);
   U923 : BUF_X1 port map( A => n38208, Z => n37729);
   U924 : BUF_X1 port map( A => n38206, Z => n37727);
   U925 : BUF_X1 port map( A => n38240, Z => n37749);
   U926 : BUF_X1 port map( A => n38232, Z => n37745);
   U927 : BUF_X1 port map( A => n38228, Z => n37741);
   U928 : BUF_X1 port map( A => n38211, Z => n37732);
   U929 : BUF_X1 port map( A => n38247, Z => n37756);
   U930 : BUF_X1 port map( A => n38245, Z => n37754);
   U931 : BUF_X1 port map( A => n38235, Z => n37748);
   U932 : BUF_X1 port map( A => n38233, Z => n37746);
   U933 : BUF_X1 port map( A => n38229, Z => n37742);
   U934 : BUF_X1 port map( A => n38223, Z => n37740);
   U935 : BUF_X1 port map( A => n38219, Z => n37736);
   U936 : BUF_X1 port map( A => n38217, Z => n37734);
   U937 : BUF_X1 port map( A => n38209, Z => n37730);
   U938 : BUF_X1 port map( A => n38234, Z => n37747);
   U939 : BUF_X1 port map( A => n38222, Z => n37739);
   U940 : BUF_X1 port map( A => n38244, Z => n37753);
   U941 : BUF_X1 port map( A => n38242, Z => n37751);
   U942 : BUF_X1 port map( A => n38220, Z => n37737);
   U943 : BUF_X1 port map( A => n38216, Z => n37733);
   U944 : BUF_X1 port map( A => n38207, Z => n37728);
   U945 : BUF_X1 port map( A => n38205, Z => n37726);
   U946 : INV_X1 port map( A => ADD_RDA(1), ZN => n37811);
   U947 : INV_X1 port map( A => ADD_RDA(3), ZN => n37817);
   U948 : INV_X1 port map( A => ADD_RDA(2), ZN => n37812);
   U949 : OR4_X1 port map( A1 => n38184, A2 => n38183, A3 => n38182, A4 => 
                           n38181, ZN => OUTA(6));
   U950 : OR4_X1 port map( A1 => n38144, A2 => n38143, A3 => n38142, A4 => 
                           n38141, ZN => OUTA(3));
   U951 : OR4_X1 port map( A1 => n38164, A2 => n38163, A3 => n38162, A4 => 
                           n38161, ZN => OUTA(5));
   U952 : OR4_X1 port map( A1 => n38124, A2 => n38123, A3 => n38122, A4 => 
                           n38121, ZN => OUTA(31));
   U953 : OR4_X1 port map( A1 => n38104, A2 => n38103, A3 => n38102, A4 => 
                           n38101, ZN => OUTA(30));
   U954 : OR4_X1 port map( A1 => n37924, A2 => n37923, A3 => n37922, A4 => 
                           n37921, ZN => OUTA(22));
   U955 : OR4_X1 port map( A1 => n37984, A2 => n37983, A3 => n37982, A4 => 
                           n37981, ZN => OUTA(25));
   U956 : OR4_X1 port map( A1 => n37964, A2 => n37963, A3 => n37962, A4 => 
                           n37961, ZN => OUTA(24));
   U957 : OR4_X1 port map( A1 => n37864, A2 => n37863, A3 => n37862, A4 => 
                           n37861, ZN => OUTA(19));
   U958 : OR4_X1 port map( A1 => n37884, A2 => n37883, A3 => n37882, A4 => 
                           n37881, ZN => OUTA(20));
   U959 : OR4_X1 port map( A1 => n37844, A2 => n37843, A3 => n37842, A4 => 
                           n37841, ZN => OUTA(18));
   U960 : OR4_X1 port map( A1 => n37944, A2 => n37943, A3 => n37942, A4 => 
                           n37941, ZN => OUTA(23));
   U961 : OR4_X1 port map( A1 => n37904, A2 => n37903, A3 => n37902, A4 => 
                           n37901, ZN => OUTA(21));
   U962 : OR4_X1 port map( A1 => n38024, A2 => n38023, A3 => n38022, A4 => 
                           n38021, ZN => OUTA(27));
   U963 : OR4_X1 port map( A1 => n38204, A2 => n38203, A3 => n38202, A4 => 
                           n38201, ZN => OUTA(8));
   U964 : OR4_X1 port map( A1 => n38084, A2 => n38083, A3 => n38082, A4 => 
                           n38081, ZN => OUTA(2));
   U965 : OR4_X1 port map( A1 => n38064, A2 => n38063, A3 => n38062, A4 => 
                           n38061, ZN => OUTA(29));
   U966 : OR4_X1 port map( A1 => n38004, A2 => n38003, A3 => n38002, A4 => 
                           n38001, ZN => OUTA(26));
   U967 : OR4_X1 port map( A1 => n38255, A2 => n38254, A3 => n38253, A4 => 
                           n38252, ZN => OUTA(9));
   U968 : OR4_X1 port map( A1 => n38044, A2 => n38043, A3 => n38042, A4 => 
                           n38041, ZN => OUTA(28));
   U969 : NOR2_X1 port map( A1 => n37809, A2 => n37818, ZN => n38211);
   U970 : BUF_X1 port map( A => N291, Z => n37771);
   U971 : BUF_X1 port map( A => N290, Z => n37772);
   U972 : BUF_X1 port map( A => N292, Z => n37770);
   U973 : BUF_X1 port map( A => N293, Z => n37769);
   U974 : BUF_X1 port map( A => N294, Z => n37768);
   U975 : BUF_X1 port map( A => N285, Z => n37777);
   U976 : BUF_X1 port map( A => N284, Z => n37778);
   U977 : BUF_X1 port map( A => N286, Z => n37776);
   U978 : BUF_X1 port map( A => N287, Z => n37775);
   U979 : BUF_X1 port map( A => N288, Z => n37774);
   U980 : BUF_X1 port map( A => N289, Z => n37773);
   U981 : BUF_X1 port map( A => N302, Z => n37760);
   U982 : BUF_X1 port map( A => N303, Z => n37759);
   U983 : BUF_X1 port map( A => N304, Z => n37758);
   U984 : BUF_X1 port map( A => N305, Z => n37757);
   U985 : BUF_X1 port map( A => N295, Z => n37767);
   U986 : BUF_X1 port map( A => N296, Z => n37766);
   U987 : BUF_X1 port map( A => N297, Z => n37765);
   U988 : BUF_X1 port map( A => N298, Z => n37764);
   U989 : BUF_X1 port map( A => N299, Z => n37763);
   U990 : BUF_X1 port map( A => N300, Z => n37762);
   U991 : BUF_X1 port map( A => N301, Z => n37761);
   U992 : BUF_X1 port map( A => N281, Z => n37781);
   U993 : BUF_X1 port map( A => N279, Z => n37783);
   U994 : BUF_X1 port map( A => N243, Z => n37787);
   U995 : BUF_X1 port map( A => N280, Z => n37782);
   U996 : BUF_X1 port map( A => N278, Z => n37784);
   U997 : BUF_X1 port map( A => N283, Z => n37779);
   U998 : BUF_X1 port map( A => N276, Z => n37786);
   U999 : BUF_X1 port map( A => N282, Z => n37780);
   U1000 : INV_X1 port map( A => ADD_WR(0), ZN => n37790);
   U1001 : BUF_X1 port map( A => N277, Z => n37785);
   U1002 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(0), ZN => N244);
   U1003 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(31), ZN => N275);
   U1004 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(1), ZN => N245);
   U1005 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(30), ZN => N274);
   U1006 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(29), ZN => N273);
   U1007 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(2), ZN => N246);
   U1008 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(28), ZN => N272);
   U1009 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(27), ZN => N271);
   U1010 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(3), ZN => N247);
   U1011 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(26), ZN => N270);
   U1012 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(25), ZN => N269);
   U1013 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(4), ZN => N248);
   U1014 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(24), ZN => N268);
   U1015 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(23), ZN => N267);
   U1016 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(5), ZN => N249);
   U1017 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(22), ZN => N266);
   U1018 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(21), ZN => N265);
   U1019 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(6), ZN => N250);
   U1020 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(20), ZN => N264);
   U1021 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(19), ZN => N263);
   U1022 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(7), ZN => N251);
   U1023 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(18), ZN => N262);
   U1024 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(17), ZN => N261);
   U1025 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(8), ZN => N252);
   U1026 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(15), ZN => N259);
   U1027 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(9), ZN => N253);
   U1028 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(16), ZN => N260);
   U1029 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(14), ZN => N258);
   U1030 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(10), ZN => N254);
   U1031 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(13), ZN => N257);
   U1032 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(11), ZN => N255);
   U1033 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(12), ZN => N256);
   U1034 : NOR2_X1 port map( A1 => n38262, A2 => n38271, ZN => n38289);
   U1035 : NOR2_X1 port map( A1 => n38267, A2 => n38271, ZN => n38277);
   U1036 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => ADD_WR(2)
                           , ZN => n37798);
   U1037 : NAND3_X1 port map( A1 => WE, A2 => ADD_WR(3), A3 => ADD_WR(4), ZN =>
                           n37792);
   U1038 : OAI21_X1 port map( B1 => n37798, B2 => n37792, A => RESET, ZN => 
                           N243);
   U1039 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n37790, 
                           ZN => n37799);
   U1040 : OAI21_X1 port map( B1 => n37792, B2 => n37799, A => RESET, ZN => 
                           N276);
   U1041 : INV_X1 port map( A => ADD_WR(1), ZN => n37788);
   U1042 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n37788, 
                           ZN => n37800);
   U1043 : OAI21_X1 port map( B1 => n37792, B2 => n37800, A => RESET, ZN => 
                           N277);
   U1044 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n37790, A3 => n37788, ZN 
                           => n37801);
   U1045 : OAI21_X1 port map( B1 => n37792, B2 => n37801, A => RESET, ZN => 
                           N278);
   U1046 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n37788, ZN => n37789);
   U1047 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n37789, ZN => n37802);
   U1048 : OAI21_X1 port map( B1 => n37792, B2 => n37802, A => RESET, ZN => 
                           N279);
   U1049 : NAND2_X1 port map( A1 => n37789, A2 => n37790, ZN => n37803);
   U1050 : OAI21_X1 port map( B1 => n37792, B2 => n37803, A => RESET, ZN => 
                           N280);
   U1051 : NOR2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), ZN => n37791);
   U1052 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n37791, ZN => n37805);
   U1053 : OAI21_X1 port map( B1 => n37792, B2 => n37805, A => RESET, ZN => 
                           N281);
   U1054 : NAND2_X1 port map( A1 => n37791, A2 => n37790, ZN => n37795);
   U1055 : OAI21_X1 port map( B1 => n37792, B2 => n37795, A => RESET, ZN => 
                           N282);
   U1056 : INV_X1 port map( A => ADD_WR(3), ZN => n37797);
   U1057 : NAND3_X1 port map( A1 => WE, A2 => ADD_WR(4), A3 => n37797, ZN => 
                           n37793);
   U1058 : OAI21_X1 port map( B1 => n37798, B2 => n37793, A => RESET, ZN => 
                           N283);
   U1059 : OAI21_X1 port map( B1 => n37799, B2 => n37793, A => RESET, ZN => 
                           N284);
   U1060 : OAI21_X1 port map( B1 => n37800, B2 => n37793, A => RESET, ZN => 
                           N285);
   U1061 : OAI21_X1 port map( B1 => n37801, B2 => n37793, A => RESET, ZN => 
                           N286);
   U1062 : OAI21_X1 port map( B1 => n37802, B2 => n37793, A => RESET, ZN => 
                           N287);
   U1063 : OAI21_X1 port map( B1 => n37803, B2 => n37793, A => RESET, ZN => 
                           N288);
   U1064 : OAI21_X1 port map( B1 => n37805, B2 => n37793, A => RESET, ZN => 
                           N289);
   U1065 : OAI21_X1 port map( B1 => n37795, B2 => n37793, A => RESET, ZN => 
                           N290);
   U1066 : INV_X1 port map( A => ADD_WR(4), ZN => n37796);
   U1067 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => WE, A3 => n37796, ZN => 
                           n37794);
   U1068 : OAI21_X1 port map( B1 => n37798, B2 => n37794, A => RESET, ZN => 
                           N291);
   U1069 : OAI21_X1 port map( B1 => n37799, B2 => n37794, A => RESET, ZN => 
                           N292);
   U1070 : OAI21_X1 port map( B1 => n37800, B2 => n37794, A => RESET, ZN => 
                           N293);
   U1071 : OAI21_X1 port map( B1 => n37801, B2 => n37794, A => RESET, ZN => 
                           N294);
   U1072 : OAI21_X1 port map( B1 => n37802, B2 => n37794, A => RESET, ZN => 
                           N295);
   U1073 : OAI21_X1 port map( B1 => n37803, B2 => n37794, A => RESET, ZN => 
                           N296);
   U1074 : OAI21_X1 port map( B1 => n37805, B2 => n37794, A => RESET, ZN => 
                           N297);
   U1075 : OAI21_X1 port map( B1 => n37795, B2 => n37794, A => RESET, ZN => 
                           N298);
   U1076 : NAND3_X1 port map( A1 => WE, A2 => n37797, A3 => n37796, ZN => 
                           n37804);
   U1077 : OAI21_X1 port map( B1 => n37798, B2 => n37804, A => RESET, ZN => 
                           N299);
   U1078 : OAI21_X1 port map( B1 => n37799, B2 => n37804, A => RESET, ZN => 
                           N300);
   U1079 : OAI21_X1 port map( B1 => n37800, B2 => n37804, A => RESET, ZN => 
                           N301);
   U1080 : OAI21_X1 port map( B1 => n37801, B2 => n37804, A => RESET, ZN => 
                           N302);
   U1081 : OAI21_X1 port map( B1 => n37802, B2 => n37804, A => RESET, ZN => 
                           N303);
   U1082 : OAI21_X1 port map( B1 => n37803, B2 => n37804, A => RESET, ZN => 
                           N304);
   U1083 : OAI21_X1 port map( B1 => n37805, B2 => n37804, A => RESET, ZN => 
                           N305);
   U1084 : INV_X1 port map( A => ADD_RDA(4), ZN => n37806);
   U1085 : NAND3_X1 port map( A1 => ADD_RDA(3), A2 => ADD_RDA(0), A3 => n37806,
                           ZN => n37809);
   U1086 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDA(1), A3 => n37812, ZN 
                           => n37824);
   U1087 : NOR2_X1 port map( A1 => n37809, A2 => n37824, ZN => n38206);
   U1088 : INV_X1 port map( A => ADD_RDA(0), ZN => n37807);
   U1089 : NAND3_X1 port map( A1 => ADD_RDA(4), A2 => n37817, A3 => n37807, ZN 
                           => n37808);
   U1090 : NAND3_X1 port map( A1 => RESET, A2 => n37812, A3 => n37811, ZN => 
                           n37820);
   U1091 : NOR2_X1 port map( A1 => n37808, A2 => n37820, ZN => n38205);
   U1092 : NAND3_X1 port map( A1 => ADD_RDA(0), A2 => n37817, A3 => n37806, ZN 
                           => n37816);
   U1093 : NOR2_X1 port map( A1 => n37820, A2 => n37816, ZN => n38208);
   U1094 : NAND3_X1 port map( A1 => ADD_RDA(4), A2 => ADD_RDA(3), A3 => n37807,
                           ZN => n37815);
   U1095 : NOR2_X1 port map( A1 => n37820, A2 => n37815, ZN => n38207);
   U1096 : NAND3_X1 port map( A1 => ADD_RDA(2), A2 => RESET, A3 => n37811, ZN 
                           => n37818);
   U1097 : NOR2_X1 port map( A1 => ADD_RDA(4), A2 => ADD_RDA(0), ZN => n37810);
   U1098 : NAND2_X1 port map( A1 => ADD_RDA(3), A2 => n37810, ZN => n37822);
   U1099 : NOR2_X1 port map( A1 => n37818, A2 => n37822, ZN => n38210);
   U1100 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDA(2), A3 => ADD_RDA(1), 
                           ZN => n37821);
   U1101 : NOR2_X1 port map( A1 => n37809, A2 => n37821, ZN => n38209);
   U1102 : NOR2_X1 port map( A1 => n37818, A2 => n37808, ZN => n38217);
   U1103 : NOR2_X1 port map( A1 => n37808, A2 => n37821, ZN => n38216);
   U1104 : NOR2_X1 port map( A1 => n37824, A2 => n37808, ZN => n38219);
   U1105 : NOR2_X1 port map( A1 => n37809, A2 => n37820, ZN => n38218);
   U1106 : NAND3_X1 port map( A1 => RESET, A2 => n37810, A3 => n37817, ZN => 
                           n37813);
   U1107 : NAND3_X1 port map( A1 => ADD_RDA(3), A2 => ADD_RDA(4), A3 => 
                           ADD_RDA(0), ZN => n37819);
   U1108 : NOR2_X1 port map( A1 => n37821, A2 => n37819, ZN => n38220);
   U1109 : NOR2_X1 port map( A1 => n37824, A2 => n37816, ZN => n38223);
   U1110 : NOR2_X1 port map( A1 => n37820, A2 => n37822, ZN => n38222);
   U1111 : NOR2_X1 port map( A1 => n37815, A2 => n37821, ZN => n38229);
   U1112 : NOR2_X1 port map( A1 => n37818, A2 => n37819, ZN => n38228);
   U1113 : NOR2_X1 port map( A1 => n37824, A2 => n37819, ZN => n38231);
   U1114 : NOR3_X1 port map( A1 => ADD_RDA(1), A2 => n37812, A3 => n37813, ZN 
                           => n38230);
   U1115 : NOR2_X1 port map( A1 => n37824, A2 => n37822, ZN => n38233);
   U1116 : NOR2_X1 port map( A1 => n37818, A2 => n37815, ZN => n38232);
   U1117 : NAND2_X1 port map( A1 => ADD_RDA(2), A2 => ADD_RDA(1), ZN => n37814)
                           ;
   U1118 : NOR2_X1 port map( A1 => n37814, A2 => n37813, ZN => n38235);
   U1119 : NOR2_X1 port map( A1 => n37816, A2 => n37821, ZN => n38234);
   U1120 : NOR2_X1 port map( A1 => n37824, A2 => n37815, ZN => n38241);
   U1121 : NOR2_X1 port map( A1 => n37818, A2 => n37816, ZN => n38240);
   U1122 : NAND3_X1 port map( A1 => ADD_RDA(4), A2 => ADD_RDA(0), A3 => n37817,
                           ZN => n37823);
   U1123 : NOR2_X1 port map( A1 => n37818, A2 => n37823, ZN => n38243);
   U1124 : NOR2_X1 port map( A1 => n37820, A2 => n37819, ZN => n38242);
   U1125 : NOR2_X1 port map( A1 => n37821, A2 => n37823, ZN => n38245);
   U1126 : NOR2_X1 port map( A1 => n37820, A2 => n37823, ZN => n38244);
   U1127 : NOR2_X1 port map( A1 => n37822, A2 => n37821, ZN => n38247);
   U1128 : NOR2_X1 port map( A1 => n37824, A2 => n37823, ZN => n38246);
   U1129 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_18_port, B1 => 
                           n37726, B2 => REGISTERS_16_18_port, ZN => n37828);
   U1130 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_18_port, B1 => 
                           n37728, B2 => REGISTERS_24_18_port, ZN => n37827);
   U1131 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_18_port, B1 => 
                           n37730, B2 => REGISTERS_15_18_port, ZN => n37826);
   U1132 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_18_port, ZN => 
                           n37825);
   U1133 : NAND4_X1 port map( A1 => n37828, A2 => n37827, A3 => n37826, A4 => 
                           n37825, ZN => n37844);
   U1134 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_18_port, B1 => 
                           n37733, B2 => REGISTERS_22_18_port, ZN => n37832);
   U1135 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_18_port, B1 => 
                           n37735, B2 => REGISTERS_9_18_port, ZN => n37831);
   U1136 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_18_port, B1 => 
                           n37737, B2 => REGISTERS_31_18_port, ZN => n37830);
   U1137 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_18_port, B1 => 
                           n37739, B2 => REGISTERS_8_18_port, ZN => n37829);
   U1138 : NAND4_X1 port map( A1 => n37832, A2 => n37831, A3 => n37830, A4 => 
                           n37829, ZN => n37843);
   U1139 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_18_port, B1 => 
                           n37741, B2 => REGISTERS_29_18_port, ZN => n37836);
   U1140 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_18_port, B1 => 
                           n37743, B2 => REGISTERS_4_18_port, ZN => n37835);
   U1141 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_18_port, B1 => 
                           n37745, B2 => REGISTERS_28_18_port, ZN => n37834);
   U1142 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_18_port, B1 => 
                           n37747, B2 => REGISTERS_7_18_port, ZN => n37833);
   U1143 : NAND4_X1 port map( A1 => n37836, A2 => n37835, A3 => n37834, A4 => 
                           n37833, ZN => n37842);
   U1144 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_18_port, B1 => 
                           n37749, B2 => REGISTERS_5_18_port, ZN => n37840);
   U1145 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_18_port, B1 => 
                           n37751, B2 => REGISTERS_25_18_port, ZN => n37839);
   U1146 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_18_port, B1 => 
                           n37753, B2 => REGISTERS_17_18_port, ZN => n37838);
   U1147 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_18_port, B1 => 
                           n37755, B2 => REGISTERS_19_18_port, ZN => n37837);
   U1148 : NAND4_X1 port map( A1 => n37840, A2 => n37839, A3 => n37838, A4 => 
                           n37837, ZN => n37841);
   U1149 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_19_port, B1 => 
                           n37726, B2 => REGISTERS_16_19_port, ZN => n37848);
   U1150 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_19_port, B1 => 
                           n37728, B2 => REGISTERS_24_19_port, ZN => n37847);
   U1151 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_19_port, B1 => 
                           n37730, B2 => REGISTERS_15_19_port, ZN => n37846);
   U1152 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_19_port, ZN => 
                           n37845);
   U1153 : NAND4_X1 port map( A1 => n37848, A2 => n37847, A3 => n37846, A4 => 
                           n37845, ZN => n37864);
   U1154 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_19_port, B1 => 
                           n37733, B2 => REGISTERS_22_19_port, ZN => n37852);
   U1155 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_19_port, B1 => 
                           n37735, B2 => REGISTERS_9_19_port, ZN => n37851);
   U1156 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_19_port, B1 => 
                           n37737, B2 => REGISTERS_31_19_port, ZN => n37850);
   U1157 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_19_port, B1 => 
                           n37739, B2 => REGISTERS_8_19_port, ZN => n37849);
   U1158 : NAND4_X1 port map( A1 => n37852, A2 => n37851, A3 => n37850, A4 => 
                           n37849, ZN => n37863);
   U1159 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_19_port, B1 => 
                           n37741, B2 => REGISTERS_29_19_port, ZN => n37856);
   U1160 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_19_port, B1 => 
                           n37743, B2 => REGISTERS_4_19_port, ZN => n37855);
   U1161 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_19_port, B1 => 
                           n37745, B2 => REGISTERS_28_19_port, ZN => n37854);
   U1162 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_19_port, B1 => 
                           n37747, B2 => REGISTERS_7_19_port, ZN => n37853);
   U1163 : NAND4_X1 port map( A1 => n37856, A2 => n37855, A3 => n37854, A4 => 
                           n37853, ZN => n37862);
   U1164 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_19_port, B1 => 
                           n37749, B2 => REGISTERS_5_19_port, ZN => n37860);
   U1165 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_19_port, B1 => 
                           n37751, B2 => REGISTERS_25_19_port, ZN => n37859);
   U1166 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_19_port, B1 => 
                           n37753, B2 => REGISTERS_17_19_port, ZN => n37858);
   U1167 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_19_port, B1 => 
                           n37755, B2 => REGISTERS_19_19_port, ZN => n37857);
   U1168 : NAND4_X1 port map( A1 => n37860, A2 => n37859, A3 => n37858, A4 => 
                           n37857, ZN => n37861);
   U1169 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_20_port, B1 => 
                           n37726, B2 => REGISTERS_16_20_port, ZN => n37868);
   U1170 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_20_port, B1 => 
                           n37728, B2 => REGISTERS_24_20_port, ZN => n37867);
   U1171 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_20_port, B1 => 
                           n37730, B2 => REGISTERS_15_20_port, ZN => n37866);
   U1172 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_20_port, ZN => 
                           n37865);
   U1173 : NAND4_X1 port map( A1 => n37868, A2 => n37867, A3 => n37866, A4 => 
                           n37865, ZN => n37884);
   U1174 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_20_port, B1 => 
                           n37733, B2 => REGISTERS_22_20_port, ZN => n37872);
   U1175 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_20_port, B1 => 
                           n37735, B2 => REGISTERS_9_20_port, ZN => n37871);
   U1176 : AOI22_X1 port map( A1 => n38221, A2 => REGISTERS_2_20_port, B1 => 
                           n37737, B2 => REGISTERS_31_20_port, ZN => n37870);
   U1177 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_20_port, B1 => 
                           n37739, B2 => REGISTERS_8_20_port, ZN => n37869);
   U1178 : NAND4_X1 port map( A1 => n37872, A2 => n37871, A3 => n37870, A4 => 
                           n37869, ZN => n37883);
   U1179 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_20_port, B1 => 
                           n37741, B2 => REGISTERS_29_20_port, ZN => n37876);
   U1180 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_20_port, B1 => 
                           n37743, B2 => REGISTERS_4_20_port, ZN => n37875);
   U1181 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_20_port, B1 => 
                           n37745, B2 => REGISTERS_28_20_port, ZN => n37874);
   U1182 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_20_port, B1 => 
                           n37747, B2 => REGISTERS_7_20_port, ZN => n37873);
   U1183 : NAND4_X1 port map( A1 => n37876, A2 => n37875, A3 => n37874, A4 => 
                           n37873, ZN => n37882);
   U1184 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_20_port, B1 => 
                           n37749, B2 => REGISTERS_5_20_port, ZN => n37880);
   U1185 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_20_port, B1 => 
                           n37751, B2 => REGISTERS_25_20_port, ZN => n37879);
   U1186 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_20_port, B1 => 
                           n37753, B2 => REGISTERS_17_20_port, ZN => n37878);
   U1187 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_20_port, B1 => 
                           n37755, B2 => REGISTERS_19_20_port, ZN => n37877);
   U1188 : NAND4_X1 port map( A1 => n37880, A2 => n37879, A3 => n37878, A4 => 
                           n37877, ZN => n37881);
   U1189 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_21_port, B1 => 
                           n37726, B2 => REGISTERS_16_21_port, ZN => n37888);
   U1190 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_21_port, B1 => 
                           n37728, B2 => REGISTERS_24_21_port, ZN => n37887);
   U1191 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_21_port, B1 => 
                           n37730, B2 => REGISTERS_15_21_port, ZN => n37886);
   U1192 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_21_port, ZN => 
                           n37885);
   U1193 : NAND4_X1 port map( A1 => n37888, A2 => n37887, A3 => n37886, A4 => 
                           n37885, ZN => n37904);
   U1194 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_21_port, B1 => 
                           n37733, B2 => REGISTERS_22_21_port, ZN => n37892);
   U1195 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_21_port, B1 => 
                           n37735, B2 => REGISTERS_9_21_port, ZN => n37891);
   U1196 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_21_port, B1 => 
                           n37737, B2 => REGISTERS_31_21_port, ZN => n37890);
   U1197 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_21_port, B1 => 
                           n37739, B2 => REGISTERS_8_21_port, ZN => n37889);
   U1198 : NAND4_X1 port map( A1 => n37892, A2 => n37891, A3 => n37890, A4 => 
                           n37889, ZN => n37903);
   U1199 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_21_port, B1 => 
                           n37741, B2 => REGISTERS_29_21_port, ZN => n37896);
   U1200 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_21_port, B1 => 
                           n37743, B2 => REGISTERS_4_21_port, ZN => n37895);
   U1201 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_21_port, B1 => 
                           n37745, B2 => REGISTERS_28_21_port, ZN => n37894);
   U1202 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_21_port, B1 => 
                           n37747, B2 => REGISTERS_7_21_port, ZN => n37893);
   U1203 : NAND4_X1 port map( A1 => n37896, A2 => n37895, A3 => n37894, A4 => 
                           n37893, ZN => n37902);
   U1204 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_21_port, B1 => 
                           n37749, B2 => REGISTERS_5_21_port, ZN => n37900);
   U1205 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_21_port, B1 => 
                           n37751, B2 => REGISTERS_25_21_port, ZN => n37899);
   U1206 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_21_port, B1 => 
                           n37753, B2 => REGISTERS_17_21_port, ZN => n37898);
   U1207 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_21_port, B1 => 
                           n37755, B2 => REGISTERS_19_21_port, ZN => n37897);
   U1208 : NAND4_X1 port map( A1 => n37900, A2 => n37899, A3 => n37898, A4 => 
                           n37897, ZN => n37901);
   U1209 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_22_port, B1 => 
                           n37726, B2 => REGISTERS_16_22_port, ZN => n37908);
   U1210 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_22_port, B1 => 
                           n37728, B2 => REGISTERS_24_22_port, ZN => n37907);
   U1211 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_22_port, B1 => 
                           n37730, B2 => REGISTERS_15_22_port, ZN => n37906);
   U1212 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_22_port, ZN => 
                           n37905);
   U1213 : NAND4_X1 port map( A1 => n37908, A2 => n37907, A3 => n37906, A4 => 
                           n37905, ZN => n37924);
   U1214 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_22_port, B1 => 
                           n37733, B2 => REGISTERS_22_22_port, ZN => n37912);
   U1215 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_22_port, B1 => 
                           n37735, B2 => REGISTERS_9_22_port, ZN => n37911);
   U1216 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_22_port, B1 => 
                           n37737, B2 => REGISTERS_31_22_port, ZN => n37910);
   U1217 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_22_port, B1 => 
                           n37739, B2 => REGISTERS_8_22_port, ZN => n37909);
   U1218 : NAND4_X1 port map( A1 => n37912, A2 => n37911, A3 => n37910, A4 => 
                           n37909, ZN => n37923);
   U1219 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_22_port, B1 => 
                           n37741, B2 => REGISTERS_29_22_port, ZN => n37916);
   U1220 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_22_port, B1 => 
                           n37743, B2 => REGISTERS_4_22_port, ZN => n37915);
   U1221 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_22_port, B1 => 
                           n37745, B2 => REGISTERS_28_22_port, ZN => n37914);
   U1222 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_22_port, B1 => 
                           n37747, B2 => REGISTERS_7_22_port, ZN => n37913);
   U1223 : NAND4_X1 port map( A1 => n37916, A2 => n37915, A3 => n37914, A4 => 
                           n37913, ZN => n37922);
   U1224 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_22_port, B1 => 
                           n37749, B2 => REGISTERS_5_22_port, ZN => n37920);
   U1225 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_22_port, B1 => 
                           n37751, B2 => REGISTERS_25_22_port, ZN => n37919);
   U1226 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_22_port, B1 => 
                           n37753, B2 => REGISTERS_17_22_port, ZN => n37918);
   U1227 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_22_port, B1 => 
                           n37755, B2 => REGISTERS_19_22_port, ZN => n37917);
   U1228 : NAND4_X1 port map( A1 => n37920, A2 => n37919, A3 => n37918, A4 => 
                           n37917, ZN => n37921);
   U1229 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_23_port, B1 => 
                           n37726, B2 => REGISTERS_16_23_port, ZN => n37928);
   U1230 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_23_port, B1 => 
                           n37728, B2 => REGISTERS_24_23_port, ZN => n37927);
   U1231 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_23_port, B1 => 
                           n37730, B2 => REGISTERS_15_23_port, ZN => n37926);
   U1232 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_23_port, ZN => 
                           n37925);
   U1233 : NAND4_X1 port map( A1 => n37928, A2 => n37927, A3 => n37926, A4 => 
                           n37925, ZN => n37944);
   U1234 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_23_port, B1 => 
                           n37733, B2 => REGISTERS_22_23_port, ZN => n37932);
   U1235 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_23_port, B1 => 
                           n37735, B2 => REGISTERS_9_23_port, ZN => n37931);
   U1236 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_23_port, B1 => 
                           n37737, B2 => REGISTERS_31_23_port, ZN => n37930);
   U1237 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_23_port, B1 => 
                           n37739, B2 => REGISTERS_8_23_port, ZN => n37929);
   U1238 : NAND4_X1 port map( A1 => n37932, A2 => n37931, A3 => n37930, A4 => 
                           n37929, ZN => n37943);
   U1239 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_23_port, B1 => 
                           n37741, B2 => REGISTERS_29_23_port, ZN => n37936);
   U1240 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_23_port, B1 => 
                           n37743, B2 => REGISTERS_4_23_port, ZN => n37935);
   U1241 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_23_port, B1 => 
                           n37745, B2 => REGISTERS_28_23_port, ZN => n37934);
   U1242 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_23_port, B1 => 
                           n37747, B2 => REGISTERS_7_23_port, ZN => n37933);
   U1243 : NAND4_X1 port map( A1 => n37936, A2 => n37935, A3 => n37934, A4 => 
                           n37933, ZN => n37942);
   U1244 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_23_port, B1 => 
                           n37749, B2 => REGISTERS_5_23_port, ZN => n37940);
   U1245 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_23_port, B1 => 
                           n37751, B2 => REGISTERS_25_23_port, ZN => n37939);
   U1246 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_23_port, B1 => 
                           n37753, B2 => REGISTERS_17_23_port, ZN => n37938);
   U1247 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_23_port, B1 => 
                           n37755, B2 => REGISTERS_19_23_port, ZN => n37937);
   U1248 : NAND4_X1 port map( A1 => n37940, A2 => n37939, A3 => n37938, A4 => 
                           n37937, ZN => n37941);
   U1249 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_24_port, B1 => 
                           n37726, B2 => REGISTERS_16_24_port, ZN => n37948);
   U1250 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_24_port, B1 => 
                           n37728, B2 => REGISTERS_24_24_port, ZN => n37947);
   U1251 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_24_port, B1 => 
                           n37730, B2 => REGISTERS_15_24_port, ZN => n37946);
   U1252 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_24_port, ZN => 
                           n37945);
   U1253 : NAND4_X1 port map( A1 => n37948, A2 => n37947, A3 => n37946, A4 => 
                           n37945, ZN => n37964);
   U1254 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_24_port, B1 => 
                           n37733, B2 => REGISTERS_22_24_port, ZN => n37952);
   U1255 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_24_port, B1 => 
                           n37735, B2 => REGISTERS_9_24_port, ZN => n37951);
   U1256 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_24_port, B1 => 
                           n37737, B2 => REGISTERS_31_24_port, ZN => n37950);
   U1257 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_24_port, B1 => 
                           n37739, B2 => REGISTERS_8_24_port, ZN => n37949);
   U1258 : NAND4_X1 port map( A1 => n37952, A2 => n37951, A3 => n37950, A4 => 
                           n37949, ZN => n37963);
   U1259 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_24_port, B1 => 
                           n37741, B2 => REGISTERS_29_24_port, ZN => n37956);
   U1260 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_24_port, B1 => 
                           n37743, B2 => REGISTERS_4_24_port, ZN => n37955);
   U1261 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_24_port, B1 => 
                           n37745, B2 => REGISTERS_28_24_port, ZN => n37954);
   U1262 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_24_port, B1 => 
                           n37747, B2 => REGISTERS_7_24_port, ZN => n37953);
   U1263 : NAND4_X1 port map( A1 => n37956, A2 => n37955, A3 => n37954, A4 => 
                           n37953, ZN => n37962);
   U1264 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_24_port, B1 => 
                           n37749, B2 => REGISTERS_5_24_port, ZN => n37960);
   U1265 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_24_port, B1 => 
                           n37751, B2 => REGISTERS_25_24_port, ZN => n37959);
   U1266 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_24_port, B1 => 
                           n37753, B2 => REGISTERS_17_24_port, ZN => n37958);
   U1267 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_24_port, B1 => 
                           n37755, B2 => REGISTERS_19_24_port, ZN => n37957);
   U1268 : NAND4_X1 port map( A1 => n37960, A2 => n37959, A3 => n37958, A4 => 
                           n37957, ZN => n37961);
   U1269 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_25_port, B1 => 
                           n37726, B2 => REGISTERS_16_25_port, ZN => n37968);
   U1270 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_25_port, B1 => 
                           n37728, B2 => REGISTERS_24_25_port, ZN => n37967);
   U1271 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_25_port, B1 => 
                           n37730, B2 => REGISTERS_15_25_port, ZN => n37966);
   U1272 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_25_port, ZN => 
                           n37965);
   U1273 : NAND4_X1 port map( A1 => n37968, A2 => n37967, A3 => n37966, A4 => 
                           n37965, ZN => n37984);
   U1274 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_25_port, B1 => 
                           n37733, B2 => REGISTERS_22_25_port, ZN => n37972);
   U1275 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_25_port, B1 => 
                           n37735, B2 => REGISTERS_9_25_port, ZN => n37971);
   U1276 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_25_port, B1 => 
                           n37737, B2 => REGISTERS_31_25_port, ZN => n37970);
   U1277 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_25_port, B1 => 
                           n37739, B2 => REGISTERS_8_25_port, ZN => n37969);
   U1278 : NAND4_X1 port map( A1 => n37972, A2 => n37971, A3 => n37970, A4 => 
                           n37969, ZN => n37983);
   U1279 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_25_port, B1 => 
                           n37741, B2 => REGISTERS_29_25_port, ZN => n37976);
   U1280 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_25_port, B1 => 
                           n37743, B2 => REGISTERS_4_25_port, ZN => n37975);
   U1281 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_25_port, B1 => 
                           n37745, B2 => REGISTERS_28_25_port, ZN => n37974);
   U1282 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_25_port, B1 => 
                           n37747, B2 => REGISTERS_7_25_port, ZN => n37973);
   U1283 : NAND4_X1 port map( A1 => n37976, A2 => n37975, A3 => n37974, A4 => 
                           n37973, ZN => n37982);
   U1284 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_25_port, B1 => 
                           n37749, B2 => REGISTERS_5_25_port, ZN => n37980);
   U1285 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_25_port, B1 => 
                           n37751, B2 => REGISTERS_25_25_port, ZN => n37979);
   U1286 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_25_port, B1 => 
                           n37753, B2 => REGISTERS_17_25_port, ZN => n37978);
   U1287 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_25_port, B1 => 
                           n37755, B2 => REGISTERS_19_25_port, ZN => n37977);
   U1288 : NAND4_X1 port map( A1 => n37980, A2 => n37979, A3 => n37978, A4 => 
                           n37977, ZN => n37981);
   U1289 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_26_port, B1 => 
                           n38205, B2 => REGISTERS_16_26_port, ZN => n37988);
   U1290 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_26_port, B1 => 
                           n38207, B2 => REGISTERS_24_26_port, ZN => n37987);
   U1291 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_26_port, B1 => 
                           n38209, B2 => REGISTERS_15_26_port, ZN => n37986);
   U1292 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_26_port, ZN => 
                           n37985);
   U1293 : NAND4_X1 port map( A1 => n37988, A2 => n37987, A3 => n37986, A4 => 
                           n37985, ZN => n38004);
   U1294 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_26_port, B1 => 
                           n38216, B2 => REGISTERS_22_26_port, ZN => n37992);
   U1295 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_26_port, B1 => 
                           n38218, B2 => REGISTERS_9_26_port, ZN => n37991);
   U1296 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_26_port, B1 => 
                           n38220, B2 => REGISTERS_31_26_port, ZN => n37990);
   U1297 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_26_port, B1 => 
                           n38222, B2 => REGISTERS_8_26_port, ZN => n37989);
   U1298 : NAND4_X1 port map( A1 => n37992, A2 => n37991, A3 => n37990, A4 => 
                           n37989, ZN => n38003);
   U1299 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_26_port, B1 => 
                           n38228, B2 => REGISTERS_29_26_port, ZN => n37996);
   U1300 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_26_port, B1 => 
                           n37743, B2 => REGISTERS_4_26_port, ZN => n37995);
   U1301 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_26_port, B1 => 
                           n38232, B2 => REGISTERS_28_26_port, ZN => n37994);
   U1302 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_26_port, B1 => 
                           n38234, B2 => REGISTERS_7_26_port, ZN => n37993);
   U1303 : NAND4_X1 port map( A1 => n37996, A2 => n37995, A3 => n37994, A4 => 
                           n37993, ZN => n38002);
   U1304 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_26_port, B1 => 
                           n38240, B2 => REGISTERS_5_26_port, ZN => n38000);
   U1305 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_26_port, B1 => 
                           n37751, B2 => REGISTERS_25_26_port, ZN => n37999);
   U1306 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_26_port, B1 => 
                           n37753, B2 => REGISTERS_17_26_port, ZN => n37998);
   U1307 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_26_port, B1 => 
                           n37755, B2 => REGISTERS_19_26_port, ZN => n37997);
   U1308 : NAND4_X1 port map( A1 => n38000, A2 => n37999, A3 => n37998, A4 => 
                           n37997, ZN => n38001);
   U1309 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_27_port, B1 => 
                           n38205, B2 => REGISTERS_16_27_port, ZN => n38008);
   U1310 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_27_port, B1 => 
                           n38207, B2 => REGISTERS_24_27_port, ZN => n38007);
   U1311 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_27_port, B1 => 
                           n38209, B2 => REGISTERS_15_27_port, ZN => n38006);
   U1312 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_27_port, ZN => 
                           n38005);
   U1313 : NAND4_X1 port map( A1 => n38008, A2 => n38007, A3 => n38006, A4 => 
                           n38005, ZN => n38024);
   U1314 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_27_port, B1 => 
                           n38216, B2 => REGISTERS_22_27_port, ZN => n38012);
   U1315 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_27_port, B1 => 
                           n37735, B2 => REGISTERS_9_27_port, ZN => n38011);
   U1316 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_27_port, B1 => 
                           n38220, B2 => REGISTERS_31_27_port, ZN => n38010);
   U1317 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_27_port, B1 => 
                           n37739, B2 => REGISTERS_8_27_port, ZN => n38009);
   U1318 : NAND4_X1 port map( A1 => n38012, A2 => n38011, A3 => n38010, A4 => 
                           n38009, ZN => n38023);
   U1319 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_27_port, B1 => 
                           n38228, B2 => REGISTERS_29_27_port, ZN => n38016);
   U1320 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_27_port, B1 => 
                           n37743, B2 => REGISTERS_4_27_port, ZN => n38015);
   U1321 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_27_port, B1 => 
                           n38232, B2 => REGISTERS_28_27_port, ZN => n38014);
   U1322 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_27_port, B1 => 
                           n37747, B2 => REGISTERS_7_27_port, ZN => n38013);
   U1323 : NAND4_X1 port map( A1 => n38016, A2 => n38015, A3 => n38014, A4 => 
                           n38013, ZN => n38022);
   U1324 : AOI22_X1 port map( A1 => n37750, A2 => REGISTERS_26_27_port, B1 => 
                           n38240, B2 => REGISTERS_5_27_port, ZN => n38020);
   U1325 : AOI22_X1 port map( A1 => n37752, A2 => REGISTERS_21_27_port, B1 => 
                           n38242, B2 => REGISTERS_25_27_port, ZN => n38019);
   U1326 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_27_port, B1 => 
                           n38244, B2 => REGISTERS_17_27_port, ZN => n38018);
   U1327 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_27_port, B1 => 
                           n38246, B2 => REGISTERS_19_27_port, ZN => n38017);
   U1328 : NAND4_X1 port map( A1 => n38020, A2 => n38019, A3 => n38018, A4 => 
                           n38017, ZN => n38021);
   U1329 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_28_port, B1 => 
                           n37726, B2 => REGISTERS_16_28_port, ZN => n38028);
   U1330 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_28_port, B1 => 
                           n37728, B2 => REGISTERS_24_28_port, ZN => n38027);
   U1331 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_28_port, B1 => 
                           n38209, B2 => REGISTERS_15_28_port, ZN => n38026);
   U1332 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_28_port, ZN => 
                           n38025);
   U1333 : NAND4_X1 port map( A1 => n38028, A2 => n38027, A3 => n38026, A4 => 
                           n38025, ZN => n38044);
   U1334 : AOI22_X1 port map( A1 => n37734, A2 => REGISTERS_20_28_port, B1 => 
                           n37733, B2 => REGISTERS_22_28_port, ZN => n38032);
   U1335 : AOI22_X1 port map( A1 => n37736, A2 => REGISTERS_18_28_port, B1 => 
                           n38218, B2 => REGISTERS_9_28_port, ZN => n38031);
   U1336 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_28_port, B1 => 
                           n38220, B2 => REGISTERS_31_28_port, ZN => n38030);
   U1337 : AOI22_X1 port map( A1 => n37740, A2 => REGISTERS_3_28_port, B1 => 
                           n38222, B2 => REGISTERS_8_28_port, ZN => n38029);
   U1338 : NAND4_X1 port map( A1 => n38032, A2 => n38031, A3 => n38030, A4 => 
                           n38029, ZN => n38043);
   U1339 : AOI22_X1 port map( A1 => n37742, A2 => REGISTERS_30_28_port, B1 => 
                           n38228, B2 => REGISTERS_29_28_port, ZN => n38036);
   U1340 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_28_port, B1 => 
                           n37743, B2 => REGISTERS_4_28_port, ZN => n38035);
   U1341 : AOI22_X1 port map( A1 => n37746, A2 => REGISTERS_10_28_port, B1 => 
                           n38232, B2 => REGISTERS_28_28_port, ZN => n38034);
   U1342 : AOI22_X1 port map( A1 => n37748, A2 => REGISTERS_6_28_port, B1 => 
                           n38234, B2 => REGISTERS_7_28_port, ZN => n38033);
   U1343 : NAND4_X1 port map( A1 => n38036, A2 => n38035, A3 => n38034, A4 => 
                           n38033, ZN => n38042);
   U1344 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_28_port, B1 => 
                           n38240, B2 => REGISTERS_5_28_port, ZN => n38040);
   U1345 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_28_port, B1 => 
                           n38242, B2 => REGISTERS_25_28_port, ZN => n38039);
   U1346 : AOI22_X1 port map( A1 => n37754, A2 => REGISTERS_23_28_port, B1 => 
                           n38244, B2 => REGISTERS_17_28_port, ZN => n38038);
   U1347 : AOI22_X1 port map( A1 => n37756, A2 => REGISTERS_14_28_port, B1 => 
                           n38246, B2 => REGISTERS_19_28_port, ZN => n38037);
   U1348 : NAND4_X1 port map( A1 => n38040, A2 => n38039, A3 => n38038, A4 => 
                           n38037, ZN => n38041);
   U1349 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_29_port, B1 => 
                           n38205, B2 => REGISTERS_16_29_port, ZN => n38048);
   U1350 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_29_port, B1 => 
                           n38207, B2 => REGISTERS_24_29_port, ZN => n38047);
   U1351 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_29_port, B1 => 
                           n38209, B2 => REGISTERS_15_29_port, ZN => n38046);
   U1352 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_29_port, ZN => 
                           n38045);
   U1353 : NAND4_X1 port map( A1 => n38048, A2 => n38047, A3 => n38046, A4 => 
                           n38045, ZN => n38064);
   U1354 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_29_port, B1 => 
                           n38216, B2 => REGISTERS_22_29_port, ZN => n38052);
   U1355 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_29_port, B1 => 
                           n38218, B2 => REGISTERS_9_29_port, ZN => n38051);
   U1356 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_29_port, B1 => 
                           n38220, B2 => REGISTERS_31_29_port, ZN => n38050);
   U1357 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_29_port, B1 => 
                           n38222, B2 => REGISTERS_8_29_port, ZN => n38049);
   U1358 : NAND4_X1 port map( A1 => n38052, A2 => n38051, A3 => n38050, A4 => 
                           n38049, ZN => n38063);
   U1359 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_29_port, B1 => 
                           n38228, B2 => REGISTERS_29_29_port, ZN => n38056);
   U1360 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_29_port, B1 => 
                           n37743, B2 => REGISTERS_4_29_port, ZN => n38055);
   U1361 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_29_port, B1 => 
                           n38232, B2 => REGISTERS_28_29_port, ZN => n38054);
   U1362 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_29_port, B1 => 
                           n38234, B2 => REGISTERS_7_29_port, ZN => n38053);
   U1363 : NAND4_X1 port map( A1 => n38056, A2 => n38055, A3 => n38054, A4 => 
                           n38053, ZN => n38062);
   U1364 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_29_port, B1 => 
                           n38240, B2 => REGISTERS_5_29_port, ZN => n38060);
   U1365 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_29_port, B1 => 
                           n38242, B2 => REGISTERS_25_29_port, ZN => n38059);
   U1366 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_29_port, B1 => 
                           n38244, B2 => REGISTERS_17_29_port, ZN => n38058);
   U1367 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_29_port, B1 => 
                           n38246, B2 => REGISTERS_19_29_port, ZN => n38057);
   U1368 : NAND4_X1 port map( A1 => n38060, A2 => n38059, A3 => n38058, A4 => 
                           n38057, ZN => n38061);
   U1369 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_2_port, B1 => 
                           n38205, B2 => REGISTERS_16_2_port, ZN => n38068);
   U1370 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_2_port, B1 => 
                           n38207, B2 => REGISTERS_24_2_port, ZN => n38067);
   U1371 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_2_port, B1 => 
                           n38209, B2 => REGISTERS_15_2_port, ZN => n38066);
   U1372 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_2_port, ZN => 
                           n38065);
   U1373 : NAND4_X1 port map( A1 => n38068, A2 => n38067, A3 => n38066, A4 => 
                           n38065, ZN => n38084);
   U1374 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_2_port, B1 => 
                           n38216, B2 => REGISTERS_22_2_port, ZN => n38072);
   U1375 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_2_port, B1 => 
                           n38218, B2 => REGISTERS_9_2_port, ZN => n38071);
   U1376 : AOI22_X1 port map( A1 => n38221, A2 => REGISTERS_2_2_port, B1 => 
                           n38220, B2 => REGISTERS_31_2_port, ZN => n38070);
   U1377 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_2_port, B1 => 
                           n38222, B2 => REGISTERS_8_2_port, ZN => n38069);
   U1378 : NAND4_X1 port map( A1 => n38072, A2 => n38071, A3 => n38070, A4 => 
                           n38069, ZN => n38083);
   U1379 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_2_port, B1 => 
                           n38228, B2 => REGISTERS_29_2_port, ZN => n38076);
   U1380 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_2_port, B1 => 
                           n37743, B2 => REGISTERS_4_2_port, ZN => n38075);
   U1381 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_2_port, B1 => 
                           n38232, B2 => REGISTERS_28_2_port, ZN => n38074);
   U1382 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_2_port, B1 => 
                           n38234, B2 => REGISTERS_7_2_port, ZN => n38073);
   U1383 : NAND4_X1 port map( A1 => n38076, A2 => n38075, A3 => n38074, A4 => 
                           n38073, ZN => n38082);
   U1384 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_2_port, B1 => 
                           n38240, B2 => REGISTERS_5_2_port, ZN => n38080);
   U1385 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_2_port, B1 => 
                           n38242, B2 => REGISTERS_25_2_port, ZN => n38079);
   U1386 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_2_port, B1 => 
                           n38244, B2 => REGISTERS_17_2_port, ZN => n38078);
   U1387 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_2_port, B1 => 
                           n38246, B2 => REGISTERS_19_2_port, ZN => n38077);
   U1388 : NAND4_X1 port map( A1 => n38080, A2 => n38079, A3 => n38078, A4 => 
                           n38077, ZN => n38081);
   U1389 : AOI22_X1 port map( A1 => n37727, A2 => REGISTERS_11_30_port, B1 => 
                           n38205, B2 => REGISTERS_16_30_port, ZN => n38088);
   U1390 : AOI22_X1 port map( A1 => n37729, A2 => REGISTERS_1_30_port, B1 => 
                           n38207, B2 => REGISTERS_24_30_port, ZN => n38087);
   U1391 : AOI22_X1 port map( A1 => n37731, A2 => REGISTERS_12_30_port, B1 => 
                           n37730, B2 => REGISTERS_15_30_port, ZN => n38086);
   U1392 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_30_port, ZN => 
                           n38085);
   U1393 : NAND4_X1 port map( A1 => n38088, A2 => n38087, A3 => n38086, A4 => 
                           n38085, ZN => n38104);
   U1394 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_30_port, B1 => 
                           n38216, B2 => REGISTERS_22_30_port, ZN => n38092);
   U1395 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_30_port, B1 => 
                           n38218, B2 => REGISTERS_9_30_port, ZN => n38091);
   U1396 : AOI22_X1 port map( A1 => n38221, A2 => REGISTERS_2_30_port, B1 => 
                           n38220, B2 => REGISTERS_31_30_port, ZN => n38090);
   U1397 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_30_port, B1 => 
                           n38222, B2 => REGISTERS_8_30_port, ZN => n38089);
   U1398 : NAND4_X1 port map( A1 => n38092, A2 => n38091, A3 => n38090, A4 => 
                           n38089, ZN => n38103);
   U1399 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_30_port, B1 => 
                           n38228, B2 => REGISTERS_29_30_port, ZN => n38096);
   U1400 : AOI22_X1 port map( A1 => n37744, A2 => REGISTERS_27_30_port, B1 => 
                           n38230, B2 => REGISTERS_4_30_port, ZN => n38095);
   U1401 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_30_port, B1 => 
                           n38232, B2 => REGISTERS_28_30_port, ZN => n38094);
   U1402 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_30_port, B1 => 
                           n38234, B2 => REGISTERS_7_30_port, ZN => n38093);
   U1403 : NAND4_X1 port map( A1 => n38096, A2 => n38095, A3 => n38094, A4 => 
                           n38093, ZN => n38102);
   U1404 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_30_port, B1 => 
                           n38240, B2 => REGISTERS_5_30_port, ZN => n38100);
   U1405 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_30_port, B1 => 
                           n38242, B2 => REGISTERS_25_30_port, ZN => n38099);
   U1406 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_30_port, B1 => 
                           n38244, B2 => REGISTERS_17_30_port, ZN => n38098);
   U1407 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_30_port, B1 => 
                           n38246, B2 => REGISTERS_19_30_port, ZN => n38097);
   U1408 : NAND4_X1 port map( A1 => n38100, A2 => n38099, A3 => n38098, A4 => 
                           n38097, ZN => n38101);
   U1409 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_31_port, B1 => 
                           n38205, B2 => REGISTERS_16_31_port, ZN => n38108);
   U1410 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_31_port, B1 => 
                           n38207, B2 => REGISTERS_24_31_port, ZN => n38107);
   U1411 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_31_port, B1 => 
                           n38209, B2 => REGISTERS_15_31_port, ZN => n38106);
   U1412 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_31_port, ZN => 
                           n38105);
   U1413 : NAND4_X1 port map( A1 => n38108, A2 => n38107, A3 => n38106, A4 => 
                           n38105, ZN => n38124);
   U1414 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_31_port, B1 => 
                           n38216, B2 => REGISTERS_22_31_port, ZN => n38112);
   U1415 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_31_port, B1 => 
                           n38218, B2 => REGISTERS_9_31_port, ZN => n38111);
   U1416 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_31_port, B1 => 
                           n38220, B2 => REGISTERS_31_31_port, ZN => n38110);
   U1417 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_31_port, B1 => 
                           n38222, B2 => REGISTERS_8_31_port, ZN => n38109);
   U1418 : NAND4_X1 port map( A1 => n38112, A2 => n38111, A3 => n38110, A4 => 
                           n38109, ZN => n38123);
   U1419 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_31_port, B1 => 
                           n38228, B2 => REGISTERS_29_31_port, ZN => n38116);
   U1420 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_31_port, B1 => 
                           n38230, B2 => REGISTERS_4_31_port, ZN => n38115);
   U1421 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_31_port, B1 => 
                           n38232, B2 => REGISTERS_28_31_port, ZN => n38114);
   U1422 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_31_port, B1 => 
                           n38234, B2 => REGISTERS_7_31_port, ZN => n38113);
   U1423 : NAND4_X1 port map( A1 => n38116, A2 => n38115, A3 => n38114, A4 => 
                           n38113, ZN => n38122);
   U1424 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_31_port, B1 => 
                           n38240, B2 => REGISTERS_5_31_port, ZN => n38120);
   U1425 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_31_port, B1 => 
                           n38242, B2 => REGISTERS_25_31_port, ZN => n38119);
   U1426 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_31_port, B1 => 
                           n38244, B2 => REGISTERS_17_31_port, ZN => n38118);
   U1427 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_31_port, B1 => 
                           n38246, B2 => REGISTERS_19_31_port, ZN => n38117);
   U1428 : NAND4_X1 port map( A1 => n38120, A2 => n38119, A3 => n38118, A4 => 
                           n38117, ZN => n38121);
   U1429 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_3_port, B1 => 
                           n38205, B2 => REGISTERS_16_3_port, ZN => n38128);
   U1430 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_3_port, B1 => 
                           n38207, B2 => REGISTERS_24_3_port, ZN => n38127);
   U1431 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_3_port, B1 => 
                           n38209, B2 => REGISTERS_15_3_port, ZN => n38126);
   U1432 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_3_port, ZN => 
                           n38125);
   U1433 : NAND4_X1 port map( A1 => n38128, A2 => n38127, A3 => n38126, A4 => 
                           n38125, ZN => n38144);
   U1434 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_3_port, B1 => 
                           n38216, B2 => REGISTERS_22_3_port, ZN => n38132);
   U1435 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_3_port, B1 => 
                           n38218, B2 => REGISTERS_9_3_port, ZN => n38131);
   U1436 : AOI22_X1 port map( A1 => n38221, A2 => REGISTERS_2_3_port, B1 => 
                           n38220, B2 => REGISTERS_31_3_port, ZN => n38130);
   U1437 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_3_port, B1 => 
                           n38222, B2 => REGISTERS_8_3_port, ZN => n38129);
   U1438 : NAND4_X1 port map( A1 => n38132, A2 => n38131, A3 => n38130, A4 => 
                           n38129, ZN => n38143);
   U1439 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_3_port, B1 => 
                           n38228, B2 => REGISTERS_29_3_port, ZN => n38136);
   U1440 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_3_port, B1 => 
                           n38230, B2 => REGISTERS_4_3_port, ZN => n38135);
   U1441 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_3_port, B1 => 
                           n38232, B2 => REGISTERS_28_3_port, ZN => n38134);
   U1442 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_3_port, B1 => 
                           n38234, B2 => REGISTERS_7_3_port, ZN => n38133);
   U1443 : NAND4_X1 port map( A1 => n38136, A2 => n38135, A3 => n38134, A4 => 
                           n38133, ZN => n38142);
   U1444 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_3_port, B1 => 
                           n38240, B2 => REGISTERS_5_3_port, ZN => n38140);
   U1445 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_3_port, B1 => 
                           n38242, B2 => REGISTERS_25_3_port, ZN => n38139);
   U1446 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_3_port, B1 => 
                           n38244, B2 => REGISTERS_17_3_port, ZN => n38138);
   U1447 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_3_port, B1 => 
                           n38246, B2 => REGISTERS_19_3_port, ZN => n38137);
   U1448 : NAND4_X1 port map( A1 => n38140, A2 => n38139, A3 => n38138, A4 => 
                           n38137, ZN => n38141);
   U1449 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_5_port, B1 => 
                           n38205, B2 => REGISTERS_16_5_port, ZN => n38148);
   U1450 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_5_port, B1 => 
                           n38207, B2 => REGISTERS_24_5_port, ZN => n38147);
   U1451 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_5_port, B1 => 
                           n38209, B2 => REGISTERS_15_5_port, ZN => n38146);
   U1452 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_5_port, ZN => 
                           n38145);
   U1453 : NAND4_X1 port map( A1 => n38148, A2 => n38147, A3 => n38146, A4 => 
                           n38145, ZN => n38164);
   U1454 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_5_port, B1 => 
                           n38216, B2 => REGISTERS_22_5_port, ZN => n38152);
   U1455 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_5_port, B1 => 
                           n38218, B2 => REGISTERS_9_5_port, ZN => n38151);
   U1456 : AOI22_X1 port map( A1 => n38221, A2 => REGISTERS_2_5_port, B1 => 
                           n38220, B2 => REGISTERS_31_5_port, ZN => n38150);
   U1457 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_5_port, B1 => 
                           n38222, B2 => REGISTERS_8_5_port, ZN => n38149);
   U1458 : NAND4_X1 port map( A1 => n38152, A2 => n38151, A3 => n38150, A4 => 
                           n38149, ZN => n38163);
   U1459 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_5_port, B1 => 
                           n38228, B2 => REGISTERS_29_5_port, ZN => n38156);
   U1460 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_5_port, B1 => 
                           n38230, B2 => REGISTERS_4_5_port, ZN => n38155);
   U1461 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_5_port, B1 => 
                           n38232, B2 => REGISTERS_28_5_port, ZN => n38154);
   U1462 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_5_port, B1 => 
                           n38234, B2 => REGISTERS_7_5_port, ZN => n38153);
   U1463 : NAND4_X1 port map( A1 => n38156, A2 => n38155, A3 => n38154, A4 => 
                           n38153, ZN => n38162);
   U1464 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_5_port, B1 => 
                           n38240, B2 => REGISTERS_5_5_port, ZN => n38160);
   U1465 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_5_port, B1 => 
                           n38242, B2 => REGISTERS_25_5_port, ZN => n38159);
   U1466 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_5_port, B1 => 
                           n38244, B2 => REGISTERS_17_5_port, ZN => n38158);
   U1467 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_5_port, B1 => 
                           n38246, B2 => REGISTERS_19_5_port, ZN => n38157);
   U1468 : NAND4_X1 port map( A1 => n38160, A2 => n38159, A3 => n38158, A4 => 
                           n38157, ZN => n38161);
   U1469 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_6_port, B1 => 
                           n38205, B2 => REGISTERS_16_6_port, ZN => n38168);
   U1470 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_6_port, B1 => 
                           n38207, B2 => REGISTERS_24_6_port, ZN => n38167);
   U1471 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_6_port, B1 => 
                           n38209, B2 => REGISTERS_15_6_port, ZN => n38166);
   U1472 : NAND2_X1 port map( A1 => n38211, A2 => REGISTERS_13_6_port, ZN => 
                           n38165);
   U1473 : NAND4_X1 port map( A1 => n38168, A2 => n38167, A3 => n38166, A4 => 
                           n38165, ZN => n38184);
   U1474 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_6_port, B1 => 
                           n38216, B2 => REGISTERS_22_6_port, ZN => n38172);
   U1475 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_6_port, B1 => 
                           n38218, B2 => REGISTERS_9_6_port, ZN => n38171);
   U1476 : AOI22_X1 port map( A1 => n38221, A2 => REGISTERS_2_6_port, B1 => 
                           n38220, B2 => REGISTERS_31_6_port, ZN => n38170);
   U1477 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_6_port, B1 => 
                           n38222, B2 => REGISTERS_8_6_port, ZN => n38169);
   U1478 : NAND4_X1 port map( A1 => n38172, A2 => n38171, A3 => n38170, A4 => 
                           n38169, ZN => n38183);
   U1479 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_6_port, B1 => 
                           n38228, B2 => REGISTERS_29_6_port, ZN => n38176);
   U1480 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_6_port, B1 => 
                           n38230, B2 => REGISTERS_4_6_port, ZN => n38175);
   U1481 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_6_port, B1 => 
                           n38232, B2 => REGISTERS_28_6_port, ZN => n38174);
   U1482 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_6_port, B1 => 
                           n38234, B2 => REGISTERS_7_6_port, ZN => n38173);
   U1483 : NAND4_X1 port map( A1 => n38176, A2 => n38175, A3 => n38174, A4 => 
                           n38173, ZN => n38182);
   U1484 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_6_port, B1 => 
                           n38240, B2 => REGISTERS_5_6_port, ZN => n38180);
   U1485 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_6_port, B1 => 
                           n38242, B2 => REGISTERS_25_6_port, ZN => n38179);
   U1486 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_6_port, B1 => 
                           n38244, B2 => REGISTERS_17_6_port, ZN => n38178);
   U1487 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_6_port, B1 => 
                           n38246, B2 => REGISTERS_19_6_port, ZN => n38177);
   U1488 : NAND4_X1 port map( A1 => n38180, A2 => n38179, A3 => n38178, A4 => 
                           n38177, ZN => n38181);
   U1489 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_8_port, B1 => 
                           n38205, B2 => REGISTERS_16_8_port, ZN => n38188);
   U1490 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_8_port, B1 => 
                           n38207, B2 => REGISTERS_24_8_port, ZN => n38187);
   U1491 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_8_port, B1 => 
                           n38209, B2 => REGISTERS_15_8_port, ZN => n38186);
   U1492 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_8_port, ZN => 
                           n38185);
   U1493 : NAND4_X1 port map( A1 => n38188, A2 => n38187, A3 => n38186, A4 => 
                           n38185, ZN => n38204);
   U1494 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_8_port, B1 => 
                           n38216, B2 => REGISTERS_22_8_port, ZN => n38192);
   U1495 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_8_port, B1 => 
                           n38218, B2 => REGISTERS_9_8_port, ZN => n38191);
   U1496 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_8_port, B1 => 
                           n38220, B2 => REGISTERS_31_8_port, ZN => n38190);
   U1497 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_8_port, B1 => 
                           n38222, B2 => REGISTERS_8_8_port, ZN => n38189);
   U1498 : NAND4_X1 port map( A1 => n38192, A2 => n38191, A3 => n38190, A4 => 
                           n38189, ZN => n38203);
   U1499 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_8_port, B1 => 
                           n38228, B2 => REGISTERS_29_8_port, ZN => n38196);
   U1500 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_8_port, B1 => 
                           n37743, B2 => REGISTERS_4_8_port, ZN => n38195);
   U1501 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_8_port, B1 => 
                           n38232, B2 => REGISTERS_28_8_port, ZN => n38194);
   U1502 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_8_port, B1 => 
                           n38234, B2 => REGISTERS_7_8_port, ZN => n38193);
   U1503 : NAND4_X1 port map( A1 => n38196, A2 => n38195, A3 => n38194, A4 => 
                           n38193, ZN => n38202);
   U1504 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_8_port, B1 => 
                           n38240, B2 => REGISTERS_5_8_port, ZN => n38200);
   U1505 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_8_port, B1 => 
                           n38242, B2 => REGISTERS_25_8_port, ZN => n38199);
   U1506 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_8_port, B1 => 
                           n38244, B2 => REGISTERS_17_8_port, ZN => n38198);
   U1507 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_8_port, B1 => 
                           n38246, B2 => REGISTERS_19_8_port, ZN => n38197);
   U1508 : NAND4_X1 port map( A1 => n38200, A2 => n38199, A3 => n38198, A4 => 
                           n38197, ZN => n38201);
   U1509 : AOI22_X1 port map( A1 => n38206, A2 => REGISTERS_11_9_port, B1 => 
                           n38205, B2 => REGISTERS_16_9_port, ZN => n38215);
   U1510 : AOI22_X1 port map( A1 => n38208, A2 => REGISTERS_1_9_port, B1 => 
                           n38207, B2 => REGISTERS_24_9_port, ZN => n38214);
   U1511 : AOI22_X1 port map( A1 => n38210, A2 => REGISTERS_12_9_port, B1 => 
                           n38209, B2 => REGISTERS_15_9_port, ZN => n38213);
   U1512 : NAND2_X1 port map( A1 => n37732, A2 => REGISTERS_13_9_port, ZN => 
                           n38212);
   U1513 : NAND4_X1 port map( A1 => n38215, A2 => n38214, A3 => n38213, A4 => 
                           n38212, ZN => n38255);
   U1514 : AOI22_X1 port map( A1 => n38217, A2 => REGISTERS_20_9_port, B1 => 
                           n38216, B2 => REGISTERS_22_9_port, ZN => n38227);
   U1515 : AOI22_X1 port map( A1 => n38219, A2 => REGISTERS_18_9_port, B1 => 
                           n38218, B2 => REGISTERS_9_9_port, ZN => n38226);
   U1516 : AOI22_X1 port map( A1 => n37738, A2 => REGISTERS_2_9_port, B1 => 
                           n37737, B2 => REGISTERS_31_9_port, ZN => n38225);
   U1517 : AOI22_X1 port map( A1 => n38223, A2 => REGISTERS_3_9_port, B1 => 
                           n38222, B2 => REGISTERS_8_9_port, ZN => n38224);
   U1518 : NAND4_X1 port map( A1 => n38227, A2 => n38226, A3 => n38225, A4 => 
                           n38224, ZN => n38254);
   U1519 : AOI22_X1 port map( A1 => n38229, A2 => REGISTERS_30_9_port, B1 => 
                           n37741, B2 => REGISTERS_29_9_port, ZN => n38239);
   U1520 : AOI22_X1 port map( A1 => n38231, A2 => REGISTERS_27_9_port, B1 => 
                           n37743, B2 => REGISTERS_4_9_port, ZN => n38238);
   U1521 : AOI22_X1 port map( A1 => n38233, A2 => REGISTERS_10_9_port, B1 => 
                           n37745, B2 => REGISTERS_28_9_port, ZN => n38237);
   U1522 : AOI22_X1 port map( A1 => n38235, A2 => REGISTERS_6_9_port, B1 => 
                           n38234, B2 => REGISTERS_7_9_port, ZN => n38236);
   U1523 : NAND4_X1 port map( A1 => n38239, A2 => n38238, A3 => n38237, A4 => 
                           n38236, ZN => n38253);
   U1524 : AOI22_X1 port map( A1 => n38241, A2 => REGISTERS_26_9_port, B1 => 
                           n37749, B2 => REGISTERS_5_9_port, ZN => n38251);
   U1525 : AOI22_X1 port map( A1 => n38243, A2 => REGISTERS_21_9_port, B1 => 
                           n38242, B2 => REGISTERS_25_9_port, ZN => n38250);
   U1526 : AOI22_X1 port map( A1 => n38245, A2 => REGISTERS_23_9_port, B1 => 
                           n38244, B2 => REGISTERS_17_9_port, ZN => n38249);
   U1527 : AOI22_X1 port map( A1 => n38247, A2 => REGISTERS_14_9_port, B1 => 
                           n38246, B2 => REGISTERS_19_9_port, ZN => n38248);
   U1528 : NAND4_X1 port map( A1 => n38251, A2 => n38250, A3 => n38249, A4 => 
                           n38248, ZN => n38252);
   U1529 : INV_X1 port map( A => ADD_RDB(2), ZN => n38260);
   U1530 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDB(1), A3 => n38260, ZN 
                           => n38270);
   U1531 : INV_X1 port map( A => ADD_RDB(4), ZN => n38259);
   U1532 : NAND3_X1 port map( A1 => ADD_RDB(3), A2 => ADD_RDB(0), A3 => n38259,
                           ZN => n38262);
   U1533 : NOR2_X1 port map( A1 => n38270, A2 => n38262, ZN => n38276);
   U1534 : NAND3_X1 port map( A1 => ADD_RDB(4), A2 => ADD_RDB(3), A3 => 
                           ADD_RDB(0), ZN => n38267);
   U1535 : INV_X1 port map( A => ADD_RDB(1), ZN => n38256);
   U1536 : NAND3_X1 port map( A1 => RESET, A2 => n38260, A3 => n38256, ZN => 
                           n38266);
   U1537 : NOR2_X1 port map( A1 => n38267, A2 => n38266, ZN => n38275);
   U1538 : NOR2_X1 port map( A1 => ADD_RDB(3), A2 => ADD_RDB(0), ZN => n38261);
   U1539 : NAND3_X1 port map( A1 => RESET, A2 => n38261, A3 => n38259, ZN => 
                           n38264);
   U1540 : NOR3_X1 port map( A1 => ADD_RDB(2), A2 => n38256, A3 => n38264, ZN 
                           => n38278);
   U1541 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDB(2), A3 => ADD_RDB(1), 
                           ZN => n38271);
   U1542 : NAND3_X1 port map( A1 => ADD_RDB(2), A2 => RESET, A3 => n38256, ZN 
                           => n38274);
   U1543 : NOR2_X1 port map( A1 => n38262, A2 => n38274, ZN => n38280);
   U1544 : NOR2_X1 port map( A1 => n38267, A2 => n38274, ZN => n38279);
   U1545 : INV_X1 port map( A => ADD_RDB(3), ZN => n38258);
   U1546 : NAND3_X1 port map( A1 => ADD_RDB(4), A2 => ADD_RDB(0), A3 => n38258,
                           ZN => n38268);
   U1547 : NOR2_X1 port map( A1 => n38270, A2 => n38268, ZN => n38281);
   U1548 : INV_X1 port map( A => ADD_RDB(0), ZN => n38257);
   U1549 : NAND3_X1 port map( A1 => ADD_RDB(3), A2 => n38259, A3 => n38257, ZN 
                           => n38265);
   U1550 : NOR2_X1 port map( A1 => n38266, A2 => n38265, ZN => n38283);
   U1551 : NAND3_X1 port map( A1 => ADD_RDB(3), A2 => ADD_RDB(4), A3 => n38257,
                           ZN => n38272);
   U1552 : NOR2_X1 port map( A1 => n38270, A2 => n38272, ZN => n38282);
   U1553 : NAND3_X1 port map( A1 => ADD_RDB(0), A2 => n38259, A3 => n38258, ZN 
                           => n38273);
   U1554 : NOR2_X1 port map( A1 => n38270, A2 => n38273, ZN => n38285);
   U1555 : NOR2_X1 port map( A1 => n38271, A2 => n38272, ZN => n38284);
   U1556 : NOR3_X1 port map( A1 => ADD_RDB(1), A2 => n38260, A3 => n38264, ZN 
                           => n38287);
   U1557 : NOR2_X1 port map( A1 => n38268, A2 => n38266, ZN => n38286);
   U1558 : NAND2_X1 port map( A1 => ADD_RDB(4), A2 => n38261, ZN => n38269);
   U1559 : NOR2_X1 port map( A1 => n38271, A2 => n38269, ZN => n38288);
   U1560 : NOR2_X1 port map( A1 => n38266, A2 => n38269, ZN => n38291);
   U1561 : NOR2_X1 port map( A1 => n38262, A2 => n38266, ZN => n38290);
   U1562 : NAND2_X1 port map( A1 => ADD_RDB(2), A2 => ADD_RDB(1), ZN => n38263)
                           ;
   U1563 : NOR2_X1 port map( A1 => n38264, A2 => n38263, ZN => n38293);
   U1564 : NOR2_X1 port map( A1 => n38268, A2 => n38271, ZN => n38292);
   U1565 : NOR2_X1 port map( A1 => n38266, A2 => n38272, ZN => n38295);
   U1566 : NOR2_X1 port map( A1 => n38271, A2 => n38265, ZN => n38294);
   U1567 : NOR2_X1 port map( A1 => n38274, A2 => n38265, ZN => n38297);
   U1568 : NOR2_X1 port map( A1 => n38270, A2 => n38265, ZN => n38296);
   U1569 : NOR2_X1 port map( A1 => n38266, A2 => n38273, ZN => n38299);
   U1570 : NOR2_X1 port map( A1 => n38270, A2 => n38267, ZN => n38298);
   U1571 : NOR2_X1 port map( A1 => n38274, A2 => n38269, ZN => n38301);
   U1572 : NOR2_X1 port map( A1 => n38268, A2 => n38274, ZN => n38300);
   U1573 : NOR2_X1 port map( A1 => n38270, A2 => n38269, ZN => n38303);
   U1574 : NOR2_X1 port map( A1 => n38271, A2 => n38273, ZN => n38302);
   U1575 : NOR2_X1 port map( A1 => n38274, A2 => n38272, ZN => n38305);
   U1576 : NOR2_X1 port map( A1 => n38274, A2 => n38273, ZN => n38304);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity DLX_syn is

   port( Clk, Rst : in std_logic;  IRAM_DATA_OUT, DRAM_DATA_OUT : in 
         std_logic_vector (31 downto 0);  DRAM_DATA_IN : out std_logic_vector 
         (31 downto 0);  DRAM_ADDRESS : out std_logic_vector (11 downto 0);  
         DRAM_ENABLE, DRAM_RW : out std_logic;  DRAM_SEL : out std_logic_vector
         (2 downto 0);  IRAM_ADDRESS : out std_logic_vector (7 downto 0));

end DLX_syn;

architecture SYN_structural of DLX_syn is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X2
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_IF_ID
      port( CLK, EN : in std_logic;  ENCLK : out std_logic;  TE : in std_logic
            );
   end component;
   
   component branch_predictor
      port( RST : in std_logic;  PC_IN, PC_FAIL, IR_IN : in std_logic_vector 
            (31 downto 0);  IR_FAIL : in std_logic_vector (15 downto 0);  
            WRONG_PRE, RIGHT_PRE : in std_logic;  NPC_OUT, LINK_ADD : out 
            std_logic_vector (31 downto 0);  SEL, TAKEN : out std_logic);
   end component;
   
   component register_file_N32_addBit5
      port( RESET, RE, WE : in std_logic;  ADD_WR, ADD_RDA, ADD_RDB : in 
            std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
            downto 0);  OUTA, OUTB : out std_logic_vector (31 downto 0));
   end component;
   
   signal DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, IR_CU_31, IR_CU_28, IR_CU_27, 
      IR_CU_26, IR_CU_9_port, IR_CU_8_port, IR_CU_7_port, IR_CU_6_port, 
      IR_CU_5_port, IR_CU_4_port, IR_CU_1_port, IR_CU_0_port, BR_EN_i, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, 
      ALU_OPCODE_i_0_port, WB_MUX_SEL_i_1_port, RF_WE_i, 
      CU_I_aluOpcode_i_0_port, CU_I_aluOpcode_i_1_port, CU_I_aluOpcode_i_2_port
      , CU_I_aluOpcode_i_3_port, CU_I_aluOpcode_i_4_port, CU_I_cw2_1_port, 
      CU_I_cw_0_port, CU_I_cw_1_port, CU_I_cw_3_port, CU_I_cw_4_port, 
      CU_I_cw_6_port, CU_I_cw_7_port, CU_I_cw_9_port, CU_I_cw_10_port, 
      DataP_LMD_out_0_port, DataP_LMD_out_1_port, DataP_LMD_out_2_port, 
      DataP_LMD_out_3_port, DataP_LMD_out_4_port, DataP_LMD_out_5_port, 
      DataP_LMD_out_6_port, DataP_LMD_out_7_port, DataP_LMD_out_8_port, 
      DataP_LMD_out_9_port, DataP_LMD_out_10_port, DataP_LMD_out_11_port, 
      DataP_LMD_out_12_port, DataP_LMD_out_13_port, DataP_LMD_out_14_port, 
      DataP_LMD_out_15_port, DataP_LMD_out_16_port, DataP_LMD_out_17_port, 
      DataP_LMD_out_18_port, DataP_LMD_out_19_port, DataP_LMD_out_20_port, 
      DataP_LMD_out_21_port, DataP_LMD_out_22_port, DataP_LMD_out_23_port, 
      DataP_LMD_out_24_port, DataP_LMD_out_25_port, DataP_LMD_out_26_port, 
      DataP_LMD_out_27_port, DataP_LMD_out_28_port, DataP_LMD_out_29_port, 
      DataP_LMD_out_30_port, DataP_LMD_out_31_port, DataP_link_addr_W_0_port, 
      DataP_link_addr_W_1_port, DataP_link_addr_W_2_port, 
      DataP_link_addr_W_3_port, DataP_link_addr_W_4_port, 
      DataP_link_addr_W_5_port, DataP_link_addr_W_6_port, 
      DataP_link_addr_W_7_port, DataP_link_addr_W_8_port, 
      DataP_link_addr_W_9_port, DataP_link_addr_W_10_port, 
      DataP_link_addr_W_11_port, DataP_link_addr_W_12_port, 
      DataP_link_addr_W_13_port, DataP_link_addr_W_14_port, 
      DataP_link_addr_W_15_port, DataP_link_addr_W_16_port, 
      DataP_link_addr_W_17_port, DataP_link_addr_W_18_port, 
      DataP_link_addr_W_19_port, DataP_link_addr_W_20_port, 
      DataP_link_addr_W_21_port, DataP_link_addr_W_22_port, 
      DataP_link_addr_W_23_port, DataP_link_addr_W_24_port, 
      DataP_link_addr_W_25_port, DataP_link_addr_W_26_port, 
      DataP_link_addr_W_27_port, DataP_link_addr_W_28_port, 
      DataP_link_addr_W_29_port, DataP_link_addr_W_30_port, 
      DataP_link_addr_W_31_port, DataP_FWD_MUX_BR_S_0_port, 
      DataP_FWD_MUX_BR_S_1_port, DataP_alu_b_in_0_port, DataP_alu_b_in_2_port, 
      DataP_alu_b_in_3_port, DataP_alu_b_in_5_port, DataP_alu_b_in_6_port, 
      DataP_alu_b_in_7_port, DataP_alu_b_in_8_port, DataP_alu_b_in_9_port, 
      DataP_alu_b_in_10_port, DataP_alu_b_in_12_port, DataP_alu_b_in_13_port, 
      DataP_alu_b_in_15_port, DataP_alu_b_in_16_port, DataP_alu_b_in_17_port, 
      DataP_alu_b_in_18_port, DataP_alu_b_in_19_port, DataP_alu_b_in_20_port, 
      DataP_alu_b_in_21_port, DataP_alu_b_in_22_port, DataP_alu_b_in_23_port, 
      DataP_alu_b_in_24_port, DataP_alu_b_in_25_port, DataP_alu_b_in_26_port, 
      DataP_alu_b_in_27_port, DataP_alu_b_in_28_port, DataP_alu_b_in_29_port, 
      DataP_alu_b_in_30_port, DataP_alu_b_in_31_port, DataP_alu_a_in_0_port, 
      DataP_alu_a_in_1_port, DataP_alu_a_in_2_port, DataP_alu_a_in_3_port, 
      DataP_alu_a_in_4_port, DataP_alu_a_in_5_port, DataP_alu_a_in_6_port, 
      DataP_alu_a_in_7_port, DataP_alu_a_in_8_port, DataP_alu_a_in_9_port, 
      DataP_alu_a_in_10_port, DataP_alu_a_in_11_port, DataP_alu_a_in_12_port, 
      DataP_alu_a_in_13_port, DataP_alu_a_in_14_port, DataP_alu_a_in_15_port, 
      DataP_alu_a_in_16_port, DataP_alu_a_in_17_port, DataP_alu_a_in_18_port, 
      DataP_alu_a_in_19_port, DataP_alu_a_in_20_port, DataP_alu_a_in_21_port, 
      DataP_alu_a_in_22_port, DataP_alu_a_in_23_port, DataP_alu_a_in_24_port, 
      DataP_alu_a_in_25_port, DataP_alu_a_in_26_port, DataP_alu_a_in_27_port, 
      DataP_alu_a_in_28_port, DataP_alu_a_in_29_port, DataP_alu_a_in_30_port, 
      DataP_alu_a_in_31_port, DataP_alu_out_W_0_port, DataP_alu_out_W_1_port, 
      DataP_alu_out_W_2_port, DataP_alu_out_W_3_port, DataP_alu_out_W_4_port, 
      DataP_alu_out_W_5_port, DataP_alu_out_W_6_port, DataP_alu_out_W_7_port, 
      DataP_alu_out_W_8_port, DataP_alu_out_W_9_port, DataP_alu_out_W_10_port, 
      DataP_alu_out_W_11_port, DataP_alu_out_W_12_port, DataP_alu_out_W_13_port
      , DataP_alu_out_W_14_port, DataP_alu_out_W_15_port, 
      DataP_alu_out_W_16_port, DataP_alu_out_W_17_port, DataP_alu_out_W_18_port
      , DataP_alu_out_W_19_port, DataP_alu_out_W_20_port, 
      DataP_alu_out_W_21_port, DataP_alu_out_W_22_port, DataP_alu_out_W_23_port
      , DataP_alu_out_W_24_port, DataP_alu_out_W_25_port, 
      DataP_alu_out_W_26_port, DataP_alu_out_W_27_port, DataP_alu_out_W_28_port
      , DataP_alu_out_W_29_port, DataP_alu_out_W_30_port, 
      DataP_alu_out_W_31_port, DataP_alu_out_M_12_port, DataP_alu_out_M_13_port
      , DataP_alu_out_M_14_port, DataP_alu_out_M_15_port, 
      DataP_alu_out_M_16_port, DataP_alu_out_M_17_port, DataP_alu_out_M_18_port
      , DataP_alu_out_M_19_port, DataP_alu_out_M_20_port, 
      DataP_alu_out_M_21_port, DataP_alu_out_M_22_port, DataP_alu_out_M_23_port
      , DataP_alu_out_M_24_port, DataP_alu_out_M_25_port, 
      DataP_alu_out_M_26_port, DataP_alu_out_M_27_port, DataP_alu_out_M_28_port
      , DataP_alu_out_M_29_port, DataP_alu_out_M_30_port, 
      DataP_alu_out_M_31_port, DataP_opcode_W_0_port, DataP_opcode_W_1_port, 
      DataP_opcode_W_2_port, DataP_opcode_W_3_port, DataP_opcode_W_4_port, 
      DataP_opcode_W_5_port, DataP_opcode_M_0_port, DataP_opcode_M_1_port, 
      DataP_opcode_M_3_port, DataP_opcode_M_4_port, DataP_opcode_M_5_port, 
      DataP_dest_M_0_port, DataP_dest_M_1_port, DataP_dest_M_2_port, 
      DataP_dest_M_3_port, DataP_dest_M_4_port, DataP_pr_E, 
      DataP_opcode_E_0_port, DataP_opcode_E_3_port, DataP_opcode_E_4_port, 
      DataP_Rs2_0_port, DataP_Rs2_1_port, DataP_Rs2_2_port, DataP_Rs2_3_port, 
      DataP_Rs2_4_port, DataP_Rs1_1_port, DataP_Rs1_2_port, DataP_IMM_s_16_port
      , DataP_IMM_s_17_port, DataP_IMM_s_18_port, DataP_IMM_s_19_port, 
      DataP_IMM_s_20_port, DataP_IMM_s_21_port, DataP_IMM_s_22_port, 
      DataP_IMM_s_23_port, DataP_IMM_s_24_port, DataP_IMM_s_31_port, 
      DataP_B_s_0_port, DataP_B_s_1_port, DataP_B_s_2_port, DataP_B_s_3_port, 
      DataP_B_s_4_port, DataP_B_s_5_port, DataP_B_s_6_port, DataP_B_s_7_port, 
      DataP_B_s_8_port, DataP_B_s_9_port, DataP_B_s_10_port, DataP_B_s_11_port,
      DataP_B_s_12_port, DataP_B_s_13_port, DataP_B_s_14_port, 
      DataP_B_s_15_port, DataP_B_s_16_port, DataP_B_s_17_port, 
      DataP_B_s_18_port, DataP_B_s_19_port, DataP_B_s_20_port, 
      DataP_B_s_21_port, DataP_B_s_22_port, DataP_B_s_23_port, 
      DataP_B_s_24_port, DataP_B_s_25_port, DataP_B_s_26_port, 
      DataP_B_s_27_port, DataP_B_s_28_port, DataP_B_s_29_port, 
      DataP_B_s_30_port, DataP_B_s_31_port, DataP_A_s_0_port, DataP_A_s_1_port,
      DataP_A_s_2_port, DataP_A_s_3_port, DataP_A_s_4_port, DataP_A_s_5_port, 
      DataP_A_s_6_port, DataP_A_s_7_port, DataP_A_s_8_port, DataP_A_s_9_port, 
      DataP_A_s_10_port, DataP_A_s_11_port, DataP_A_s_12_port, 
      DataP_A_s_13_port, DataP_A_s_14_port, DataP_A_s_15_port, 
      DataP_A_s_16_port, DataP_A_s_17_port, DataP_A_s_18_port, 
      DataP_A_s_19_port, DataP_A_s_20_port, DataP_A_s_21_port, 
      DataP_A_s_22_port, DataP_A_s_23_port, DataP_A_s_24_port, 
      DataP_A_s_25_port, DataP_A_s_26_port, DataP_A_s_27_port, 
      DataP_A_s_28_port, DataP_A_s_29_port, DataP_A_s_30_port, 
      DataP_A_s_31_port, DataP_imm_out_16_port, DataP_imm_out_17_port, 
      DataP_imm_out_18_port, DataP_imm_out_19_port, DataP_imm_out_20_port, 
      DataP_imm_out_21_port, DataP_imm_out_22_port, DataP_imm_out_23_port, 
      DataP_imm_out_24_port, DataP_imm_out_31_port, DataP_b_out_0_port, 
      DataP_b_out_1_port, DataP_b_out_2_port, DataP_b_out_3_port, 
      DataP_b_out_4_port, DataP_b_out_5_port, DataP_b_out_6_port, 
      DataP_b_out_7_port, DataP_b_out_8_port, DataP_b_out_9_port, 
      DataP_b_out_10_port, DataP_b_out_11_port, DataP_b_out_12_port, 
      DataP_b_out_13_port, DataP_b_out_14_port, DataP_b_out_15_port, 
      DataP_b_out_16_port, DataP_b_out_17_port, DataP_b_out_18_port, 
      DataP_b_out_19_port, DataP_b_out_20_port, DataP_b_out_21_port, 
      DataP_b_out_22_port, DataP_b_out_23_port, DataP_b_out_24_port, 
      DataP_b_out_25_port, DataP_b_out_26_port, DataP_b_out_27_port, 
      DataP_b_out_28_port, DataP_b_out_29_port, DataP_b_out_30_port, 
      DataP_b_out_31_port, DataP_a_out_0_port, DataP_a_out_1_port, 
      DataP_a_out_2_port, DataP_a_out_3_port, DataP_a_out_4_port, 
      DataP_a_out_5_port, DataP_a_out_6_port, DataP_a_out_7_port, 
      DataP_a_out_8_port, DataP_a_out_9_port, DataP_a_out_10_port, 
      DataP_a_out_11_port, DataP_a_out_12_port, DataP_a_out_13_port, 
      DataP_a_out_14_port, DataP_a_out_15_port, DataP_a_out_16_port, 
      DataP_a_out_17_port, DataP_a_out_18_port, DataP_a_out_19_port, 
      DataP_a_out_20_port, DataP_a_out_21_port, DataP_a_out_22_port, 
      DataP_a_out_23_port, DataP_a_out_24_port, DataP_a_out_25_port, 
      DataP_a_out_26_port, DataP_a_out_27_port, DataP_a_out_28_port, 
      DataP_a_out_29_port, DataP_a_out_30_port, DataP_a_out_31_port, 
      DataP_WB_0_port, DataP_WB_1_port, DataP_WB_2_port, DataP_WB_3_port, 
      DataP_WB_4_port, DataP_WB_5_port, DataP_WB_6_port, DataP_WB_7_port, 
      DataP_WB_8_port, DataP_WB_9_port, DataP_WB_10_port, DataP_WB_11_port, 
      DataP_WB_12_port, DataP_WB_13_port, DataP_WB_14_port, DataP_WB_15_port, 
      DataP_WB_16_port, DataP_WB_17_port, DataP_WB_18_port, DataP_WB_19_port, 
      DataP_WB_20_port, DataP_WB_21_port, DataP_WB_22_port, DataP_WB_23_port, 
      DataP_WB_24_port, DataP_WB_25_port, DataP_WB_26_port, DataP_WB_27_port, 
      DataP_WB_28_port, DataP_WB_29_port, DataP_WB_30_port, DataP_WB_31_port, 
      DataP_add_D_0_port, DataP_add_D_1_port, DataP_add_D_2_port, 
      DataP_add_D_3_port, DataP_add_D_4_port, DataP_dest_D_0_port, 
      DataP_dest_D_1_port, DataP_dest_D_2_port, DataP_dest_D_3_port, 
      DataP_dest_D_4_port, DataP_add_S2_0_port, DataP_add_S2_1_port, 
      DataP_add_S2_2_port, DataP_add_S2_3_port, DataP_add_S2_4_port, 
      DataP_prediction, DataP_npc_mux_sel, DataP_link_addr_F_0_port, 
      DataP_link_addr_F_1_port, DataP_link_addr_F_2_port, 
      DataP_link_addr_F_3_port, DataP_link_addr_F_4_port, 
      DataP_link_addr_F_5_port, DataP_link_addr_F_6_port, 
      DataP_link_addr_F_7_port, DataP_link_addr_F_8_port, 
      DataP_link_addr_F_9_port, DataP_link_addr_F_10_port, 
      DataP_link_addr_F_11_port, DataP_link_addr_F_12_port, 
      DataP_link_addr_F_13_port, DataP_link_addr_F_14_port, 
      DataP_link_addr_F_15_port, DataP_link_addr_F_16_port, 
      DataP_link_addr_F_17_port, DataP_link_addr_F_18_port, 
      DataP_link_addr_F_19_port, DataP_link_addr_F_20_port, 
      DataP_link_addr_F_21_port, DataP_link_addr_F_22_port, 
      DataP_link_addr_F_23_port, DataP_link_addr_F_24_port, 
      DataP_link_addr_F_25_port, DataP_link_addr_F_26_port, 
      DataP_link_addr_F_27_port, DataP_link_addr_F_28_port, 
      DataP_link_addr_F_29_port, DataP_link_addr_F_30_port, 
      DataP_link_addr_F_31_port, DataP_npc_pre_0_port, DataP_npc_pre_1_port, 
      DataP_npc_pre_2_port, DataP_npc_pre_3_port, DataP_npc_pre_4_port, 
      DataP_npc_pre_5_port, DataP_npc_pre_6_port, DataP_npc_pre_7_port, 
      DataP_npc_pre_8_port, DataP_npc_pre_9_port, DataP_npc_pre_10_port, 
      DataP_npc_pre_11_port, DataP_npc_pre_12_port, DataP_npc_pre_13_port, 
      DataP_npc_pre_14_port, DataP_npc_pre_15_port, DataP_npc_pre_16_port, 
      DataP_npc_pre_17_port, DataP_npc_pre_18_port, DataP_npc_pre_19_port, 
      DataP_npc_pre_20_port, DataP_npc_pre_21_port, DataP_npc_pre_22_port, 
      DataP_npc_pre_23_port, DataP_npc_pre_24_port, DataP_npc_pre_25_port, 
      DataP_npc_pre_26_port, DataP_npc_pre_27_port, DataP_npc_pre_28_port, 
      DataP_npc_pre_29_port, DataP_npc_pre_30_port, DataP_npc_pre_31_port, 
      DataP_right_br, DataP_wrong_br, DataP_ir_E_0_port, DataP_ir_E_1_port, 
      DataP_ir_E_2_port, DataP_ir_E_3_port, DataP_ir_E_4_port, 
      DataP_ir_E_5_port, DataP_ir_E_6_port, DataP_ir_E_7_port, 
      DataP_ir_E_8_port, DataP_ir_E_9_port, DataP_ir_E_10_port, 
      DataP_ir_E_11_port, DataP_ir_E_12_port, DataP_ir_E_13_port, 
      DataP_ir_E_14_port, DataP_ir_E_15_port, DataP_npc_M_0_port, 
      DataP_npc_M_1_port, DataP_npc_M_2_port, DataP_npc_M_3_port, 
      DataP_npc_M_4_port, DataP_npc_M_5_port, DataP_npc_M_6_port, 
      DataP_npc_M_7_port, DataP_npc_M_8_port, DataP_npc_M_9_port, 
      DataP_npc_M_10_port, DataP_npc_M_11_port, DataP_npc_M_12_port, 
      DataP_npc_M_13_port, DataP_npc_M_14_port, DataP_npc_M_15_port, 
      DataP_npc_M_16_port, DataP_npc_M_17_port, DataP_npc_M_18_port, 
      DataP_npc_M_19_port, DataP_npc_M_20_port, DataP_npc_M_21_port, 
      DataP_npc_M_22_port, DataP_npc_M_23_port, DataP_npc_M_24_port, 
      DataP_npc_M_25_port, DataP_npc_M_26_port, DataP_npc_M_27_port, 
      DataP_npc_M_28_port, DataP_npc_M_29_port, DataP_npc_M_30_port, 
      DataP_npc_M_31_port, DataP_pc_out_0, DataP_pc_out_1, DataP_pc_out_10_port
      , DataP_pc_out_11_port, DataP_pc_out_12_port, DataP_pc_out_13_port, 
      DataP_pc_out_14_port, DataP_pc_out_15_port, DataP_pc_out_16_port, 
      DataP_pc_out_17_port, DataP_pc_out_18_port, DataP_pc_out_19_port, 
      DataP_pc_out_20_port, DataP_pc_out_21_port, DataP_pc_out_22_port, 
      DataP_pc_out_23_port, DataP_pc_out_24_port, DataP_pc_out_25_port, 
      DataP_pc_out_26_port, DataP_pc_out_27_port, DataP_pc_out_28_port, 
      DataP_pc_out_29_port, DataP_pc_out_30_port, DataP_pc_out_31_port, 
      DataP_npc_0_port, DataP_npc_1_port, DataP_npc_2_port, DataP_npc_3_port, 
      DataP_npc_4_port, DataP_npc_5_port, DataP_npc_6_port, DataP_npc_7_port, 
      DataP_npc_8_port, DataP_npc_9_port, DataP_npc_10_port, DataP_npc_11_port,
      DataP_npc_12_port, DataP_npc_13_port, DataP_npc_14_port, 
      DataP_npc_15_port, DataP_npc_16_port, DataP_npc_17_port, 
      DataP_npc_18_port, DataP_npc_19_port, DataP_npc_20_port, 
      DataP_npc_21_port, DataP_npc_22_port, DataP_npc_23_port, 
      DataP_npc_24_port, DataP_npc_25_port, DataP_npc_26_port, 
      DataP_npc_27_port, DataP_npc_28_port, DataP_npc_29_port, 
      DataP_npc_30_port, DataP_npc_31_port, DataP_IR1_11_port, 
      DataP_IR1_12_port, DataP_IR1_13_port, DataP_IR1_14_port, 
      DataP_IR1_15_port, DataP_IR1_21_port, DataP_IR1_22_port, 
      DataP_IR1_23_port, DataP_IR1_24_port, DataP_IR1_25_port, DataP_PC_reg_N33
      , DataP_PC_reg_N32, DataP_PC_reg_N31, DataP_PC_reg_N30, DataP_PC_reg_N29,
      DataP_PC_reg_N28, DataP_PC_reg_N27, DataP_PC_reg_N26, DataP_PC_reg_N25, 
      DataP_PC_reg_N24, DataP_PC_reg_N23, DataP_PC_reg_N22, DataP_PC_reg_N21, 
      DataP_PC_reg_N20, DataP_PC_reg_N19, DataP_PC_reg_N18, DataP_PC_reg_N17, 
      DataP_PC_reg_N16, DataP_PC_reg_N15, DataP_PC_reg_N14, DataP_PC_reg_N13, 
      DataP_PC_reg_N12, DataP_PC_reg_N11, DataP_PC_reg_N10, DataP_PC_reg_N9, 
      DataP_PC_reg_N8, DataP_PC_reg_N7, DataP_PC_reg_N6, DataP_PC_reg_N5, 
      DataP_PC_reg_N4, DataP_PC_reg_N3, DataP_PC_reg_N2, DataP_NPC_add_N32, 
      DataP_NPC_add_N31, DataP_NPC_add_N30, DataP_NPC_add_N29, 
      DataP_NPC_add_N28, DataP_NPC_add_N27, DataP_NPC_add_N26, 
      DataP_NPC_add_N25, DataP_NPC_add_N24, DataP_NPC_add_N23, 
      DataP_NPC_add_N22, DataP_NPC_add_N21, DataP_NPC_add_N20, 
      DataP_NPC_add_N19, DataP_NPC_add_N18, DataP_NPC_add_N17, 
      DataP_NPC_add_N16, DataP_NPC_add_N15, DataP_NPC_add_N14, 
      DataP_NPC_add_N13, DataP_NPC_add_N12, DataP_NPC_add_N11, 
      DataP_NPC_add_N10, DataP_NPC_add_N9, DataP_NPC_add_N8, DataP_NPC_add_N7, 
      DataP_NPC_add_N6, DataP_NPC_add_N5, DataP_NPC_add_N4, DataP_NPC_add_N3, 
      DataP_NPC_add_N2, DataP_NPC_add_N1, DataP_NPC_add_N0, 
      DataP_IF_IDs_net834167, DataP_FORWARDING_BR_N12, DataP_ALU_C_shifter_N107
      , DataP_ALU_C_shifter_N106, DataP_ALU_C_shifter_N105, 
      DataP_ALU_C_shifter_N104, DataP_ALU_C_shifter_N103, 
      DataP_ALU_C_shifter_N102, DataP_ALU_C_shifter_N101, 
      DataP_ALU_C_shifter_N100, DataP_ALU_C_shifter_N99, 
      DataP_ALU_C_shifter_N98, DataP_ALU_C_shifter_N97, DataP_ALU_C_shifter_N96
      , DataP_ALU_C_shifter_N95, DataP_ALU_C_shifter_N94, 
      DataP_ALU_C_shifter_N93, DataP_ALU_C_shifter_N92, DataP_ALU_C_shifter_N89
      , DataP_ALU_C_shifter_N83, DataP_ALU_C_shifter_N82, 
      DataP_ALU_C_shifter_N81, DataP_ALU_C_shifter_N80, DataP_ALU_C_shifter_N79
      , DataP_ALU_C_shifter_N78, DataP_ALU_C_shifter_N77, 
      DataP_ALU_C_shifter_N76, DataP_ALU_C_shifter_N75, DataP_ALU_C_shifter_N74
      , DataP_ALU_C_shifter_N73, DataP_ALU_C_shifter_N72, 
      DataP_ALU_C_shifter_N71, DataP_ALU_C_shifter_N70, DataP_ALU_C_shifter_N69
      , DataP_ALU_C_shifter_N68, DataP_ALU_C_shifter_N67, 
      DataP_ALU_C_shifter_N66, DataP_ALU_C_shifter_N65, DataP_ALU_C_shifter_N64
      , DataP_ALU_C_shifter_N63, DataP_ALU_C_shifter_N62, 
      DataP_ALU_C_shifter_N61, DataP_ALU_C_shifter_N60, DataP_ALU_C_shifter_N51
      , DataP_ALU_C_shifter_N50, DataP_ALU_C_shifter_N49, 
      DataP_ALU_C_shifter_N48, DataP_ALU_C_shifter_N47, DataP_ALU_C_shifter_N46
      , DataP_ALU_C_shifter_N43, DataP_ALU_C_shifter_N42, 
      DataP_ALU_C_shifter_N40, DataP_ALU_C_shifter_N39, DataP_ALU_C_shifter_N38
      , DataP_ALU_C_shifter_N37, DataP_ALU_C_shifter_N36, 
      DataP_ALU_C_shifter_N34, DataP_ALU_C_shifter_N33, DataP_ALU_C_shifter_N32
      , DataP_ALU_C_shifter_N31, DataP_ALU_C_shifter_N30, 
      DataP_ALU_C_shifter_N29, DataP_ALU_C_shifter_N28, DataP_ALU_C_shifter_N19
      , DataP_ALU_C_comp_N24, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
      n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n296, n297, n299, n300, n301, n303, n304, n308, n309, n311, n313, 
      n317, n319, n322, n323, n326, n330, n332, n333, n337, n340, n341, n345, 
      n350, n353, n354, n355, n356, n357, n358, n399, n432, n443, n476, n477, 
      n478, n479, n480, n482, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n497, n504, n510, n514, n515, n516, n520, n521, n523, 
      n524, n528, n529, n530, n536, n538, n540, n606, n1357, n1371, n1448, 
      n1513, sra_131_SH_4_port, sra_131_SH_1_port, lt_x_135_B_4_port, 
      lt_x_134_B_5_port, lt_x_134_B_4_port, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
      n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
      n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
      n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
      n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
      n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
      n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
      n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
      n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
      n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
      n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
      n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
      n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
      n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
      n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
      n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
      n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
      n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
      n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
      n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
      n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
      n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
      n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, 
      n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
      n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
      n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
      n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
      n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, 
      n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
      n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, 
      n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, 
      n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, 
      n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, 
      n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, 
      n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
      n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
      n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
      n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
      n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
      n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, 
      n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, 
      n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, 
      n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
      n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
      n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, 
      n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
      n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
      n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
      n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, 
      n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, 
      n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
      n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
      n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, 
      n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, 
      n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
      n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
      n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
      n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
      n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, 
      n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, 
      n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
      n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, 
      n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
      n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
      n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
      n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
      n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
      n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
      n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
      n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
      n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
      n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
      n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
      n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
      n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, 
      n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
      n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
      n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
      n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
      n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
      n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
      n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
      n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
      n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
      n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
      n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
      n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, 
      n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, 
      n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
      n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
      n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
      n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
      n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
      n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
      n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
      n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
      n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
      n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
      n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
      n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
      n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
      n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
      n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
      n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
      n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
      n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
      n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
      n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
      n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
      n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
      n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
      n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
      n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
      n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
      n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, 
      n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
      n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
      n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
      n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
      n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
      n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
      n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
      n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, 
      n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
      n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
      n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
      n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, 
      n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, 
      n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
      n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
      n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
      n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, 
      n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
      n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, 
      n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, 
      n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, 
      n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, 
      n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, 
      n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, 
      n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, 
      n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, 
      n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, 
      n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, 
      n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, 
      n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, 
      n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, 
      n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, 
      n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, 
      n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
      n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, 
      n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, 
      n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, 
      n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
      n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
      n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, 
      n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, 
      n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, 
      n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, 
      n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, 
      n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, 
      n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, 
      n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, 
      n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
      n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, 
      n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, 
      n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, 
      n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, 
      n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, 
      n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, 
      n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, 
      n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, 
      n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, 
      n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, 
      n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, 
      n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, 
      n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, 
      n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, 
      n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
      n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
      n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
      n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
      n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, 
      n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, 
      n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, 
      n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, 
      n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, 
      n4020, n4021, n4022, n4023, n4024, n_1004, n_1005, n_1006, n_1007, n_1008
      , n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017,
      n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, 
      n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, 
      n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, 
      n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, 
      n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, 
      n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, 
      n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, 
      n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, 
      n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, 
      n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, 
      n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, 
      n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, 
      n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, 
      n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, 
      n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, 
      n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, 
      n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, 
      n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, 
      n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, 
      n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, 
      n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, 
      n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, 
      n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, 
      n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, 
      n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, 
      n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, 
      n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, 
      n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, 
      n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, 
      n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, 
      n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, 
      n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, 
      n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, 
      n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, 
      n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, 
      n_1396, n_1397 : std_logic;

begin
   DRAM_ADDRESS <= ( DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, 
      DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, 
      DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, 
      DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, 
      DRAM_ADDRESS_0_port );
   IRAM_ADDRESS <= ( IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   
   DataP_Reg_F : register_file_N32_addBit5 port map( RESET => Rst, RE => n1513,
                           WE => RF_WE_i, ADD_WR(4) => DataP_add_D_4_port, 
                           ADD_WR(3) => DataP_add_D_3_port, ADD_WR(2) => n1955,
                           ADD_WR(1) => n1892, ADD_WR(0) => n1852, ADD_RDA(4) 
                           => n494, ADD_RDA(3) => n493, ADD_RDA(2) => n492, 
                           ADD_RDA(1) => n491, ADD_RDA(0) => n490, ADD_RDB(4) 
                           => DataP_add_S2_4_port, ADD_RDB(3) => 
                           DataP_add_S2_3_port, ADD_RDB(2) => 
                           DataP_add_S2_2_port, ADD_RDB(1) => 
                           DataP_add_S2_1_port, ADD_RDB(0) => 
                           DataP_add_S2_0_port, DATAIN(31) => DataP_WB_31_port,
                           DATAIN(30) => DataP_WB_30_port, DATAIN(29) => 
                           DataP_WB_29_port, DATAIN(28) => DataP_WB_28_port, 
                           DATAIN(27) => DataP_WB_27_port, DATAIN(26) => 
                           DataP_WB_26_port, DATAIN(25) => DataP_WB_25_port, 
                           DATAIN(24) => DataP_WB_24_port, DATAIN(23) => 
                           DataP_WB_23_port, DATAIN(22) => DataP_WB_22_port, 
                           DATAIN(21) => DataP_WB_21_port, DATAIN(20) => 
                           DataP_WB_20_port, DATAIN(19) => DataP_WB_19_port, 
                           DATAIN(18) => DataP_WB_18_port, DATAIN(17) => 
                           DataP_WB_17_port, DATAIN(16) => DataP_WB_16_port, 
                           DATAIN(15) => DataP_WB_15_port, DATAIN(14) => 
                           DataP_WB_14_port, DATAIN(13) => DataP_WB_13_port, 
                           DATAIN(12) => DataP_WB_12_port, DATAIN(11) => 
                           DataP_WB_11_port, DATAIN(10) => DataP_WB_10_port, 
                           DATAIN(9) => DataP_WB_9_port, DATAIN(8) => 
                           DataP_WB_8_port, DATAIN(7) => DataP_WB_7_port, 
                           DATAIN(6) => DataP_WB_6_port, DATAIN(5) => 
                           DataP_WB_5_port, DATAIN(4) => DataP_WB_4_port, 
                           DATAIN(3) => DataP_WB_3_port, DATAIN(2) => 
                           DataP_WB_2_port, DATAIN(1) => DataP_WB_1_port, 
                           DATAIN(0) => DataP_WB_0_port, OUTA(31) => 
                           DataP_a_out_31_port, OUTA(30) => DataP_a_out_30_port
                           , OUTA(29) => DataP_a_out_29_port, OUTA(28) => 
                           DataP_a_out_28_port, OUTA(27) => DataP_a_out_27_port
                           , OUTA(26) => DataP_a_out_26_port, OUTA(25) => 
                           DataP_a_out_25_port, OUTA(24) => DataP_a_out_24_port
                           , OUTA(23) => DataP_a_out_23_port, OUTA(22) => 
                           DataP_a_out_22_port, OUTA(21) => DataP_a_out_21_port
                           , OUTA(20) => DataP_a_out_20_port, OUTA(19) => 
                           DataP_a_out_19_port, OUTA(18) => DataP_a_out_18_port
                           , OUTA(17) => DataP_a_out_17_port, OUTA(16) => 
                           DataP_a_out_16_port, OUTA(15) => DataP_a_out_15_port
                           , OUTA(14) => DataP_a_out_14_port, OUTA(13) => 
                           DataP_a_out_13_port, OUTA(12) => DataP_a_out_12_port
                           , OUTA(11) => DataP_a_out_11_port, OUTA(10) => 
                           DataP_a_out_10_port, OUTA(9) => DataP_a_out_9_port, 
                           OUTA(8) => DataP_a_out_8_port, OUTA(7) => 
                           DataP_a_out_7_port, OUTA(6) => DataP_a_out_6_port, 
                           OUTA(5) => DataP_a_out_5_port, OUTA(4) => 
                           DataP_a_out_4_port, OUTA(3) => DataP_a_out_3_port, 
                           OUTA(2) => DataP_a_out_2_port, OUTA(1) => 
                           DataP_a_out_1_port, OUTA(0) => DataP_a_out_0_port, 
                           OUTB(31) => DataP_b_out_31_port, OUTB(30) => 
                           DataP_b_out_30_port, OUTB(29) => DataP_b_out_29_port
                           , OUTB(28) => DataP_b_out_28_port, OUTB(27) => 
                           DataP_b_out_27_port, OUTB(26) => DataP_b_out_26_port
                           , OUTB(25) => DataP_b_out_25_port, OUTB(24) => 
                           DataP_b_out_24_port, OUTB(23) => DataP_b_out_23_port
                           , OUTB(22) => DataP_b_out_22_port, OUTB(21) => 
                           DataP_b_out_21_port, OUTB(20) => DataP_b_out_20_port
                           , OUTB(19) => DataP_b_out_19_port, OUTB(18) => 
                           DataP_b_out_18_port, OUTB(17) => DataP_b_out_17_port
                           , OUTB(16) => DataP_b_out_16_port, OUTB(15) => 
                           DataP_b_out_15_port, OUTB(14) => DataP_b_out_14_port
                           , OUTB(13) => DataP_b_out_13_port, OUTB(12) => 
                           DataP_b_out_12_port, OUTB(11) => DataP_b_out_11_port
                           , OUTB(10) => DataP_b_out_10_port, OUTB(9) => 
                           DataP_b_out_9_port, OUTB(8) => DataP_b_out_8_port, 
                           OUTB(7) => DataP_b_out_7_port, OUTB(6) => 
                           DataP_b_out_6_port, OUTB(5) => DataP_b_out_5_port, 
                           OUTB(4) => DataP_b_out_4_port, OUTB(3) => 
                           DataP_b_out_3_port, OUTB(2) => DataP_b_out_2_port, 
                           OUTB(1) => DataP_b_out_1_port, OUTB(0) => 
                           DataP_b_out_0_port);
   DataP_BR_pred : branch_predictor port map( RST => Rst, PC_IN(31) => 
                           DataP_pc_out_31_port, PC_IN(30) => 
                           DataP_pc_out_30_port, PC_IN(29) => 
                           DataP_pc_out_29_port, PC_IN(28) => 
                           DataP_pc_out_28_port, PC_IN(27) => 
                           DataP_pc_out_27_port, PC_IN(26) => 
                           DataP_pc_out_26_port, PC_IN(25) => 
                           DataP_pc_out_25_port, PC_IN(24) => 
                           DataP_pc_out_24_port, PC_IN(23) => 
                           DataP_pc_out_23_port, PC_IN(22) => 
                           DataP_pc_out_22_port, PC_IN(21) => 
                           DataP_pc_out_21_port, PC_IN(20) => 
                           DataP_pc_out_20_port, PC_IN(19) => 
                           DataP_pc_out_19_port, PC_IN(18) => 
                           DataP_pc_out_18_port, PC_IN(17) => 
                           DataP_pc_out_17_port, PC_IN(16) => 
                           DataP_pc_out_16_port, PC_IN(15) => 
                           DataP_pc_out_15_port, PC_IN(14) => 
                           DataP_pc_out_14_port, PC_IN(13) => 
                           DataP_pc_out_13_port, PC_IN(12) => 
                           DataP_pc_out_12_port, PC_IN(11) => 
                           DataP_pc_out_11_port, PC_IN(10) => 
                           DataP_pc_out_10_port, PC_IN(9) => 
                           IRAM_ADDRESS_7_port, PC_IN(8) => IRAM_ADDRESS_6_port
                           , PC_IN(7) => IRAM_ADDRESS_5_port, PC_IN(6) => 
                           IRAM_ADDRESS_4_port, PC_IN(5) => IRAM_ADDRESS_3_port
                           , PC_IN(4) => IRAM_ADDRESS_2_port, PC_IN(3) => 
                           IRAM_ADDRESS_1_port, PC_IN(2) => IRAM_ADDRESS_0_port
                           , PC_IN(1) => DataP_pc_out_1, PC_IN(0) => 
                           DataP_pc_out_0, PC_FAIL(31) => DataP_npc_M_31_port, 
                           PC_FAIL(30) => DataP_npc_M_30_port, PC_FAIL(29) => 
                           DataP_npc_M_29_port, PC_FAIL(28) => 
                           DataP_npc_M_28_port, PC_FAIL(27) => 
                           DataP_npc_M_27_port, PC_FAIL(26) => 
                           DataP_npc_M_26_port, PC_FAIL(25) => 
                           DataP_npc_M_25_port, PC_FAIL(24) => 
                           DataP_npc_M_24_port, PC_FAIL(23) => 
                           DataP_npc_M_23_port, PC_FAIL(22) => 
                           DataP_npc_M_22_port, PC_FAIL(21) => 
                           DataP_npc_M_21_port, PC_FAIL(20) => 
                           DataP_npc_M_20_port, PC_FAIL(19) => 
                           DataP_npc_M_19_port, PC_FAIL(18) => 
                           DataP_npc_M_18_port, PC_FAIL(17) => 
                           DataP_npc_M_17_port, PC_FAIL(16) => 
                           DataP_npc_M_16_port, PC_FAIL(15) => 
                           DataP_npc_M_15_port, PC_FAIL(14) => 
                           DataP_npc_M_14_port, PC_FAIL(13) => 
                           DataP_npc_M_13_port, PC_FAIL(12) => 
                           DataP_npc_M_12_port, PC_FAIL(11) => 
                           DataP_npc_M_11_port, PC_FAIL(10) => 
                           DataP_npc_M_10_port, PC_FAIL(9) => 
                           DataP_npc_M_9_port, PC_FAIL(8) => DataP_npc_M_8_port
                           , PC_FAIL(7) => DataP_npc_M_7_port, PC_FAIL(6) => 
                           DataP_npc_M_6_port, PC_FAIL(5) => DataP_npc_M_5_port
                           , PC_FAIL(4) => DataP_npc_M_4_port, PC_FAIL(3) => 
                           DataP_npc_M_3_port, PC_FAIL(2) => DataP_npc_M_2_port
                           , PC_FAIL(1) => DataP_npc_M_1_port, PC_FAIL(0) => 
                           DataP_npc_M_0_port, IR_IN(31) => IRAM_DATA_OUT(31), 
                           IR_IN(30) => IRAM_DATA_OUT(30), IR_IN(29) => 
                           IRAM_DATA_OUT(29), IR_IN(28) => IRAM_DATA_OUT(28), 
                           IR_IN(27) => IRAM_DATA_OUT(27), IR_IN(26) => n4024, 
                           IR_IN(25) => IRAM_DATA_OUT(25), IR_IN(24) => 
                           IRAM_DATA_OUT(24), IR_IN(23) => IRAM_DATA_OUT(23), 
                           IR_IN(22) => IRAM_DATA_OUT(22), IR_IN(21) => 
                           IRAM_DATA_OUT(21), IR_IN(20) => IRAM_DATA_OUT(20), 
                           IR_IN(19) => IRAM_DATA_OUT(19), IR_IN(18) => 
                           IRAM_DATA_OUT(18), IR_IN(17) => IRAM_DATA_OUT(17), 
                           IR_IN(16) => IRAM_DATA_OUT(16), IR_IN(15) => 
                           IRAM_DATA_OUT(15), IR_IN(14) => IRAM_DATA_OUT(14), 
                           IR_IN(13) => IRAM_DATA_OUT(13), IR_IN(12) => 
                           IRAM_DATA_OUT(12), IR_IN(11) => IRAM_DATA_OUT(11), 
                           IR_IN(10) => IRAM_DATA_OUT(10), IR_IN(9) => 
                           IRAM_DATA_OUT(9), IR_IN(8) => IRAM_DATA_OUT(8), 
                           IR_IN(7) => IRAM_DATA_OUT(7), IR_IN(6) => 
                           IRAM_DATA_OUT(6), IR_IN(5) => IRAM_DATA_OUT(5), 
                           IR_IN(4) => IRAM_DATA_OUT(4), IR_IN(3) => 
                           IRAM_DATA_OUT(3), IR_IN(2) => IRAM_DATA_OUT(2), 
                           IR_IN(1) => IRAM_DATA_OUT(1), IR_IN(0) => 
                           IRAM_DATA_OUT(0), IR_FAIL(15) => DataP_ir_E_15_port,
                           IR_FAIL(14) => DataP_ir_E_14_port, IR_FAIL(13) => 
                           DataP_ir_E_13_port, IR_FAIL(12) => 
                           DataP_ir_E_12_port, IR_FAIL(11) => 
                           DataP_ir_E_11_port, IR_FAIL(10) => 
                           DataP_ir_E_10_port, IR_FAIL(9) => DataP_ir_E_9_port,
                           IR_FAIL(8) => DataP_ir_E_8_port, IR_FAIL(7) => 
                           DataP_ir_E_7_port, IR_FAIL(6) => DataP_ir_E_6_port, 
                           IR_FAIL(5) => DataP_ir_E_5_port, IR_FAIL(4) => 
                           DataP_ir_E_4_port, IR_FAIL(3) => DataP_ir_E_3_port, 
                           IR_FAIL(2) => DataP_ir_E_2_port, IR_FAIL(1) => 
                           DataP_ir_E_1_port, IR_FAIL(0) => DataP_ir_E_0_port, 
                           WRONG_PRE => DataP_wrong_br, RIGHT_PRE => 
                           DataP_right_br, NPC_OUT(31) => DataP_npc_pre_31_port
                           , NPC_OUT(30) => DataP_npc_pre_30_port, NPC_OUT(29) 
                           => DataP_npc_pre_29_port, NPC_OUT(28) => 
                           DataP_npc_pre_28_port, NPC_OUT(27) => 
                           DataP_npc_pre_27_port, NPC_OUT(26) => 
                           DataP_npc_pre_26_port, NPC_OUT(25) => 
                           DataP_npc_pre_25_port, NPC_OUT(24) => 
                           DataP_npc_pre_24_port, NPC_OUT(23) => 
                           DataP_npc_pre_23_port, NPC_OUT(22) => 
                           DataP_npc_pre_22_port, NPC_OUT(21) => 
                           DataP_npc_pre_21_port, NPC_OUT(20) => 
                           DataP_npc_pre_20_port, NPC_OUT(19) => 
                           DataP_npc_pre_19_port, NPC_OUT(18) => 
                           DataP_npc_pre_18_port, NPC_OUT(17) => 
                           DataP_npc_pre_17_port, NPC_OUT(16) => 
                           DataP_npc_pre_16_port, NPC_OUT(15) => 
                           DataP_npc_pre_15_port, NPC_OUT(14) => 
                           DataP_npc_pre_14_port, NPC_OUT(13) => 
                           DataP_npc_pre_13_port, NPC_OUT(12) => 
                           DataP_npc_pre_12_port, NPC_OUT(11) => 
                           DataP_npc_pre_11_port, NPC_OUT(10) => 
                           DataP_npc_pre_10_port, NPC_OUT(9) => 
                           DataP_npc_pre_9_port, NPC_OUT(8) => 
                           DataP_npc_pre_8_port, NPC_OUT(7) => 
                           DataP_npc_pre_7_port, NPC_OUT(6) => 
                           DataP_npc_pre_6_port, NPC_OUT(5) => 
                           DataP_npc_pre_5_port, NPC_OUT(4) => 
                           DataP_npc_pre_4_port, NPC_OUT(3) => 
                           DataP_npc_pre_3_port, NPC_OUT(2) => 
                           DataP_npc_pre_2_port, NPC_OUT(1) => 
                           DataP_npc_pre_1_port, NPC_OUT(0) => 
                           DataP_npc_pre_0_port, LINK_ADD(31) => 
                           DataP_link_addr_F_31_port, LINK_ADD(30) => 
                           DataP_link_addr_F_30_port, LINK_ADD(29) => 
                           DataP_link_addr_F_29_port, LINK_ADD(28) => 
                           DataP_link_addr_F_28_port, LINK_ADD(27) => 
                           DataP_link_addr_F_27_port, LINK_ADD(26) => 
                           DataP_link_addr_F_26_port, LINK_ADD(25) => 
                           DataP_link_addr_F_25_port, LINK_ADD(24) => 
                           DataP_link_addr_F_24_port, LINK_ADD(23) => 
                           DataP_link_addr_F_23_port, LINK_ADD(22) => 
                           DataP_link_addr_F_22_port, LINK_ADD(21) => 
                           DataP_link_addr_F_21_port, LINK_ADD(20) => 
                           DataP_link_addr_F_20_port, LINK_ADD(19) => 
                           DataP_link_addr_F_19_port, LINK_ADD(18) => 
                           DataP_link_addr_F_18_port, LINK_ADD(17) => 
                           DataP_link_addr_F_17_port, LINK_ADD(16) => 
                           DataP_link_addr_F_16_port, LINK_ADD(15) => 
                           DataP_link_addr_F_15_port, LINK_ADD(14) => 
                           DataP_link_addr_F_14_port, LINK_ADD(13) => 
                           DataP_link_addr_F_13_port, LINK_ADD(12) => 
                           DataP_link_addr_F_12_port, LINK_ADD(11) => 
                           DataP_link_addr_F_11_port, LINK_ADD(10) => 
                           DataP_link_addr_F_10_port, LINK_ADD(9) => 
                           DataP_link_addr_F_9_port, LINK_ADD(8) => 
                           DataP_link_addr_F_8_port, LINK_ADD(7) => 
                           DataP_link_addr_F_7_port, LINK_ADD(6) => 
                           DataP_link_addr_F_6_port, LINK_ADD(5) => 
                           DataP_link_addr_F_5_port, LINK_ADD(4) => 
                           DataP_link_addr_F_4_port, LINK_ADD(3) => 
                           DataP_link_addr_F_3_port, LINK_ADD(2) => 
                           DataP_link_addr_F_2_port, LINK_ADD(1) => 
                           DataP_link_addr_F_1_port, LINK_ADD(0) => 
                           DataP_link_addr_F_0_port, SEL => DataP_npc_mux_sel, 
                           TAKEN => DataP_prediction);
   DataP_IF_IDs_clk_gate_PR_OUT_reg : SNPS_CLOCK_GATE_HIGH_IF_ID port map( CLK 
                           => Clk, EN => n1448, ENCLK => DataP_IF_IDs_net834167
                           , TE => n4024);
   DataP_NPC_add_outPC_reg_0_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N1, Q => DataP_npc_0_port);
   DataP_NPC_add_outPC_reg_1_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N2, Q => DataP_npc_1_port);
   DataP_NPC_add_outPC_reg_2_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N3, Q => DataP_npc_2_port);
   DataP_NPC_add_outPC_reg_3_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N4, Q => DataP_npc_3_port);
   DataP_NPC_add_outPC_reg_4_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N5, Q => DataP_npc_4_port);
   DataP_NPC_add_outPC_reg_5_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N6, Q => DataP_npc_5_port);
   DataP_NPC_add_outPC_reg_6_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N7, Q => DataP_npc_6_port);
   DataP_NPC_add_outPC_reg_7_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N8, Q => DataP_npc_7_port);
   DataP_NPC_add_outPC_reg_8_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N9, Q => DataP_npc_8_port);
   DataP_NPC_add_outPC_reg_9_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N10, Q => DataP_npc_9_port);
   DataP_NPC_add_outPC_reg_10_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N11, Q => DataP_npc_10_port);
   DataP_NPC_add_outPC_reg_11_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N12, Q => DataP_npc_11_port);
   DataP_NPC_add_outPC_reg_12_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N13, Q => DataP_npc_12_port);
   DataP_NPC_add_outPC_reg_13_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N14, Q => DataP_npc_13_port);
   DataP_NPC_add_outPC_reg_14_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N15, Q => DataP_npc_14_port);
   DataP_NPC_add_outPC_reg_15_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N16, Q => DataP_npc_15_port);
   DataP_NPC_add_outPC_reg_16_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N17, Q => DataP_npc_16_port);
   DataP_NPC_add_outPC_reg_17_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N18, Q => DataP_npc_17_port);
   DataP_NPC_add_outPC_reg_18_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N19, Q => DataP_npc_18_port);
   DataP_NPC_add_outPC_reg_19_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N20, Q => DataP_npc_19_port);
   DataP_NPC_add_outPC_reg_20_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N21, Q => DataP_npc_20_port);
   DataP_NPC_add_outPC_reg_21_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N22, Q => DataP_npc_21_port);
   DataP_NPC_add_outPC_reg_22_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N23, Q => DataP_npc_22_port);
   DataP_NPC_add_outPC_reg_23_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N24, Q => DataP_npc_23_port);
   DataP_NPC_add_outPC_reg_24_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N25, Q => DataP_npc_24_port);
   DataP_NPC_add_outPC_reg_25_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N26, Q => DataP_npc_25_port);
   DataP_NPC_add_outPC_reg_26_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N27, Q => DataP_npc_26_port);
   DataP_NPC_add_outPC_reg_27_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N28, Q => DataP_npc_27_port);
   DataP_NPC_add_outPC_reg_28_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N29, Q => DataP_npc_28_port);
   DataP_NPC_add_outPC_reg_29_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N30, Q => DataP_npc_29_port);
   DataP_NPC_add_outPC_reg_30_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N31, Q => DataP_npc_30_port);
   DataP_NPC_add_outPC_reg_31_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N32, Q => DataP_npc_31_port);
   DataP_MEM_WB_s_LMD_OUT_reg_0_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(0),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_0_port, QN 
                           => n_1004);
   DataP_MEM_WB_s_LMD_OUT_reg_1_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(1),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_1_port, QN 
                           => n_1005);
   DataP_MEM_WB_s_LMD_OUT_reg_2_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(2),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_2_port, QN 
                           => n_1006);
   DataP_MEM_WB_s_LMD_OUT_reg_3_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(3),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_3_port, QN 
                           => n_1007);
   DataP_MEM_WB_s_LMD_OUT_reg_4_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(4),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_4_port, QN 
                           => n_1008);
   DataP_MEM_WB_s_LMD_OUT_reg_5_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(5),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_5_port, QN 
                           => n_1009);
   DataP_MEM_WB_s_LMD_OUT_reg_6_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(6),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_6_port, QN 
                           => n_1010);
   DataP_MEM_WB_s_LMD_OUT_reg_7_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(7),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_7_port, QN 
                           => n_1011);
   DataP_MEM_WB_s_LMD_OUT_reg_8_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(8),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_8_port, QN 
                           => n_1012);
   DataP_MEM_WB_s_LMD_OUT_reg_9_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(9),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_9_port, QN 
                           => n_1013);
   DataP_MEM_WB_s_LMD_OUT_reg_10_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(10), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_10_port, QN => n_1014);
   DataP_MEM_WB_s_LMD_OUT_reg_11_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(11), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_11_port, QN => n_1015);
   DataP_MEM_WB_s_LMD_OUT_reg_12_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(12), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_12_port, QN => n_1016);
   DataP_MEM_WB_s_LMD_OUT_reg_13_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(13), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_13_port, QN => n_1017);
   DataP_MEM_WB_s_LMD_OUT_reg_14_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(14), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_14_port, QN => n_1018);
   DataP_MEM_WB_s_LMD_OUT_reg_15_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(15), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_15_port, QN => n_1019);
   DataP_MEM_WB_s_LMD_OUT_reg_16_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(16), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_16_port, QN => n_1020);
   DataP_MEM_WB_s_LMD_OUT_reg_17_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(17), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_17_port, QN => n_1021);
   DataP_MEM_WB_s_LMD_OUT_reg_18_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(18), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_18_port, QN => n_1022);
   DataP_MEM_WB_s_LMD_OUT_reg_19_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(19), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_19_port, QN => n_1023);
   DataP_MEM_WB_s_LMD_OUT_reg_20_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(20), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_20_port, QN => n_1024);
   DataP_MEM_WB_s_LMD_OUT_reg_21_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(21), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_21_port, QN => n_1025);
   DataP_MEM_WB_s_LMD_OUT_reg_22_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(22), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_22_port, QN => n_1026);
   DataP_MEM_WB_s_LMD_OUT_reg_23_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(23), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_23_port, QN => n_1027);
   DataP_MEM_WB_s_LMD_OUT_reg_24_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(24), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_24_port, QN => n_1028);
   DataP_MEM_WB_s_LMD_OUT_reg_25_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(25), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_25_port, QN => n_1029);
   DataP_MEM_WB_s_LMD_OUT_reg_26_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(26), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_26_port, QN => n_1030);
   DataP_MEM_WB_s_LMD_OUT_reg_27_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(27), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_27_port, QN => n_1031);
   DataP_MEM_WB_s_LMD_OUT_reg_28_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(28), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_28_port, QN => n_1032);
   DataP_MEM_WB_s_LMD_OUT_reg_29_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(29), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_29_port, QN => n_1033);
   DataP_MEM_WB_s_LMD_OUT_reg_30_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(30), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_30_port, QN => n_1034);
   DataP_MEM_WB_s_LMD_OUT_reg_31_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(31), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_31_port, QN => n_1035);
   DataP_MEM_WB_s_ALU_OUT_reg_31_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_31_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_31_port, QN => n2267);
   DataP_IF_IDs_NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_31_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1036, QN 
                           => n293);
   DataP_ID_EXs_NPC_L_OUT_reg_31_inst : DFFS_X1 port map( D => n293, CK => Clk,
                           SN => Rst, Q => n292, QN => n_1037);
   DataP_EX_MEM_s_NPC_L_OUT_reg_31_inst : DFFS_X1 port map( D => n292, CK => 
                           Clk, SN => Rst, Q => n291, QN => n_1038);
   DataP_MEM_WB_s_NPC_L_OUT_reg_31_inst : DFFS_X1 port map( D => n291, CK => 
                           Clk, SN => Rst, Q => n_1039, QN => 
                           DataP_link_addr_W_31_port);
   DataP_ID_EXs_B_OUT_reg_0_inst : DFFR_X1 port map( D => DataP_b_out_0_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_0_port, QN => 
                           n290);
   DataP_EX_MEM_s_B_OUT_reg_0_inst : DFFS_X1 port map( D => n290, CK => Clk, SN
                           => Rst, Q => n_1040, QN => DRAM_DATA_IN(0));
   DataP_ID_EXs_B_OUT_reg_1_inst : DFFR_X1 port map( D => DataP_b_out_1_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_1_port, QN => 
                           n289);
   DataP_EX_MEM_s_B_OUT_reg_1_inst : DFFS_X1 port map( D => n289, CK => Clk, SN
                           => Rst, Q => n_1041, QN => DRAM_DATA_IN(1));
   DataP_ID_EXs_B_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_b_out_2_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_2_port, QN => 
                           n288);
   DataP_EX_MEM_s_B_OUT_reg_2_inst : DFFS_X1 port map( D => n288, CK => Clk, SN
                           => Rst, Q => n_1042, QN => DRAM_DATA_IN(2));
   DataP_ID_EXs_B_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_b_out_3_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_3_port, QN => 
                           n287);
   DataP_EX_MEM_s_B_OUT_reg_3_inst : DFFS_X1 port map( D => n287, CK => Clk, SN
                           => Rst, Q => n_1043, QN => DRAM_DATA_IN(3));
   DataP_ID_EXs_B_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_b_out_4_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_4_port, QN => 
                           n286);
   DataP_EX_MEM_s_B_OUT_reg_4_inst : DFFS_X1 port map( D => n286, CK => Clk, SN
                           => Rst, Q => n_1044, QN => DRAM_DATA_IN(4));
   DataP_ID_EXs_B_OUT_reg_5_inst : DFFR_X1 port map( D => DataP_b_out_5_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_5_port, QN => 
                           n285);
   DataP_EX_MEM_s_B_OUT_reg_5_inst : DFFS_X1 port map( D => n285, CK => Clk, SN
                           => Rst, Q => n_1045, QN => DRAM_DATA_IN(5));
   DataP_ID_EXs_B_OUT_reg_6_inst : DFFR_X1 port map( D => DataP_b_out_6_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_6_port, QN => 
                           n284);
   DataP_EX_MEM_s_B_OUT_reg_6_inst : DFFS_X1 port map( D => n284, CK => Clk, SN
                           => Rst, Q => n_1046, QN => DRAM_DATA_IN(6));
   DataP_ID_EXs_B_OUT_reg_7_inst : DFFR_X1 port map( D => DataP_b_out_7_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_7_port, QN => 
                           n283);
   DataP_EX_MEM_s_B_OUT_reg_7_inst : DFFS_X1 port map( D => n283, CK => Clk, SN
                           => Rst, Q => n_1047, QN => DRAM_DATA_IN(7));
   DataP_ID_EXs_B_OUT_reg_8_inst : DFFR_X1 port map( D => DataP_b_out_8_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_8_port, QN => 
                           n282);
   DataP_EX_MEM_s_B_OUT_reg_8_inst : DFFS_X1 port map( D => n282, CK => Clk, SN
                           => Rst, Q => n_1048, QN => DRAM_DATA_IN(8));
   DataP_ID_EXs_B_OUT_reg_9_inst : DFFR_X1 port map( D => DataP_b_out_9_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_9_port, QN => 
                           n281);
   DataP_EX_MEM_s_B_OUT_reg_9_inst : DFFS_X1 port map( D => n281, CK => Clk, SN
                           => Rst, Q => n_1049, QN => DRAM_DATA_IN(9));
   DataP_ID_EXs_B_OUT_reg_10_inst : DFFR_X1 port map( D => DataP_b_out_10_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_10_port, QN => 
                           n280);
   DataP_EX_MEM_s_B_OUT_reg_10_inst : DFFS_X1 port map( D => n280, CK => Clk, 
                           SN => Rst, Q => n_1050, QN => DRAM_DATA_IN(10));
   DataP_ID_EXs_B_OUT_reg_11_inst : DFFR_X1 port map( D => DataP_b_out_11_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_11_port, QN => 
                           n279);
   DataP_EX_MEM_s_B_OUT_reg_11_inst : DFFS_X1 port map( D => n279, CK => Clk, 
                           SN => Rst, Q => n_1051, QN => DRAM_DATA_IN(11));
   DataP_ID_EXs_B_OUT_reg_12_inst : DFFR_X1 port map( D => DataP_b_out_12_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_12_port, QN => 
                           n278);
   DataP_EX_MEM_s_B_OUT_reg_12_inst : DFFS_X1 port map( D => n278, CK => Clk, 
                           SN => Rst, Q => n_1052, QN => DRAM_DATA_IN(12));
   DataP_ID_EXs_B_OUT_reg_13_inst : DFFR_X1 port map( D => DataP_b_out_13_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_13_port, QN => 
                           n277);
   DataP_EX_MEM_s_B_OUT_reg_13_inst : DFFS_X1 port map( D => n277, CK => Clk, 
                           SN => Rst, Q => n_1053, QN => DRAM_DATA_IN(13));
   DataP_ID_EXs_B_OUT_reg_14_inst : DFFR_X1 port map( D => DataP_b_out_14_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_14_port, QN => 
                           n276);
   DataP_EX_MEM_s_B_OUT_reg_14_inst : DFFS_X1 port map( D => n276, CK => Clk, 
                           SN => Rst, Q => n_1054, QN => DRAM_DATA_IN(14));
   DataP_ID_EXs_B_OUT_reg_15_inst : DFFR_X1 port map( D => DataP_b_out_15_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_15_port, QN => 
                           n275);
   DataP_EX_MEM_s_B_OUT_reg_15_inst : DFFS_X1 port map( D => n275, CK => Clk, 
                           SN => Rst, Q => n_1055, QN => DRAM_DATA_IN(15));
   DataP_ID_EXs_B_OUT_reg_16_inst : DFFR_X1 port map( D => DataP_b_out_16_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_16_port, QN => 
                           n274);
   DataP_EX_MEM_s_B_OUT_reg_16_inst : DFFS_X1 port map( D => n274, CK => Clk, 
                           SN => Rst, Q => n_1056, QN => DRAM_DATA_IN(16));
   DataP_ID_EXs_B_OUT_reg_17_inst : DFFR_X1 port map( D => DataP_b_out_17_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_17_port, QN => 
                           n273);
   DataP_EX_MEM_s_B_OUT_reg_17_inst : DFFS_X1 port map( D => n273, CK => Clk, 
                           SN => Rst, Q => n_1057, QN => DRAM_DATA_IN(17));
   DataP_ID_EXs_B_OUT_reg_18_inst : DFFR_X1 port map( D => DataP_b_out_18_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_18_port, QN => 
                           n272);
   DataP_EX_MEM_s_B_OUT_reg_18_inst : DFFS_X1 port map( D => n272, CK => Clk, 
                           SN => Rst, Q => n_1058, QN => DRAM_DATA_IN(18));
   DataP_ID_EXs_B_OUT_reg_19_inst : DFFR_X1 port map( D => DataP_b_out_19_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_19_port, QN => 
                           n271);
   DataP_EX_MEM_s_B_OUT_reg_19_inst : DFFS_X1 port map( D => n271, CK => Clk, 
                           SN => Rst, Q => n_1059, QN => DRAM_DATA_IN(19));
   DataP_ID_EXs_B_OUT_reg_20_inst : DFFR_X1 port map( D => DataP_b_out_20_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_20_port, QN => 
                           n270);
   DataP_EX_MEM_s_B_OUT_reg_20_inst : DFFS_X1 port map( D => n270, CK => Clk, 
                           SN => Rst, Q => n_1060, QN => DRAM_DATA_IN(20));
   DataP_ID_EXs_B_OUT_reg_21_inst : DFFR_X1 port map( D => DataP_b_out_21_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_21_port, QN => 
                           n269);
   DataP_EX_MEM_s_B_OUT_reg_21_inst : DFFS_X1 port map( D => n269, CK => Clk, 
                           SN => Rst, Q => n_1061, QN => DRAM_DATA_IN(21));
   DataP_ID_EXs_B_OUT_reg_22_inst : DFFR_X1 port map( D => DataP_b_out_22_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_22_port, QN => 
                           n268);
   DataP_EX_MEM_s_B_OUT_reg_22_inst : DFFS_X1 port map( D => n268, CK => Clk, 
                           SN => Rst, Q => n_1062, QN => DRAM_DATA_IN(22));
   DataP_ID_EXs_B_OUT_reg_23_inst : DFFR_X1 port map( D => DataP_b_out_23_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_23_port, QN => 
                           n267);
   DataP_EX_MEM_s_B_OUT_reg_23_inst : DFFS_X1 port map( D => n267, CK => Clk, 
                           SN => Rst, Q => n_1063, QN => DRAM_DATA_IN(23));
   DataP_ID_EXs_B_OUT_reg_24_inst : DFFR_X1 port map( D => DataP_b_out_24_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_24_port, QN => 
                           n266);
   DataP_EX_MEM_s_B_OUT_reg_24_inst : DFFS_X1 port map( D => n266, CK => Clk, 
                           SN => Rst, Q => n_1064, QN => DRAM_DATA_IN(24));
   DataP_ID_EXs_B_OUT_reg_25_inst : DFFR_X1 port map( D => DataP_b_out_25_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_25_port, QN => 
                           n265);
   DataP_EX_MEM_s_B_OUT_reg_25_inst : DFFS_X1 port map( D => n265, CK => Clk, 
                           SN => Rst, Q => n_1065, QN => DRAM_DATA_IN(25));
   DataP_ID_EXs_B_OUT_reg_26_inst : DFFR_X1 port map( D => DataP_b_out_26_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_26_port, QN => 
                           n264);
   DataP_EX_MEM_s_B_OUT_reg_26_inst : DFFS_X1 port map( D => n264, CK => Clk, 
                           SN => Rst, Q => n_1066, QN => DRAM_DATA_IN(26));
   DataP_ID_EXs_B_OUT_reg_27_inst : DFFR_X1 port map( D => DataP_b_out_27_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_27_port, QN => 
                           n263);
   DataP_EX_MEM_s_B_OUT_reg_27_inst : DFFS_X1 port map( D => n263, CK => Clk, 
                           SN => Rst, Q => n_1067, QN => DRAM_DATA_IN(27));
   DataP_ID_EXs_B_OUT_reg_28_inst : DFFR_X1 port map( D => DataP_b_out_28_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_28_port, QN => 
                           n262);
   DataP_EX_MEM_s_B_OUT_reg_28_inst : DFFS_X1 port map( D => n262, CK => Clk, 
                           SN => Rst, Q => n_1068, QN => DRAM_DATA_IN(28));
   DataP_ID_EXs_B_OUT_reg_29_inst : DFFR_X1 port map( D => DataP_b_out_29_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_29_port, QN => 
                           n261);
   DataP_EX_MEM_s_B_OUT_reg_29_inst : DFFS_X1 port map( D => n261, CK => Clk, 
                           SN => Rst, Q => n_1069, QN => DRAM_DATA_IN(29));
   DataP_ID_EXs_B_OUT_reg_30_inst : DFFR_X1 port map( D => DataP_b_out_30_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_30_port, QN => 
                           n260);
   DataP_EX_MEM_s_B_OUT_reg_30_inst : DFFS_X1 port map( D => n260, CK => Clk, 
                           SN => Rst, Q => n_1070, QN => DRAM_DATA_IN(30));
   DataP_ID_EXs_B_OUT_reg_31_inst : DFFR_X1 port map( D => DataP_b_out_31_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_31_port, QN => 
                           n259);
   DataP_EX_MEM_s_B_OUT_reg_31_inst : DFFS_X1 port map( D => n259, CK => Clk, 
                           SN => Rst, Q => n_1071, QN => DRAM_DATA_IN(31));
   DataP_ID_EXs_A_OUT_reg_0_inst : DFFR_X1 port map( D => DataP_a_out_0_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_0_port, QN => 
                           n2214);
   DataP_ID_EXs_A_OUT_reg_1_inst : DFFR_X1 port map( D => DataP_a_out_1_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_1_port, QN => 
                           n2215);
   DataP_ID_EXs_A_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_a_out_2_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_2_port, QN => 
                           n2213);
   DataP_ID_EXs_A_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_a_out_3_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_3_port, QN => 
                           n2212);
   DataP_ID_EXs_A_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_a_out_4_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_4_port, QN => 
                           n2221);
   DataP_ID_EXs_A_OUT_reg_5_inst : DFFR_X1 port map( D => DataP_a_out_5_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_5_port, QN => 
                           n2198);
   DataP_ID_EXs_A_OUT_reg_6_inst : DFFR_X1 port map( D => DataP_a_out_6_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_6_port, QN => 
                           n2216);
   DataP_ID_EXs_A_OUT_reg_7_inst : DFFR_X1 port map( D => DataP_a_out_7_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_7_port, QN => 
                           n2205);
   DataP_ID_EXs_A_OUT_reg_8_inst : DFFR_X1 port map( D => DataP_a_out_8_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_8_port, QN => 
                           n2220);
   DataP_ID_EXs_A_OUT_reg_9_inst : DFFR_X1 port map( D => DataP_a_out_9_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_9_port, QN => 
                           n2190);
   DataP_ID_EXs_A_OUT_reg_10_inst : DFFR_X1 port map( D => DataP_a_out_10_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_10_port, QN => 
                           n2211);
   DataP_ID_EXs_A_OUT_reg_11_inst : DFFR_X1 port map( D => DataP_a_out_11_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_11_port, QN => 
                           n2204);
   DataP_ID_EXs_A_OUT_reg_12_inst : DFFR_X1 port map( D => DataP_a_out_12_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_12_port, QN => 
                           n2197);
   DataP_ID_EXs_A_OUT_reg_13_inst : DFFR_X1 port map( D => DataP_a_out_13_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_13_port, QN => 
                           n2210);
   DataP_ID_EXs_A_OUT_reg_14_inst : DFFR_X1 port map( D => DataP_a_out_14_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_14_port, QN => 
                           n2203);
   DataP_ID_EXs_A_OUT_reg_15_inst : DFFR_X1 port map( D => DataP_a_out_15_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_15_port, QN => 
                           n2196);
   DataP_ID_EXs_A_OUT_reg_16_inst : DFFR_X1 port map( D => DataP_a_out_16_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_16_port, QN => 
                           n2219);
   DataP_ID_EXs_A_OUT_reg_17_inst : DFFR_X1 port map( D => DataP_a_out_17_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_17_port, QN => 
                           n2195);
   DataP_ID_EXs_A_OUT_reg_18_inst : DFFR_X1 port map( D => DataP_a_out_18_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_18_port, QN => 
                           n2209);
   DataP_ID_EXs_A_OUT_reg_19_inst : DFFR_X1 port map( D => DataP_a_out_19_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_19_port, QN => 
                           n2202);
   DataP_ID_EXs_A_OUT_reg_20_inst : DFFR_X1 port map( D => DataP_a_out_20_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_20_port, QN => 
                           n2208);
   DataP_ID_EXs_A_OUT_reg_21_inst : DFFR_X1 port map( D => DataP_a_out_21_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_21_port, QN => 
                           n2201);
   DataP_ID_EXs_A_OUT_reg_22_inst : DFFR_X1 port map( D => DataP_a_out_22_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_22_port, QN => 
                           n2218);
   DataP_ID_EXs_A_OUT_reg_23_inst : DFFR_X1 port map( D => DataP_a_out_23_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_23_port, QN => 
                           n2194);
   DataP_ID_EXs_A_OUT_reg_24_inst : DFFR_X1 port map( D => DataP_a_out_24_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_24_port, QN => 
                           n2217);
   DataP_ID_EXs_A_OUT_reg_25_inst : DFFR_X1 port map( D => DataP_a_out_25_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_25_port, QN => 
                           n2207);
   DataP_ID_EXs_A_OUT_reg_26_inst : DFFR_X1 port map( D => DataP_a_out_26_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_26_port, QN => 
                           n2200);
   DataP_ID_EXs_A_OUT_reg_27_inst : DFFR_X1 port map( D => DataP_a_out_27_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_27_port, QN => 
                           n2193);
   DataP_ID_EXs_A_OUT_reg_28_inst : DFFR_X1 port map( D => DataP_a_out_28_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_28_port, QN => 
                           n2206);
   DataP_ID_EXs_A_OUT_reg_29_inst : DFFR_X1 port map( D => DataP_a_out_29_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_29_port, QN => 
                           n2199);
   DataP_ID_EXs_A_OUT_reg_30_inst : DFFR_X1 port map( D => DataP_a_out_30_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_30_port, QN => 
                           n2192);
   DataP_ID_EXs_A_OUT_reg_31_inst : DFFR_X1 port map( D => DataP_a_out_31_port,
                           CK => Clk, RN => Rst, Q => DataP_A_s_31_port, QN => 
                           n2191);
   DataP_EX_MEM_s_ALU_OUT_reg_0_inst : DFFS_X1 port map( D => n296, CK => Clk, 
                           SN => Rst, Q => n2234, QN => DRAM_ADDRESS_0_port);
   DataP_MEM_WB_s_ALU_OUT_reg_0_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_0_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_0_port, QN => n2272);
   DataP_EX_MEM_s_ALU_OUT_reg_7_inst : DFFS_X1 port map( D => n350, CK => Clk, 
                           SN => Rst, Q => n2230, QN => DRAM_ADDRESS_7_port);
   DataP_MEM_WB_s_ALU_OUT_reg_7_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_7_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_7_port, QN => n2275);
   DataP_MEM_WB_s_ALU_OUT_reg_15_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_15_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_15_port, QN => n2247);
   DataP_MEM_WB_s_ALU_OUT_reg_19_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_19_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_19_port, QN => n2253);
   DataP_MEM_WB_s_ALU_OUT_reg_23_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_23_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_23_port, QN => n2249);
   DataP_EX_MEM_s_ALU_OUT_reg_27_inst : DFFS_X1 port map( D => n301, CK => Clk,
                           SN => Rst, Q => n2165, QN => DataP_alu_out_M_27_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_27_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_27_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_27_port, QN => n2250);
   DataP_MEM_WB_s_ALU_OUT_reg_30_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_30_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_30_port, QN => n2266);
   DataP_ID_EXs_PR_OUT_reg : DFFS_X1 port map( D => n258, CK => Clk, SN => Rst,
                           Q => n_1072, QN => DataP_pr_E);
   DataP_IF_IDs_NPC_L_OUT_reg_30_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_30_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1073, QN 
                           => n257);
   DataP_ID_EXs_NPC_L_OUT_reg_30_inst : DFFS_X1 port map( D => n257, CK => Clk,
                           SN => Rst, Q => n256, QN => n_1074);
   DataP_EX_MEM_s_NPC_L_OUT_reg_30_inst : DFFS_X1 port map( D => n256, CK => 
                           Clk, SN => Rst, Q => n255, QN => n_1075);
   DataP_MEM_WB_s_NPC_L_OUT_reg_30_inst : DFFS_X1 port map( D => n255, CK => 
                           Clk, SN => Rst, Q => n_1076, QN => 
                           DataP_link_addr_W_30_port);
   DataP_IF_IDs_NPC_L_OUT_reg_29_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_29_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1077, QN 
                           => n254);
   DataP_ID_EXs_NPC_L_OUT_reg_29_inst : DFFS_X1 port map( D => n254, CK => Clk,
                           SN => Rst, Q => n253, QN => n_1078);
   DataP_EX_MEM_s_NPC_L_OUT_reg_29_inst : DFFS_X1 port map( D => n253, CK => 
                           Clk, SN => Rst, Q => n252, QN => n_1079);
   DataP_MEM_WB_s_NPC_L_OUT_reg_29_inst : DFFS_X1 port map( D => n252, CK => 
                           Clk, SN => Rst, Q => n_1080, QN => 
                           DataP_link_addr_W_29_port);
   DataP_IF_IDs_NPC_L_OUT_reg_28_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_28_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1081, QN 
                           => n251);
   DataP_ID_EXs_NPC_L_OUT_reg_28_inst : DFFS_X1 port map( D => n251, CK => Clk,
                           SN => Rst, Q => n250, QN => n_1082);
   DataP_EX_MEM_s_NPC_L_OUT_reg_28_inst : DFFS_X1 port map( D => n250, CK => 
                           Clk, SN => Rst, Q => n249, QN => n_1083);
   DataP_MEM_WB_s_NPC_L_OUT_reg_28_inst : DFFS_X1 port map( D => n249, CK => 
                           Clk, SN => Rst, Q => n_1084, QN => 
                           DataP_link_addr_W_28_port);
   DataP_IF_IDs_NPC_L_OUT_reg_27_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_27_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1085, QN 
                           => n248);
   DataP_ID_EXs_NPC_L_OUT_reg_27_inst : DFFS_X1 port map( D => n248, CK => Clk,
                           SN => Rst, Q => n247, QN => n_1086);
   DataP_EX_MEM_s_NPC_L_OUT_reg_27_inst : DFFS_X1 port map( D => n247, CK => 
                           Clk, SN => Rst, Q => n246, QN => n_1087);
   DataP_MEM_WB_s_NPC_L_OUT_reg_27_inst : DFFS_X1 port map( D => n246, CK => 
                           Clk, SN => Rst, Q => n_1088, QN => 
                           DataP_link_addr_W_27_port);
   DataP_IF_IDs_NPC_L_OUT_reg_26_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_26_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1089, QN 
                           => n245);
   DataP_ID_EXs_NPC_L_OUT_reg_26_inst : DFFS_X1 port map( D => n245, CK => Clk,
                           SN => Rst, Q => n244, QN => n_1090);
   DataP_EX_MEM_s_NPC_L_OUT_reg_26_inst : DFFS_X1 port map( D => n244, CK => 
                           Clk, SN => Rst, Q => n243, QN => n_1091);
   DataP_MEM_WB_s_NPC_L_OUT_reg_26_inst : DFFS_X1 port map( D => n243, CK => 
                           Clk, SN => Rst, Q => n_1092, QN => 
                           DataP_link_addr_W_26_port);
   DataP_IF_IDs_NPC_L_OUT_reg_25_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_25_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1093, QN 
                           => n242);
   DataP_ID_EXs_NPC_L_OUT_reg_25_inst : DFFS_X1 port map( D => n242, CK => Clk,
                           SN => Rst, Q => n241, QN => n_1094);
   DataP_EX_MEM_s_NPC_L_OUT_reg_25_inst : DFFS_X1 port map( D => n241, CK => 
                           Clk, SN => Rst, Q => n240, QN => n_1095);
   DataP_MEM_WB_s_NPC_L_OUT_reg_25_inst : DFFS_X1 port map( D => n240, CK => 
                           Clk, SN => Rst, Q => n_1096, QN => 
                           DataP_link_addr_W_25_port);
   DataP_IF_IDs_NPC_L_OUT_reg_24_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_24_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1097, QN 
                           => n239);
   DataP_ID_EXs_NPC_L_OUT_reg_24_inst : DFFS_X1 port map( D => n239, CK => Clk,
                           SN => Rst, Q => n238, QN => n_1098);
   DataP_EX_MEM_s_NPC_L_OUT_reg_24_inst : DFFS_X1 port map( D => n238, CK => 
                           Clk, SN => Rst, Q => n237, QN => n_1099);
   DataP_MEM_WB_s_NPC_L_OUT_reg_24_inst : DFFS_X1 port map( D => n237, CK => 
                           Clk, SN => Rst, Q => n_1100, QN => 
                           DataP_link_addr_W_24_port);
   DataP_IF_IDs_NPC_L_OUT_reg_23_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_23_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1101, QN 
                           => n236);
   DataP_ID_EXs_NPC_L_OUT_reg_23_inst : DFFS_X1 port map( D => n236, CK => Clk,
                           SN => Rst, Q => n235, QN => n_1102);
   DataP_EX_MEM_s_NPC_L_OUT_reg_23_inst : DFFS_X1 port map( D => n235, CK => 
                           Clk, SN => Rst, Q => n234, QN => n_1103);
   DataP_MEM_WB_s_NPC_L_OUT_reg_23_inst : DFFS_X1 port map( D => n234, CK => 
                           Clk, SN => Rst, Q => n_1104, QN => 
                           DataP_link_addr_W_23_port);
   DataP_IF_IDs_NPC_L_OUT_reg_22_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_22_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1105, QN 
                           => n233);
   DataP_ID_EXs_NPC_L_OUT_reg_22_inst : DFFS_X1 port map( D => n233, CK => Clk,
                           SN => Rst, Q => n232, QN => n_1106);
   DataP_EX_MEM_s_NPC_L_OUT_reg_22_inst : DFFS_X1 port map( D => n232, CK => 
                           Clk, SN => Rst, Q => n231, QN => n_1107);
   DataP_MEM_WB_s_NPC_L_OUT_reg_22_inst : DFFS_X1 port map( D => n231, CK => 
                           Clk, SN => Rst, Q => n_1108, QN => 
                           DataP_link_addr_W_22_port);
   DataP_IF_IDs_NPC_L_OUT_reg_21_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_21_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1109, QN 
                           => n230);
   DataP_ID_EXs_NPC_L_OUT_reg_21_inst : DFFS_X1 port map( D => n230, CK => Clk,
                           SN => Rst, Q => n229, QN => n_1110);
   DataP_EX_MEM_s_NPC_L_OUT_reg_21_inst : DFFS_X1 port map( D => n229, CK => 
                           Clk, SN => Rst, Q => n228, QN => n_1111);
   DataP_MEM_WB_s_NPC_L_OUT_reg_21_inst : DFFS_X1 port map( D => n228, CK => 
                           Clk, SN => Rst, Q => n_1112, QN => 
                           DataP_link_addr_W_21_port);
   DataP_IF_IDs_NPC_L_OUT_reg_20_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_20_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1113, QN 
                           => n227);
   DataP_ID_EXs_NPC_L_OUT_reg_20_inst : DFFS_X1 port map( D => n227, CK => Clk,
                           SN => Rst, Q => n226, QN => n_1114);
   DataP_EX_MEM_s_NPC_L_OUT_reg_20_inst : DFFS_X1 port map( D => n226, CK => 
                           Clk, SN => Rst, Q => n225, QN => n_1115);
   DataP_MEM_WB_s_NPC_L_OUT_reg_20_inst : DFFS_X1 port map( D => n225, CK => 
                           Clk, SN => Rst, Q => n_1116, QN => 
                           DataP_link_addr_W_20_port);
   DataP_IF_IDs_NPC_L_OUT_reg_19_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_19_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1117, QN 
                           => n224);
   DataP_ID_EXs_NPC_L_OUT_reg_19_inst : DFFS_X1 port map( D => n224, CK => Clk,
                           SN => Rst, Q => n223, QN => n_1118);
   DataP_EX_MEM_s_NPC_L_OUT_reg_19_inst : DFFS_X1 port map( D => n223, CK => 
                           Clk, SN => Rst, Q => n222, QN => n_1119);
   DataP_MEM_WB_s_NPC_L_OUT_reg_19_inst : DFFS_X1 port map( D => n222, CK => 
                           Clk, SN => Rst, Q => n_1120, QN => 
                           DataP_link_addr_W_19_port);
   DataP_IF_IDs_NPC_L_OUT_reg_18_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_18_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1121, QN 
                           => n221);
   DataP_ID_EXs_NPC_L_OUT_reg_18_inst : DFFS_X1 port map( D => n221, CK => Clk,
                           SN => Rst, Q => n220, QN => n_1122);
   DataP_EX_MEM_s_NPC_L_OUT_reg_18_inst : DFFS_X1 port map( D => n220, CK => 
                           Clk, SN => Rst, Q => n219, QN => n_1123);
   DataP_MEM_WB_s_NPC_L_OUT_reg_18_inst : DFFS_X1 port map( D => n219, CK => 
                           Clk, SN => Rst, Q => n_1124, QN => 
                           DataP_link_addr_W_18_port);
   DataP_IF_IDs_NPC_L_OUT_reg_17_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_17_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1125, QN 
                           => n218);
   DataP_ID_EXs_NPC_L_OUT_reg_17_inst : DFFS_X1 port map( D => n218, CK => Clk,
                           SN => Rst, Q => n217, QN => n_1126);
   DataP_EX_MEM_s_NPC_L_OUT_reg_17_inst : DFFS_X1 port map( D => n217, CK => 
                           Clk, SN => Rst, Q => n216, QN => n_1127);
   DataP_MEM_WB_s_NPC_L_OUT_reg_17_inst : DFFS_X1 port map( D => n216, CK => 
                           Clk, SN => Rst, Q => n_1128, QN => 
                           DataP_link_addr_W_17_port);
   DataP_IF_IDs_NPC_L_OUT_reg_16_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_16_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1129, QN 
                           => n215);
   DataP_ID_EXs_NPC_L_OUT_reg_16_inst : DFFS_X1 port map( D => n215, CK => Clk,
                           SN => Rst, Q => n214, QN => n_1130);
   DataP_EX_MEM_s_NPC_L_OUT_reg_16_inst : DFFS_X1 port map( D => n214, CK => 
                           Clk, SN => Rst, Q => n213, QN => n_1131);
   DataP_MEM_WB_s_NPC_L_OUT_reg_16_inst : DFFS_X1 port map( D => n213, CK => 
                           Clk, SN => Rst, Q => n_1132, QN => 
                           DataP_link_addr_W_16_port);
   DataP_IF_IDs_NPC_L_OUT_reg_15_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_15_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1133, QN 
                           => n212);
   DataP_ID_EXs_NPC_L_OUT_reg_15_inst : DFFS_X1 port map( D => n212, CK => Clk,
                           SN => Rst, Q => n211, QN => n_1134);
   DataP_EX_MEM_s_NPC_L_OUT_reg_15_inst : DFFS_X1 port map( D => n211, CK => 
                           Clk, SN => Rst, Q => n210, QN => n_1135);
   DataP_MEM_WB_s_NPC_L_OUT_reg_15_inst : DFFS_X1 port map( D => n210, CK => 
                           Clk, SN => Rst, Q => n_1136, QN => 
                           DataP_link_addr_W_15_port);
   DataP_IF_IDs_NPC_L_OUT_reg_14_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_14_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1137, QN 
                           => n209);
   DataP_ID_EXs_NPC_L_OUT_reg_14_inst : DFFS_X1 port map( D => n209, CK => Clk,
                           SN => Rst, Q => n208, QN => n_1138);
   DataP_EX_MEM_s_NPC_L_OUT_reg_14_inst : DFFS_X1 port map( D => n208, CK => 
                           Clk, SN => Rst, Q => n207, QN => n_1139);
   DataP_MEM_WB_s_NPC_L_OUT_reg_14_inst : DFFS_X1 port map( D => n207, CK => 
                           Clk, SN => Rst, Q => n_1140, QN => 
                           DataP_link_addr_W_14_port);
   DataP_IF_IDs_NPC_L_OUT_reg_13_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_13_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1141, QN 
                           => n206);
   DataP_ID_EXs_NPC_L_OUT_reg_13_inst : DFFS_X1 port map( D => n206, CK => Clk,
                           SN => Rst, Q => n205, QN => n_1142);
   DataP_EX_MEM_s_NPC_L_OUT_reg_13_inst : DFFS_X1 port map( D => n205, CK => 
                           Clk, SN => Rst, Q => n204, QN => n_1143);
   DataP_MEM_WB_s_NPC_L_OUT_reg_13_inst : DFFS_X1 port map( D => n204, CK => 
                           Clk, SN => Rst, Q => n_1144, QN => 
                           DataP_link_addr_W_13_port);
   DataP_IF_IDs_NPC_L_OUT_reg_12_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_12_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1145, QN 
                           => n203);
   DataP_ID_EXs_NPC_L_OUT_reg_12_inst : DFFS_X1 port map( D => n203, CK => Clk,
                           SN => Rst, Q => n202, QN => n_1146);
   DataP_EX_MEM_s_NPC_L_OUT_reg_12_inst : DFFS_X1 port map( D => n202, CK => 
                           Clk, SN => Rst, Q => n201, QN => n_1147);
   DataP_MEM_WB_s_NPC_L_OUT_reg_12_inst : DFFS_X1 port map( D => n201, CK => 
                           Clk, SN => Rst, Q => n_1148, QN => 
                           DataP_link_addr_W_12_port);
   DataP_IF_IDs_NPC_L_OUT_reg_11_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_11_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1149, QN 
                           => n200);
   DataP_ID_EXs_NPC_L_OUT_reg_11_inst : DFFS_X1 port map( D => n200, CK => Clk,
                           SN => Rst, Q => n199, QN => n_1150);
   DataP_EX_MEM_s_NPC_L_OUT_reg_11_inst : DFFS_X1 port map( D => n199, CK => 
                           Clk, SN => Rst, Q => n198, QN => n_1151);
   DataP_MEM_WB_s_NPC_L_OUT_reg_11_inst : DFFS_X1 port map( D => n198, CK => 
                           Clk, SN => Rst, Q => n_1152, QN => 
                           DataP_link_addr_W_11_port);
   DataP_IF_IDs_NPC_L_OUT_reg_10_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_10_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1153, QN 
                           => n197);
   DataP_ID_EXs_NPC_L_OUT_reg_10_inst : DFFS_X1 port map( D => n197, CK => Clk,
                           SN => Rst, Q => n196, QN => n_1154);
   DataP_EX_MEM_s_NPC_L_OUT_reg_10_inst : DFFS_X1 port map( D => n196, CK => 
                           Clk, SN => Rst, Q => n195, QN => n_1155);
   DataP_MEM_WB_s_NPC_L_OUT_reg_10_inst : DFFS_X1 port map( D => n195, CK => 
                           Clk, SN => Rst, Q => n_1156, QN => 
                           DataP_link_addr_W_10_port);
   DataP_IF_IDs_NPC_L_OUT_reg_9_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_9_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1157, QN 
                           => n194);
   DataP_ID_EXs_NPC_L_OUT_reg_9_inst : DFFS_X1 port map( D => n194, CK => Clk, 
                           SN => Rst, Q => n193, QN => n_1158);
   DataP_EX_MEM_s_NPC_L_OUT_reg_9_inst : DFFS_X1 port map( D => n193, CK => Clk
                           , SN => Rst, Q => n192, QN => n_1159);
   DataP_MEM_WB_s_NPC_L_OUT_reg_9_inst : DFFS_X1 port map( D => n192, CK => Clk
                           , SN => Rst, Q => n_1160, QN => 
                           DataP_link_addr_W_9_port);
   DataP_IF_IDs_NPC_L_OUT_reg_8_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_8_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1161, QN 
                           => n191);
   DataP_ID_EXs_NPC_L_OUT_reg_8_inst : DFFS_X1 port map( D => n191, CK => Clk, 
                           SN => Rst, Q => n190, QN => n_1162);
   DataP_EX_MEM_s_NPC_L_OUT_reg_8_inst : DFFS_X1 port map( D => n190, CK => Clk
                           , SN => Rst, Q => n189, QN => n_1163);
   DataP_MEM_WB_s_NPC_L_OUT_reg_8_inst : DFFS_X1 port map( D => n189, CK => Clk
                           , SN => Rst, Q => n_1164, QN => 
                           DataP_link_addr_W_8_port);
   DataP_IF_IDs_NPC_L_OUT_reg_7_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_7_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1165, QN 
                           => n188);
   DataP_ID_EXs_NPC_L_OUT_reg_7_inst : DFFS_X1 port map( D => n188, CK => Clk, 
                           SN => Rst, Q => n187, QN => n_1166);
   DataP_EX_MEM_s_NPC_L_OUT_reg_7_inst : DFFS_X1 port map( D => n187, CK => Clk
                           , SN => Rst, Q => n186, QN => n_1167);
   DataP_MEM_WB_s_NPC_L_OUT_reg_7_inst : DFFS_X1 port map( D => n186, CK => Clk
                           , SN => Rst, Q => n_1168, QN => 
                           DataP_link_addr_W_7_port);
   DataP_IF_IDs_NPC_L_OUT_reg_6_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_6_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1169, QN 
                           => n185);
   DataP_ID_EXs_NPC_L_OUT_reg_6_inst : DFFS_X1 port map( D => n185, CK => Clk, 
                           SN => Rst, Q => n184, QN => n_1170);
   DataP_EX_MEM_s_NPC_L_OUT_reg_6_inst : DFFS_X1 port map( D => n184, CK => Clk
                           , SN => Rst, Q => n183, QN => n_1171);
   DataP_MEM_WB_s_NPC_L_OUT_reg_6_inst : DFFS_X1 port map( D => n183, CK => Clk
                           , SN => Rst, Q => n_1172, QN => 
                           DataP_link_addr_W_6_port);
   DataP_IF_IDs_NPC_L_OUT_reg_5_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_5_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1173, QN 
                           => n182);
   DataP_ID_EXs_NPC_L_OUT_reg_5_inst : DFFS_X1 port map( D => n182, CK => Clk, 
                           SN => Rst, Q => n181, QN => n_1174);
   DataP_EX_MEM_s_NPC_L_OUT_reg_5_inst : DFFS_X1 port map( D => n181, CK => Clk
                           , SN => Rst, Q => n180, QN => n_1175);
   DataP_MEM_WB_s_NPC_L_OUT_reg_5_inst : DFFS_X1 port map( D => n180, CK => Clk
                           , SN => Rst, Q => n_1176, QN => 
                           DataP_link_addr_W_5_port);
   DataP_IF_IDs_NPC_L_OUT_reg_4_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_4_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1177, QN 
                           => n179);
   DataP_ID_EXs_NPC_L_OUT_reg_4_inst : DFFS_X1 port map( D => n179, CK => Clk, 
                           SN => Rst, Q => n178, QN => n_1178);
   DataP_EX_MEM_s_NPC_L_OUT_reg_4_inst : DFFS_X1 port map( D => n178, CK => Clk
                           , SN => Rst, Q => n177, QN => n_1179);
   DataP_MEM_WB_s_NPC_L_OUT_reg_4_inst : DFFS_X1 port map( D => n177, CK => Clk
                           , SN => Rst, Q => n_1180, QN => 
                           DataP_link_addr_W_4_port);
   DataP_IF_IDs_NPC_L_OUT_reg_3_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_3_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1181, QN 
                           => n176);
   DataP_ID_EXs_NPC_L_OUT_reg_3_inst : DFFS_X1 port map( D => n176, CK => Clk, 
                           SN => Rst, Q => n175, QN => n_1182);
   DataP_EX_MEM_s_NPC_L_OUT_reg_3_inst : DFFS_X1 port map( D => n175, CK => Clk
                           , SN => Rst, Q => n174, QN => n_1183);
   DataP_MEM_WB_s_NPC_L_OUT_reg_3_inst : DFFS_X1 port map( D => n174, CK => Clk
                           , SN => Rst, Q => n_1184, QN => 
                           DataP_link_addr_W_3_port);
   DataP_IF_IDs_NPC_L_OUT_reg_2_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_2_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1185, QN 
                           => n173);
   DataP_ID_EXs_NPC_L_OUT_reg_2_inst : DFFS_X1 port map( D => n173, CK => Clk, 
                           SN => Rst, Q => n172, QN => n_1186);
   DataP_EX_MEM_s_NPC_L_OUT_reg_2_inst : DFFS_X1 port map( D => n172, CK => Clk
                           , SN => Rst, Q => n171, QN => n_1187);
   DataP_MEM_WB_s_NPC_L_OUT_reg_2_inst : DFFS_X1 port map( D => n171, CK => Clk
                           , SN => Rst, Q => n_1188, QN => 
                           DataP_link_addr_W_2_port);
   DataP_IF_IDs_NPC_L_OUT_reg_1_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_1_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1189, QN 
                           => n170);
   DataP_ID_EXs_NPC_L_OUT_reg_1_inst : DFFS_X1 port map( D => n170, CK => Clk, 
                           SN => Rst, Q => n169, QN => n_1190);
   DataP_EX_MEM_s_NPC_L_OUT_reg_1_inst : DFFS_X1 port map( D => n169, CK => Clk
                           , SN => Rst, Q => n168, QN => n_1191);
   DataP_MEM_WB_s_NPC_L_OUT_reg_1_inst : DFFS_X1 port map( D => n168, CK => Clk
                           , SN => Rst, Q => n_1192, QN => 
                           DataP_link_addr_W_1_port);
   DataP_IF_IDs_NPC_L_OUT_reg_0_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_F_0_port, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1193, QN 
                           => n167);
   DataP_ID_EXs_NPC_L_OUT_reg_0_inst : DFFS_X1 port map( D => n167, CK => Clk, 
                           SN => Rst, Q => n166, QN => n_1194);
   DataP_EX_MEM_s_NPC_L_OUT_reg_0_inst : DFFS_X1 port map( D => n166, CK => Clk
                           , SN => Rst, Q => n165, QN => n_1195);
   DataP_MEM_WB_s_NPC_L_OUT_reg_0_inst : DFFS_X1 port map( D => n165, CK => Clk
                           , SN => Rst, Q => n_1196, QN => 
                           DataP_link_addr_W_0_port);
   DataP_IF_IDs_IR_OUT_reg_0_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(0), CK
                           => Clk, RN => n164, Q => IR_CU_0_port, QN => n476);
   DataP_ID_EXs_IR_OUT_reg_0_inst : DFFS_X1 port map( D => n476, CK => Clk, SN 
                           => Rst, Q => n_1197, QN => DataP_ir_E_0_port);
   DataP_IF_IDs_IR_OUT_reg_1_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(1), CK
                           => Clk, RN => n164, Q => IR_CU_1_port, QN => n477);
   DataP_ID_EXs_IR_OUT_reg_1_inst : DFFS_X1 port map( D => n477, CK => Clk, SN 
                           => Rst, Q => n_1198, QN => DataP_ir_E_1_port);
   DataP_IF_IDs_IR_OUT_reg_2_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(2), CK
                           => Clk, RN => n164, Q => n2128, QN => n478);
   DataP_ID_EXs_IR_OUT_reg_2_inst : DFFS_X1 port map( D => n478, CK => Clk, SN 
                           => Rst, Q => n_1199, QN => DataP_ir_E_2_port);
   DataP_IF_IDs_IR_OUT_reg_3_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(3), CK
                           => Clk, RN => n164, Q => n2135, QN => n479);
   DataP_ID_EXs_IR_OUT_reg_3_inst : DFFS_X1 port map( D => n479, CK => Clk, SN 
                           => Rst, Q => n_1200, QN => DataP_ir_E_3_port);
   DataP_IF_IDs_IR_OUT_reg_4_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(4), CK
                           => Clk, RN => n164, Q => IR_CU_4_port, QN => n480);
   DataP_ID_EXs_IR_OUT_reg_4_inst : DFFS_X1 port map( D => n480, CK => Clk, SN 
                           => Rst, Q => n_1201, QN => DataP_ir_E_4_port);
   DataP_IF_IDs_IR_OUT_reg_5_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(5), CK
                           => Clk, RN => n164, Q => IR_CU_5_port, QN => n482);
   DataP_ID_EXs_IR_OUT_reg_5_inst : DFFS_X1 port map( D => n482, CK => Clk, SN 
                           => Rst, Q => n_1202, QN => DataP_ir_E_5_port);
   DataP_IF_IDs_IR_OUT_reg_6_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(6), CK
                           => Clk, RN => n164, Q => IR_CU_6_port, QN => n163);
   DataP_ID_EXs_IR_OUT_reg_6_inst : DFFS_X1 port map( D => n163, CK => Clk, SN 
                           => Rst, Q => n_1203, QN => DataP_ir_E_6_port);
   DataP_IF_IDs_IR_OUT_reg_7_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(7), CK
                           => Clk, RN => n164, Q => IR_CU_7_port, QN => n162);
   DataP_ID_EXs_IR_OUT_reg_7_inst : DFFS_X1 port map( D => n162, CK => Clk, SN 
                           => Rst, Q => n_1204, QN => DataP_ir_E_7_port);
   DataP_IF_IDs_IR_OUT_reg_8_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(8), CK
                           => Clk, RN => n164, Q => IR_CU_8_port, QN => n161);
   DataP_ID_EXs_IR_OUT_reg_8_inst : DFFS_X1 port map( D => n161, CK => Clk, SN 
                           => Rst, Q => n_1205, QN => DataP_ir_E_8_port);
   DataP_IF_IDs_IR_OUT_reg_9_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(9), CK
                           => Clk, RN => n164, Q => IR_CU_9_port, QN => n160);
   DataP_ID_EXs_IR_OUT_reg_9_inst : DFFS_X1 port map( D => n160, CK => Clk, SN 
                           => Rst, Q => n_1206, QN => DataP_ir_E_9_port);
   DataP_IF_IDs_IR_OUT_reg_10_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(10), 
                           CK => Clk, RN => n164, Q => n_1207, QN => n484);
   DataP_ID_EXs_IR_OUT_reg_10_inst : DFFS_X1 port map( D => n484, CK => Clk, SN
                           => Rst, Q => n_1208, QN => DataP_ir_E_10_port);
   DataP_IF_IDs_IR_OUT_reg_11_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(11), 
                           CK => Clk, RN => n164, Q => DataP_IR1_11_port, QN =>
                           n159);
   DataP_ID_EXs_IR_OUT_reg_11_inst : DFFS_X1 port map( D => n159, CK => Clk, SN
                           => Rst, Q => n_1209, QN => DataP_ir_E_11_port);
   DataP_IF_IDs_IR_OUT_reg_12_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(12), 
                           CK => Clk, RN => n164, Q => DataP_IR1_12_port, QN =>
                           n158);
   DataP_ID_EXs_IR_OUT_reg_12_inst : DFFS_X1 port map( D => n158, CK => Clk, SN
                           => Rst, Q => n_1210, QN => DataP_ir_E_12_port);
   DataP_IF_IDs_IR_OUT_reg_13_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(13), 
                           CK => Clk, RN => n164, Q => DataP_IR1_13_port, QN =>
                           n157);
   DataP_ID_EXs_IR_OUT_reg_13_inst : DFFS_X1 port map( D => n157, CK => Clk, SN
                           => Rst, Q => n_1211, QN => DataP_ir_E_13_port);
   DataP_IF_IDs_IR_OUT_reg_14_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(14), 
                           CK => Clk, RN => n164, Q => DataP_IR1_14_port, QN =>
                           n156);
   DataP_ID_EXs_IR_OUT_reg_14_inst : DFFS_X1 port map( D => n156, CK => Clk, SN
                           => Rst, Q => n_1212, QN => DataP_ir_E_14_port);
   DataP_IF_IDs_IR_OUT_reg_15_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(15), 
                           CK => Clk, RN => n164, Q => DataP_IR1_15_port, QN =>
                           n155);
   DataP_ID_EXs_IR_OUT_reg_15_inst : DFFS_X1 port map( D => n155, CK => Clk, SN
                           => Rst, Q => n_1213, QN => DataP_ir_E_15_port);
   DataP_IF_IDs_IR_OUT_reg_16_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(16), 
                           CK => Clk, RN => n164, Q => n_1214, QN => n485);
   DataP_IF_IDs_IR_OUT_reg_17_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(17), 
                           CK => Clk, RN => n164, Q => n_1215, QN => n486);
   DataP_IF_IDs_IR_OUT_reg_18_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(18), 
                           CK => Clk, RN => n164, Q => n_1216, QN => n487);
   DataP_IF_IDs_IR_OUT_reg_19_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(19), 
                           CK => Clk, RN => n164, Q => n_1217, QN => n488);
   DataP_IF_IDs_IR_OUT_reg_20_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(20), 
                           CK => Clk, RN => n164, Q => n_1218, QN => n489);
   DataP_IF_IDs_IR_OUT_reg_21_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(21), 
                           CK => Clk, RN => n164, Q => DataP_IR1_21_port, QN =>
                           n_1219);
   DataP_IF_IDs_IR_OUT_reg_22_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(22), 
                           CK => Clk, RN => n164, Q => DataP_IR1_22_port, QN =>
                           n153);
   DataP_IF_IDs_IR_OUT_reg_23_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(23), 
                           CK => Clk, RN => n164, Q => DataP_IR1_23_port, QN =>
                           n152);
   DataP_ID_EXs_RS1_OUT_reg_2_inst : DFFS_X1 port map( D => n152, CK => Clk, SN
                           => Rst, Q => n2156, QN => DataP_Rs1_2_port);
   DataP_IF_IDs_IR_OUT_reg_24_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(24), 
                           CK => Clk, RN => n164, Q => DataP_IR1_24_port, QN =>
                           n_1220);
   DataP_IF_IDs_IR_OUT_reg_25_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(25), 
                           CK => Clk, RN => n164, Q => DataP_IR1_25_port, QN =>
                           n_1221);
   DataP_ID_EXs_RS1_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_IR1_25_port, 
                           CK => Clk, RN => Rst, Q => n_1222, QN => n524);
   DataP_IF_IDs_IR_OUT_reg_26_inst : DFFS_X1 port map( D => IRAM_DATA_OUT(26), 
                           CK => Clk, SN => n164, Q => IR_CU_26, QN => n497);
   DataP_MEM_WB_s_OPCODE_OUT_reg_0_inst : DFFS_X1 port map( D => n150, CK => 
                           Clk, SN => Rst, Q => n2162, QN => 
                           DataP_opcode_W_0_port);
   DataP_IF_IDs_IR_OUT_reg_27_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(27), 
                           CK => Clk, RN => n164, Q => IR_CU_27, QN => n504);
   DataP_EX_MEM_s_OPCODE_OUT_reg_1_inst : DFFS_X1 port map( D => n520, CK => 
                           Clk, SN => Rst, Q => n2576, QN => 
                           DataP_opcode_M_1_port);
   DataP_ID_EXs_OPCODE_OUT_reg_2_inst : DFFS_X1 port map( D => n510, CK => Clk,
                           SN => Rst, Q => n521, QN => n2574);
   DataP_IF_IDs_IR_OUT_reg_29_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(29), 
                           CK => Clk, RN => n164, Q => n2141, QN => n514);
   DataP_ID_EXs_OPCODE_OUT_reg_3_inst : DFFS_X1 port map( D => n514, CK => Clk,
                           SN => Rst, Q => n149, QN => DataP_opcode_E_3_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_3_inst : DFFS_X1 port map( D => n149, CK => 
                           Clk, SN => Rst, Q => n148, QN => 
                           DataP_opcode_M_3_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_3_inst : DFFS_X1 port map( D => n148, CK => 
                           Clk, SN => Rst, Q => n2159, QN => 
                           DataP_opcode_W_3_port);
   DataP_ID_EXs_OPCODE_OUT_reg_4_inst : DFFS_X1 port map( D => n515, CK => Clk,
                           SN => Rst, Q => n147, QN => DataP_opcode_E_4_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_4_inst : DFFS_X1 port map( D => n146, CK => 
                           Clk, SN => Rst, Q => n2151, QN => 
                           DataP_opcode_W_4_port);
   DataP_IF_IDs_IR_OUT_reg_31_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(31), 
                           CK => Clk, RN => n164, Q => IR_CU_31, QN => n516);
   DataP_ID_EXs_OPCODE_OUT_reg_5_inst : DFFS_X1 port map( D => n516, CK => Clk,
                           SN => Rst, Q => n145, QN => n_1223);
   DataP_EX_MEM_s_OPCODE_OUT_reg_5_inst : DFFS_X1 port map( D => n145, CK => 
                           Clk, SN => Rst, Q => n2161, QN => 
                           DataP_opcode_M_5_port);
   DataP_FORWARDING_BR_SEL_reg_1_inst : DLH_X1 port map( G => 
                           DataP_FORWARDING_BR_N12, D => n3710, Q => 
                           DataP_FWD_MUX_BR_S_1_port);
   CU_I_cw1_reg_8_inst : SDFFR_X1 port map( D => n144, SI => n606, SE => n504, 
                           CK => Clk, RN => Rst, Q => BR_EN_i, QN => n_1224);
   CU_I_aluOpcode1_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_3_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_3_port, QN 
                           => n2146);
   CU_I_cw1_reg_10_inst : DFFR_X1 port map( D => CU_I_cw_10_port, CK => Clk, RN
                           => Rst, Q => n2155, QN => n432);
   CU_I_cw2_reg_7_inst : DFFS_X1 port map( D => n143, CK => Clk, SN => Rst, Q 
                           => n_1225, QN => DRAM_RW);
   DataP_ID_EXs_RS2_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_add_S2_2_port
                           , CK => Clk, RN => Rst, Q => DataP_Rs2_2_port, QN =>
                           n_1226);
   DataP_EX_MEM_s_RD_OUT_reg_4_inst : DFFS_X1 port map( D => n142, CK => Clk, 
                           SN => Rst, Q => n2569, QN => DataP_dest_M_4_port);
   DataP_MEM_WB_s_RD_OUT_reg_4_inst : DFFR_X1 port map( D => 
                           DataP_dest_M_4_port, CK => Clk, RN => Rst, Q => 
                           DataP_add_D_4_port, QN => n540);
   DataP_EX_MEM_s_RD_OUT_reg_3_inst : DFFS_X1 port map( D => n141, CK => Clk, 
                           SN => Rst, Q => n2570, QN => DataP_dest_M_3_port);
   DataP_EX_MEM_s_RD_OUT_reg_2_inst : DFFS_X1 port map( D => n140, CK => Clk, 
                           SN => Rst, Q => n530, QN => DataP_dest_M_2_port);
   DataP_EX_MEM_s_RD_OUT_reg_1_inst : DFFS_X1 port map( D => n139, CK => Clk, 
                           SN => Rst, Q => n529, QN => DataP_dest_M_1_port);
   DataP_MEM_WB_s_RD_OUT_reg_0_inst : DFFR_X1 port map( D => 
                           DataP_dest_M_0_port, CK => Clk, RN => Rst, Q => 
                           DataP_add_D_0_port, QN => n536);
   DataP_FORWARDING_BR_SEL_reg_0_inst : DLH_X1 port map( G => 
                           DataP_FORWARDING_BR_N12, D => n2469, Q => 
                           DataP_FWD_MUX_BR_S_0_port);
   CU_I_aluOpcode1_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_0_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_0_port, QN 
                           => n2150);
   CU_I_aluOpcode1_reg_4_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_4_port,
                           CK => Clk, RN => Rst, Q => n2134, QN => n443);
   CU_I_aluOpcode1_reg_2_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_2_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_2_port, QN 
                           => n2144);
   CU_I_aluOpcode1_reg_1_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_1_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_1_port, QN 
                           => n2132);
   CU_I_cw1_reg_5_inst : DFFS_X1 port map( D => n1357, CK => Clk, SN => Rst, Q 
                           => n137, QN => n_1227);
   CU_I_cw2_reg_5_inst : DFFS_X1 port map( D => n137, CK => Clk, SN => Rst, Q 
                           => n_1228, QN => DRAM_SEL(2));
   CU_I_cw2_reg_0_inst : DFFS_X1 port map( D => n136, CK => Clk, SN => Rst, Q 
                           => n135, QN => n_1229);
   CU_I_cw3_reg_0_inst : DFFS_X1 port map( D => n135, CK => Clk, SN => Rst, Q 
                           => n_1230, QN => RF_WE_i);
   CU_I_cw1_reg_2_inst : DFFS_X1 port map( D => n1371, CK => Clk, SN => Rst, Q 
                           => n134, QN => n_1231);
   CU_I_cw2_reg_2_inst : DFFS_X1 port map( D => n134, CK => Clk, SN => Rst, Q 
                           => n133, QN => n_1232);
   CU_I_cw3_reg_2_inst : DFFS_X1 port map( D => n133, CK => Clk, SN => Rst, Q 
                           => n_1233, QN => WB_MUX_SEL_i_1_port);
   CU_I_cw2_reg_4_inst : DFFS_X1 port map( D => n132, CK => Clk, SN => Rst, Q 
                           => n_1234, QN => DRAM_SEL(1));
   CU_I_cw2_reg_3_inst : DFFS_X1 port map( D => n131, CK => Clk, SN => Rst, Q 
                           => n_1235, QN => DRAM_SEL(0));
   CU_I_cw2_reg_6_inst : DFFS_X1 port map( D => n130, CK => Clk, SN => Rst, Q 
                           => n_1236, QN => DRAM_ENABLE);
   CU_I_cw1_reg_9_inst : DFFR_X1 port map( D => CU_I_cw_9_port, CK => Clk, RN 
                           => Rst, Q => n2189, QN => n399);
   CU_I_cw2_reg_1_inst : DFFS_X1 port map( D => n129, CK => Clk, SN => Rst, Q 
                           => n_1237, QN => CU_I_cw2_1_port);
   CU_I_cw3_reg_1_inst : DFFR_X1 port map( D => CU_I_cw2_1_port, CK => Clk, RN 
                           => Rst, Q => n_1238, QN => n294);
   DataP_ID_EXs_IMM_OUT_reg_31_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_31_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_31_port, QN => n_1239);
   DataP_ID_EXs_IMM_OUT_reg_24_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_24_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_24_port, QN => n_1240);
   DataP_ID_EXs_IMM_OUT_reg_23_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_23_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_23_port, QN => n_1241);
   DataP_ID_EXs_IMM_OUT_reg_22_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_22_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_22_port, QN => n_1242);
   DataP_ID_EXs_IMM_OUT_reg_21_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_21_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_21_port, QN => n_1243);
   DataP_ID_EXs_IMM_OUT_reg_20_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_20_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_20_port, QN => n_1244);
   DataP_ID_EXs_IMM_OUT_reg_19_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_19_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_19_port, QN => n_1245);
   DataP_ID_EXs_IMM_OUT_reg_18_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_18_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_18_port, QN => n_1246);
   DataP_ID_EXs_IMM_OUT_reg_17_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_17_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_17_port, QN => n_1247);
   DataP_ID_EXs_IMM_OUT_reg_16_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_16_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_16_port, QN => n_1248);
   DataP_IF_IDs_NPC_OUT_reg_0_inst : DFFRS_X1 port map( D => DataP_npc_0_port, 
                           CK => Clk, RN => n126, SN => n127, Q => n_1249, QN 
                           => n128);
   DataP_ID_EXs_NPC_OUT_reg_0_inst : DFFS_X1 port map( D => n128, CK => Clk, SN
                           => Rst, Q => n125, QN => n_1250);
   DataP_EX_MEM_s_NPC_OUT_reg_0_inst : DFFS_X1 port map( D => n125, CK => Clk, 
                           SN => Rst, Q => n_1251, QN => DataP_npc_M_0_port);
   DataP_IF_IDs_NPC_OUT_reg_1_inst : DFFRS_X1 port map( D => DataP_npc_1_port, 
                           CK => Clk, RN => n122, SN => n123, Q => n_1252, QN 
                           => n124);
   DataP_ID_EXs_NPC_OUT_reg_1_inst : DFFS_X1 port map( D => n124, CK => Clk, SN
                           => Rst, Q => n121, QN => n_1253);
   DataP_EX_MEM_s_NPC_OUT_reg_1_inst : DFFS_X1 port map( D => n121, CK => Clk, 
                           SN => Rst, Q => n_1254, QN => DataP_npc_M_1_port);
   DataP_EX_MEM_s_ALU_OUT_reg_1_inst : DFFS_X1 port map( D => n358, CK => Clk, 
                           SN => Rst, Q => n2233, QN => DRAM_ADDRESS_1_port);
   DataP_MEM_WB_s_ALU_OUT_reg_1_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_1_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_1_port, QN => n2273);
   DataP_PC_reg_O_reg_1_inst : DFF_X1 port map( D => DataP_PC_reg_N3, CK => Clk
                           , Q => DataP_pc_out_1, QN => n_1255);
   DataP_IF_IDs_NPC_OUT_reg_2_inst : DFFRS_X1 port map( D => DataP_npc_2_port, 
                           CK => Clk, RN => n118, SN => n119, Q => n_1256, QN 
                           => n120);
   DataP_ID_EXs_NPC_OUT_reg_2_inst : DFFS_X1 port map( D => n120, CK => Clk, SN
                           => Rst, Q => n117, QN => n_1257);
   DataP_EX_MEM_s_NPC_OUT_reg_2_inst : DFFS_X1 port map( D => n117, CK => Clk, 
                           SN => Rst, Q => n_1258, QN => DataP_npc_M_2_port);
   DataP_EX_MEM_s_ALU_OUT_reg_2_inst : DFFS_X1 port map( D => n357, CK => Clk, 
                           SN => Rst, Q => n2232, QN => DRAM_ADDRESS_2_port);
   DataP_MEM_WB_s_ALU_OUT_reg_2_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_2_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_2_port, QN => n2276);
   DataP_PC_reg_O_reg_2_inst : DFF_X1 port map( D => DataP_PC_reg_N4, CK => Clk
                           , Q => IRAM_ADDRESS_0_port, QN => n_1259);
   DataP_IF_IDs_NPC_OUT_reg_3_inst : DFFRS_X1 port map( D => DataP_npc_3_port, 
                           CK => Clk, RN => n114, SN => n115, Q => n_1260, QN 
                           => n116);
   DataP_ID_EXs_NPC_OUT_reg_3_inst : DFFS_X1 port map( D => n116, CK => Clk, SN
                           => Rst, Q => n113, QN => n_1261);
   DataP_EX_MEM_s_NPC_OUT_reg_3_inst : DFFS_X1 port map( D => n113, CK => Clk, 
                           SN => Rst, Q => n_1262, QN => DataP_npc_M_3_port);
   DataP_EX_MEM_s_ALU_OUT_reg_3_inst : DFFS_X1 port map( D => n356, CK => Clk, 
                           SN => Rst, Q => n2231, QN => DRAM_ADDRESS_3_port);
   DataP_MEM_WB_s_ALU_OUT_reg_3_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_3_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_3_port, QN => n2277);
   DataP_PC_reg_O_reg_3_inst : DFF_X1 port map( D => DataP_PC_reg_N5, CK => Clk
                           , Q => IRAM_ADDRESS_1_port, QN => n_1263);
   DataP_IF_IDs_NPC_OUT_reg_4_inst : DFFRS_X1 port map( D => DataP_npc_4_port, 
                           CK => Clk, RN => n110, SN => n111, Q => n_1264, QN 
                           => n112);
   DataP_ID_EXs_NPC_OUT_reg_4_inst : DFFS_X1 port map( D => n112, CK => Clk, SN
                           => Rst, Q => n109, QN => n_1265);
   DataP_EX_MEM_s_NPC_OUT_reg_4_inst : DFFS_X1 port map( D => n109, CK => Clk, 
                           SN => Rst, Q => n_1266, QN => DataP_npc_M_4_port);
   DataP_EX_MEM_s_ALU_OUT_reg_4_inst : DFFS_X1 port map( D => n355, CK => Clk, 
                           SN => Rst, Q => n2229, QN => DRAM_ADDRESS_4_port);
   DataP_MEM_WB_s_ALU_OUT_reg_4_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_4_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_4_port, QN => n2274);
   DataP_PC_reg_O_reg_4_inst : DFF_X1 port map( D => DataP_PC_reg_N6, CK => Clk
                           , Q => IRAM_ADDRESS_2_port, QN => n_1267);
   DataP_IF_IDs_NPC_OUT_reg_5_inst : DFFRS_X1 port map( D => DataP_npc_5_port, 
                           CK => Clk, RN => n106, SN => n107, Q => n_1268, QN 
                           => n108);
   DataP_ID_EXs_NPC_OUT_reg_5_inst : DFFS_X1 port map( D => n108, CK => Clk, SN
                           => Rst, Q => n105, QN => n_1269);
   DataP_EX_MEM_s_NPC_OUT_reg_5_inst : DFFS_X1 port map( D => n105, CK => Clk, 
                           SN => Rst, Q => n_1270, QN => DataP_npc_M_5_port);
   DataP_EX_MEM_s_ALU_OUT_reg_5_inst : DFFS_X1 port map( D => n354, CK => Clk, 
                           SN => Rst, Q => n2227, QN => DRAM_ADDRESS_5_port);
   DataP_MEM_WB_s_ALU_OUT_reg_5_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_5_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_5_port, QN => n2270);
   DataP_PC_reg_O_reg_5_inst : DFF_X1 port map( D => DataP_PC_reg_N7, CK => Clk
                           , Q => IRAM_ADDRESS_3_port, QN => n_1271);
   DataP_IF_IDs_NPC_OUT_reg_6_inst : DFFRS_X1 port map( D => DataP_npc_6_port, 
                           CK => Clk, RN => n102, SN => n103, Q => n_1272, QN 
                           => n104);
   DataP_ID_EXs_NPC_OUT_reg_6_inst : DFFS_X1 port map( D => n104, CK => Clk, SN
                           => Rst, Q => n101, QN => n_1273);
   DataP_EX_MEM_s_NPC_OUT_reg_6_inst : DFFS_X1 port map( D => n101, CK => Clk, 
                           SN => Rst, Q => n_1274, QN => DataP_npc_M_6_port);
   DataP_EX_MEM_s_ALU_OUT_reg_6_inst : DFFS_X1 port map( D => n353, CK => Clk, 
                           SN => Rst, Q => n2182, QN => DRAM_ADDRESS_6_port);
   DataP_MEM_WB_s_ALU_OUT_reg_6_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_6_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_6_port, QN => n2268);
   DataP_PC_reg_O_reg_6_inst : DFF_X1 port map( D => DataP_PC_reg_N8, CK => Clk
                           , Q => IRAM_ADDRESS_4_port, QN => n_1275);
   DataP_IF_IDs_NPC_OUT_reg_7_inst : DFFRS_X1 port map( D => DataP_npc_7_port, 
                           CK => Clk, RN => n98, SN => n99, Q => n_1276, QN => 
                           n100);
   DataP_ID_EXs_NPC_OUT_reg_7_inst : DFFS_X1 port map( D => n100, CK => Clk, SN
                           => Rst, Q => n97, QN => n_1277);
   DataP_EX_MEM_s_NPC_OUT_reg_7_inst : DFFS_X1 port map( D => n97, CK => Clk, 
                           SN => Rst, Q => n_1278, QN => DataP_npc_M_7_port);
   DataP_IF_IDs_NPC_OUT_reg_8_inst : DFFRS_X1 port map( D => DataP_npc_8_port, 
                           CK => Clk, RN => n94, SN => n95, Q => n_1279, QN => 
                           n96);
   DataP_ID_EXs_NPC_OUT_reg_8_inst : DFFS_X1 port map( D => n96, CK => Clk, SN 
                           => Rst, Q => n93, QN => n_1280);
   DataP_EX_MEM_s_NPC_OUT_reg_8_inst : DFFS_X1 port map( D => n93, CK => Clk, 
                           SN => Rst, Q => n_1281, QN => DataP_npc_M_8_port);
   DataP_EX_MEM_s_ALU_OUT_reg_8_inst : DFFS_X1 port map( D => n345, CK => Clk, 
                           SN => Rst, Q => n_1282, QN => DRAM_ADDRESS_8_port);
   DataP_MEM_WB_s_ALU_OUT_reg_8_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_8_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_8_port, QN => n2271);
   DataP_PC_reg_O_reg_8_inst : DFF_X1 port map( D => DataP_PC_reg_N10, CK => 
                           Clk, Q => IRAM_ADDRESS_6_port, QN => n_1283);
   DataP_IF_IDs_NPC_OUT_reg_9_inst : DFFRS_X1 port map( D => DataP_npc_9_port, 
                           CK => Clk, RN => n90, SN => n91, Q => n_1284, QN => 
                           n92);
   DataP_ID_EXs_NPC_OUT_reg_9_inst : DFFS_X1 port map( D => n92, CK => Clk, SN 
                           => Rst, Q => n89, QN => n_1285);
   DataP_EX_MEM_s_NPC_OUT_reg_9_inst : DFFS_X1 port map( D => n89, CK => Clk, 
                           SN => Rst, Q => n_1286, QN => DataP_npc_M_9_port);
   DataP_EX_MEM_s_ALU_OUT_reg_9_inst : DFFS_X1 port map( D => n341, CK => Clk, 
                           SN => Rst, Q => n2228, QN => DRAM_ADDRESS_9_port);
   DataP_MEM_WB_s_ALU_OUT_reg_9_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_9_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_9_port, QN => n2269);
   DataP_PC_reg_O_reg_9_inst : DFF_X1 port map( D => DataP_PC_reg_N11, CK => 
                           Clk, Q => IRAM_ADDRESS_7_port, QN => n_1287);
   DataP_IF_IDs_NPC_OUT_reg_10_inst : DFFRS_X1 port map( D => DataP_npc_10_port
                           , CK => Clk, RN => n86, SN => n87, Q => n_1288, QN 
                           => n88);
   DataP_ID_EXs_NPC_OUT_reg_10_inst : DFFS_X1 port map( D => n88, CK => Clk, SN
                           => Rst, Q => n85, QN => n_1289);
   DataP_EX_MEM_s_NPC_OUT_reg_10_inst : DFFS_X1 port map( D => n85, CK => Clk, 
                           SN => Rst, Q => n_1290, QN => DataP_npc_M_10_port);
   DataP_EX_MEM_s_ALU_OUT_reg_10_inst : DFFS_X1 port map( D => n340, CK => Clk,
                           SN => Rst, Q => n_1291, QN => DRAM_ADDRESS_10_port);
   DataP_MEM_WB_s_ALU_OUT_reg_10_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_10_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_10_port, QN => n2257);
   DataP_PC_reg_O_reg_10_inst : DFF_X1 port map( D => DataP_PC_reg_N12, CK => 
                           Clk, Q => DataP_pc_out_10_port, QN => n_1292);
   DataP_IF_IDs_NPC_OUT_reg_11_inst : DFFRS_X1 port map( D => DataP_npc_11_port
                           , CK => Clk, RN => n82, SN => n83, Q => n_1293, QN 
                           => n84);
   DataP_ID_EXs_NPC_OUT_reg_11_inst : DFFS_X1 port map( D => n84, CK => Clk, SN
                           => Rst, Q => n81, QN => n_1294);
   DataP_EX_MEM_s_NPC_OUT_reg_11_inst : DFFS_X1 port map( D => n81, CK => Clk, 
                           SN => Rst, Q => n_1295, QN => DataP_npc_M_11_port);
   DataP_EX_MEM_s_ALU_OUT_reg_11_inst : DFFS_X1 port map( D => n2137, CK => Clk
                           , SN => Rst, Q => n2164, QN => DRAM_ADDRESS_11_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_11_inst : DFFR_X1 port map( D => 
                           DRAM_ADDRESS_11_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_11_port, QN => n2251);
   DataP_PC_reg_O_reg_11_inst : DFF_X1 port map( D => DataP_PC_reg_N13, CK => 
                           Clk, Q => DataP_pc_out_11_port, QN => n_1296);
   DataP_IF_IDs_NPC_OUT_reg_12_inst : DFFRS_X1 port map( D => DataP_npc_12_port
                           , CK => Clk, RN => n78, SN => n79, Q => n_1297, QN 
                           => n80);
   DataP_ID_EXs_NPC_OUT_reg_12_inst : DFFS_X1 port map( D => n80, CK => Clk, SN
                           => Rst, Q => n77, QN => n_1298);
   DataP_EX_MEM_s_NPC_OUT_reg_12_inst : DFFS_X1 port map( D => n77, CK => Clk, 
                           SN => Rst, Q => n_1299, QN => DataP_npc_M_12_port);
   DataP_EX_MEM_s_ALU_OUT_reg_12_inst : DFFS_X1 port map( D => n337, CK => Clk,
                           SN => Rst, Q => n2177, QN => DataP_alu_out_M_12_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_12_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_12_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_12_port, QN => n2246);
   DataP_PC_reg_O_reg_12_inst : DFF_X1 port map( D => DataP_PC_reg_N14, CK => 
                           Clk, Q => DataP_pc_out_12_port, QN => n_1300);
   DataP_IF_IDs_NPC_OUT_reg_13_inst : DFFRS_X1 port map( D => DataP_npc_13_port
                           , CK => Clk, RN => n74, SN => n75, Q => n_1301, QN 
                           => n76);
   DataP_ID_EXs_NPC_OUT_reg_13_inst : DFFS_X1 port map( D => n76, CK => Clk, SN
                           => Rst, Q => n73, QN => n_1302);
   DataP_EX_MEM_s_NPC_OUT_reg_13_inst : DFFS_X1 port map( D => n73, CK => Clk, 
                           SN => Rst, Q => n_1303, QN => DataP_npc_M_13_port);
   DataP_EX_MEM_s_ALU_OUT_reg_13_inst : DFFS_X1 port map( D => n333, CK => Clk,
                           SN => Rst, Q => n2176, QN => DataP_alu_out_M_13_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_13_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_13_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_13_port, QN => n2258);
   DataP_IF_IDs_NPC_OUT_reg_14_inst : DFFRS_X1 port map( D => DataP_npc_14_port
                           , CK => Clk, RN => n70, SN => n71, Q => n_1304, QN 
                           => n72);
   DataP_ID_EXs_NPC_OUT_reg_14_inst : DFFS_X1 port map( D => n72, CK => Clk, SN
                           => Rst, Q => n69, QN => n_1305);
   DataP_EX_MEM_s_NPC_OUT_reg_14_inst : DFFS_X1 port map( D => n69, CK => Clk, 
                           SN => Rst, Q => n_1306, QN => DataP_npc_M_14_port);
   DataP_EX_MEM_s_ALU_OUT_reg_14_inst : DFFS_X1 port map( D => n332, CK => Clk,
                           SN => Rst, Q => n2171, QN => DataP_alu_out_M_14_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_14_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_14_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_14_port, QN => n2252);
   DataP_PC_reg_O_reg_14_inst : DFF_X1 port map( D => DataP_PC_reg_N16, CK => 
                           Clk, Q => DataP_pc_out_14_port, QN => n_1307);
   DataP_IF_IDs_NPC_OUT_reg_15_inst : DFFRS_X1 port map( D => DataP_npc_15_port
                           , CK => Clk, RN => n66, SN => n67, Q => n_1308, QN 
                           => n68);
   DataP_ID_EXs_NPC_OUT_reg_15_inst : DFFS_X1 port map( D => n68, CK => Clk, SN
                           => Rst, Q => n65, QN => n_1309);
   DataP_EX_MEM_s_NPC_OUT_reg_15_inst : DFFS_X1 port map( D => n65, CK => Clk, 
                           SN => Rst, Q => n_1310, QN => DataP_npc_M_15_port);
   DataP_IF_IDs_NPC_OUT_reg_16_inst : DFFRS_X1 port map( D => DataP_npc_16_port
                           , CK => Clk, RN => n62, SN => n63, Q => n_1311, QN 
                           => n64);
   DataP_ID_EXs_NPC_OUT_reg_16_inst : DFFS_X1 port map( D => n64, CK => Clk, SN
                           => Rst, Q => n61, QN => n_1312);
   DataP_EX_MEM_s_NPC_OUT_reg_16_inst : DFFS_X1 port map( D => n61, CK => Clk, 
                           SN => Rst, Q => n_1313, QN => DataP_npc_M_16_port);
   DataP_EX_MEM_s_ALU_OUT_reg_16_inst : DFFS_X1 port map( D => n326, CK => Clk,
                           SN => Rst, Q => n2167, QN => DataP_alu_out_M_16_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_16_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_16_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_16_port, QN => n2263);
   DataP_PC_reg_O_reg_16_inst : DFF_X1 port map( D => DataP_PC_reg_N18, CK => 
                           Clk, Q => DataP_pc_out_16_port, QN => n_1314);
   DataP_IF_IDs_NPC_OUT_reg_17_inst : DFFRS_X1 port map( D => DataP_npc_17_port
                           , CK => Clk, RN => n58, SN => n59, Q => n_1315, QN 
                           => n60);
   DataP_ID_EXs_NPC_OUT_reg_17_inst : DFFS_X1 port map( D => n60, CK => Clk, SN
                           => Rst, Q => n57, QN => n_1316);
   DataP_EX_MEM_s_NPC_OUT_reg_17_inst : DFFS_X1 port map( D => n57, CK => Clk, 
                           SN => Rst, Q => n_1317, QN => DataP_npc_M_17_port);
   DataP_MEM_WB_s_ALU_OUT_reg_17_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_17_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_17_port, QN => n2248);
   DataP_PC_reg_O_reg_17_inst : DFF_X1 port map( D => DataP_PC_reg_N19, CK => 
                           Clk, Q => DataP_pc_out_17_port, QN => n_1318);
   DataP_IF_IDs_NPC_OUT_reg_18_inst : DFFRS_X1 port map( D => DataP_npc_18_port
                           , CK => Clk, RN => n54, SN => n55, Q => n_1319, QN 
                           => n56);
   DataP_ID_EXs_NPC_OUT_reg_18_inst : DFFS_X1 port map( D => n56, CK => Clk, SN
                           => Rst, Q => n53, QN => n_1320);
   DataP_EX_MEM_s_NPC_OUT_reg_18_inst : DFFS_X1 port map( D => n53, CK => Clk, 
                           SN => Rst, Q => n_1321, QN => DataP_npc_M_18_port);
   DataP_EX_MEM_s_ALU_OUT_reg_18_inst : DFFS_X1 port map( D => n322, CK => Clk,
                           SN => Rst, Q => n_1322, QN => 
                           DataP_alu_out_M_18_port);
   DataP_MEM_WB_s_ALU_OUT_reg_18_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_18_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_18_port, QN => n2259);
   DataP_PC_reg_O_reg_18_inst : DFF_X1 port map( D => DataP_PC_reg_N20, CK => 
                           Clk, Q => DataP_pc_out_18_port, QN => n_1323);
   DataP_IF_IDs_NPC_OUT_reg_19_inst : DFFRS_X1 port map( D => DataP_npc_19_port
                           , CK => Clk, RN => n50, SN => n51, Q => n_1324, QN 
                           => n52);
   DataP_ID_EXs_NPC_OUT_reg_19_inst : DFFS_X1 port map( D => n52, CK => Clk, SN
                           => Rst, Q => n49, QN => n_1325);
   DataP_EX_MEM_s_NPC_OUT_reg_19_inst : DFFS_X1 port map( D => n49, CK => Clk, 
                           SN => Rst, Q => n_1326, QN => DataP_npc_M_19_port);
   DataP_IF_IDs_NPC_OUT_reg_20_inst : DFFRS_X1 port map( D => DataP_npc_20_port
                           , CK => Clk, RN => n46, SN => n47, Q => n_1327, QN 
                           => n48);
   DataP_ID_EXs_NPC_OUT_reg_20_inst : DFFS_X1 port map( D => n48, CK => Clk, SN
                           => Rst, Q => n45, QN => n_1328);
   DataP_EX_MEM_s_NPC_OUT_reg_20_inst : DFFS_X1 port map( D => n45, CK => Clk, 
                           SN => Rst, Q => n_1329, QN => DataP_npc_M_20_port);
   DataP_EX_MEM_s_ALU_OUT_reg_20_inst : DFFS_X1 port map( D => n317, CK => Clk,
                           SN => Rst, Q => n2173, QN => DataP_alu_out_M_20_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_20_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_20_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_20_port, QN => n2260);
   DataP_PC_reg_O_reg_20_inst : DFF_X1 port map( D => DataP_PC_reg_N22, CK => 
                           Clk, Q => DataP_pc_out_20_port, QN => n_1330);
   DataP_IF_IDs_NPC_OUT_reg_21_inst : DFFRS_X1 port map( D => DataP_npc_21_port
                           , CK => Clk, RN => n42, SN => n43, Q => n_1331, QN 
                           => n44);
   DataP_ID_EXs_NPC_OUT_reg_21_inst : DFFS_X1 port map( D => n44, CK => Clk, SN
                           => Rst, Q => n41, QN => n_1332);
   DataP_EX_MEM_s_NPC_OUT_reg_21_inst : DFFS_X1 port map( D => n41, CK => Clk, 
                           SN => Rst, Q => n_1333, QN => DataP_npc_M_21_port);
   DataP_EX_MEM_s_ALU_OUT_reg_21_inst : DFFS_X1 port map( D => n313, CK => Clk,
                           SN => Rst, Q => n2172, QN => DataP_alu_out_M_21_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_21_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_21_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_21_port, QN => n2254);
   DataP_PC_reg_O_reg_21_inst : DFF_X1 port map( D => DataP_PC_reg_N23, CK => 
                           Clk, Q => DataP_pc_out_21_port, QN => n_1334);
   DataP_IF_IDs_NPC_OUT_reg_22_inst : DFFRS_X1 port map( D => DataP_npc_22_port
                           , CK => Clk, RN => n38, SN => n39, Q => n_1335, QN 
                           => n40);
   DataP_ID_EXs_NPC_OUT_reg_22_inst : DFFS_X1 port map( D => n40, CK => Clk, SN
                           => Rst, Q => n37, QN => n_1336);
   DataP_EX_MEM_s_NPC_OUT_reg_22_inst : DFFS_X1 port map( D => n37, CK => Clk, 
                           SN => Rst, Q => n_1337, QN => DataP_npc_M_22_port);
   DataP_MEM_WB_s_ALU_OUT_reg_22_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_22_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_22_port, QN => n2264);
   DataP_IF_IDs_NPC_OUT_reg_23_inst : DFFRS_X1 port map( D => DataP_npc_23_port
                           , CK => Clk, RN => n34, SN => n35, Q => n_1338, QN 
                           => n36);
   DataP_ID_EXs_NPC_OUT_reg_23_inst : DFFS_X1 port map( D => n36, CK => Clk, SN
                           => Rst, Q => n33, QN => n_1339);
   DataP_EX_MEM_s_NPC_OUT_reg_23_inst : DFFS_X1 port map( D => n33, CK => Clk, 
                           SN => Rst, Q => n_1340, QN => DataP_npc_M_23_port);
   DataP_IF_IDs_NPC_OUT_reg_24_inst : DFFRS_X1 port map( D => DataP_npc_24_port
                           , CK => Clk, RN => n30, SN => n31, Q => n_1341, QN 
                           => n32);
   DataP_ID_EXs_NPC_OUT_reg_24_inst : DFFS_X1 port map( D => n32, CK => Clk, SN
                           => Rst, Q => n29, QN => n_1342);
   DataP_EX_MEM_s_NPC_OUT_reg_24_inst : DFFS_X1 port map( D => n29, CK => Clk, 
                           SN => Rst, Q => n_1343, QN => DataP_npc_M_24_port);
   DataP_EX_MEM_s_ALU_OUT_reg_24_inst : DFFS_X1 port map( D => n308, CK => Clk,
                           SN => Rst, Q => n2179, QN => DataP_alu_out_M_24_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_24_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_24_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_24_port, QN => n2265);
   DataP_PC_reg_O_reg_24_inst : DFF_X1 port map( D => DataP_PC_reg_N26, CK => 
                           Clk, Q => DataP_pc_out_24_port, QN => n_1344);
   DataP_IF_IDs_NPC_OUT_reg_25_inst : DFFRS_X1 port map( D => DataP_npc_25_port
                           , CK => Clk, RN => n26, SN => n27, Q => n_1345, QN 
                           => n28);
   DataP_ID_EXs_NPC_OUT_reg_25_inst : DFFS_X1 port map( D => n28, CK => Clk, SN
                           => Rst, Q => n25, QN => n_1346);
   DataP_EX_MEM_s_NPC_OUT_reg_25_inst : DFFS_X1 port map( D => n25, CK => Clk, 
                           SN => Rst, Q => n_1347, QN => DataP_npc_M_25_port);
   DataP_EX_MEM_s_ALU_OUT_reg_25_inst : DFFS_X1 port map( D => n304, CK => Clk,
                           SN => Rst, Q => n2175, QN => DataP_alu_out_M_25_port
                           );
   DataP_MEM_WB_s_ALU_OUT_reg_25_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_25_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_25_port, QN => n2261);
   DataP_PC_reg_O_reg_25_inst : DFF_X1 port map( D => DataP_PC_reg_N27, CK => 
                           Clk, Q => DataP_pc_out_25_port, QN => n_1348);
   DataP_IF_IDs_NPC_OUT_reg_26_inst : DFFRS_X1 port map( D => DataP_npc_26_port
                           , CK => Clk, RN => n22, SN => n23, Q => n_1349, QN 
                           => n24);
   DataP_ID_EXs_NPC_OUT_reg_26_inst : DFFS_X1 port map( D => n24, CK => Clk, SN
                           => Rst, Q => n21, QN => n_1350);
   DataP_EX_MEM_s_NPC_OUT_reg_26_inst : DFFS_X1 port map( D => n21, CK => Clk, 
                           SN => Rst, Q => n_1351, QN => DataP_npc_M_26_port);
   DataP_MEM_WB_s_ALU_OUT_reg_26_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_26_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_26_port, QN => n2255);
   DataP_IF_IDs_NPC_OUT_reg_27_inst : DFFRS_X1 port map( D => DataP_npc_27_port
                           , CK => Clk, RN => n18, SN => n19, Q => n_1352, QN 
                           => n20);
   DataP_ID_EXs_NPC_OUT_reg_27_inst : DFFS_X1 port map( D => n20, CK => Clk, SN
                           => Rst, Q => n17, QN => n_1353);
   DataP_EX_MEM_s_NPC_OUT_reg_27_inst : DFFS_X1 port map( D => n17, CK => Clk, 
                           SN => Rst, Q => n_1354, QN => DataP_npc_M_27_port);
   DataP_IF_IDs_NPC_OUT_reg_28_inst : DFFRS_X1 port map( D => DataP_npc_28_port
                           , CK => Clk, RN => n14, SN => n15, Q => n_1355, QN 
                           => n16);
   DataP_ID_EXs_NPC_OUT_reg_28_inst : DFFS_X1 port map( D => n16, CK => Clk, SN
                           => Rst, Q => n13, QN => n_1356);
   DataP_EX_MEM_s_NPC_OUT_reg_28_inst : DFFS_X1 port map( D => n13, CK => Clk, 
                           SN => Rst, Q => n_1357, QN => DataP_npc_M_28_port);
   DataP_MEM_WB_s_ALU_OUT_reg_28_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_28_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_28_port, QN => n2262);
   DataP_IF_IDs_NPC_OUT_reg_29_inst : DFFRS_X1 port map( D => DataP_npc_29_port
                           , CK => Clk, RN => n10, SN => n11, Q => n_1358, QN 
                           => n12);
   DataP_ID_EXs_NPC_OUT_reg_29_inst : DFFS_X1 port map( D => n12, CK => Clk, SN
                           => Rst, Q => n9, QN => n_1359);
   DataP_EX_MEM_s_NPC_OUT_reg_29_inst : DFFS_X1 port map( D => n9, CK => Clk, 
                           SN => Rst, Q => n_1360, QN => DataP_npc_M_29_port);
   DataP_EX_MEM_s_ALU_OUT_reg_29_inst : DFFS_X1 port map( D => n299, CK => Clk,
                           SN => Rst, Q => n_1361, QN => 
                           DataP_alu_out_M_29_port);
   DataP_MEM_WB_s_ALU_OUT_reg_29_inst : DFFR_X1 port map( D => 
                           DataP_alu_out_M_29_port, CK => Clk, RN => Rst, Q => 
                           DataP_alu_out_W_29_port, QN => n2256);
   DataP_IF_IDs_NPC_OUT_reg_30_inst : DFFRS_X1 port map( D => DataP_npc_30_port
                           , CK => Clk, RN => n6, SN => n7, Q => n_1362, QN => 
                           n8);
   DataP_ID_EXs_NPC_OUT_reg_30_inst : DFFS_X1 port map( D => n8, CK => Clk, SN 
                           => Rst, Q => n5, QN => n_1363);
   DataP_EX_MEM_s_NPC_OUT_reg_30_inst : DFFS_X1 port map( D => n5, CK => Clk, 
                           SN => Rst, Q => n_1364, QN => DataP_npc_M_30_port);
   DataP_IF_IDs_NPC_OUT_reg_31_inst : DFFRS_X1 port map( D => DataP_npc_31_port
                           , CK => Clk, RN => n2, SN => n3, Q => n_1365, QN => 
                           n4);
   DataP_ID_EXs_NPC_OUT_reg_31_inst : DFFS_X1 port map( D => n4, CK => Clk, SN 
                           => Rst, Q => n1, QN => n_1366);
   DataP_EX_MEM_s_NPC_OUT_reg_31_inst : DFFS_X1 port map( D => n1, CK => Clk, 
                           SN => Rst, Q => n_1367, QN => DataP_npc_M_31_port);
   DataP_PC_reg_O_reg_27_inst : DFF_X1 port map( D => DataP_PC_reg_N29, CK => 
                           Clk, Q => DataP_pc_out_27_port, QN => n_1368);
   DataP_PC_reg_O_reg_23_inst : DFF_X1 port map( D => DataP_PC_reg_N25, CK => 
                           Clk, Q => DataP_pc_out_23_port, QN => n_1369);
   DataP_PC_reg_O_reg_7_inst : DFF_X1 port map( D => DataP_PC_reg_N9, CK => Clk
                           , Q => IRAM_ADDRESS_5_port, QN => n_1370);
   DataP_PC_reg_O_reg_0_inst : DFF_X1 port map( D => DataP_PC_reg_N2, CK => Clk
                           , Q => DataP_pc_out_0, QN => n_1371);
   sra_131_cell_849188 : AOI21_X1 port map( B1 => n2065, B2 => n2929, A => 
                           n2981, ZN => n2930);
   sra_131_cell_849192 : AOI21_X1 port map( B1 => n2065, B2 => n2925, A => 
                           n2981, ZN => n2926);
   sra_131_cell_849318 : AOI22_X1 port map( A1 => n2713, A2 => n2857, B1 => 
                           n2860, B2 => n2988, ZN => n2869);
   sra_131_cell_849321 : AOI22_X1 port map( A1 => n2713, A2 => n2855, B1 => 
                           n2858, B2 => n2988, ZN => n2866);
   sra_131_cell_849322 : AOI22_X1 port map( A1 => n2986, A2 => 
                           DataP_alu_a_in_21_port, B1 => DataP_alu_a_in_20_port
                           , B2 => n2985, ZN => n2858);
   sra_131_cell_849327 : AOI22_X1 port map( A1 => n2986, A2 => 
                           DataP_alu_a_in_25_port, B1 => DataP_alu_a_in_24_port
                           , B2 => n2985, ZN => n2856);
   sra_131_cell_849328 : AOI22_X1 port map( A1 => n2986, A2 => 
                           DataP_alu_a_in_27_port, B1 => DataP_alu_a_in_26_port
                           , B2 => n2985, ZN => n2853);
   sra_131_cell_849329 : AOI22_X1 port map( A1 => n2839, A2 => n2852, B1 => 
                           n2854, B2 => n2988, ZN => n2865);
   sra_131_cell_849331 : AOI22_X1 port map( A1 => n2986, A2 => 
                           DataP_alu_a_in_29_port, B1 => DataP_alu_a_in_28_port
                           , B2 => n2985, ZN => n2854);
   sra_131_cell_849332 : AOI22_X1 port map( A1 => n2986, A2 => 
                           DataP_alu_a_in_31_port, B1 => DataP_alu_a_in_30_port
                           , B2 => n2985, ZN => n2852);
   ashr_130_cell_849337 : AOI22_X1 port map( A1 => n1915, A2 => n2835, B1 => 
                           n2834, B2 => n2845, ZN => n2837);
   ashr_130_cell_849339 : AOI22_X1 port map( A1 => n1915, A2 => n2831, B1 => 
                           n2830, B2 => n2064, ZN => n2833);
   ashr_130_cell_849345 : AOI22_X1 port map( A1 => n2841, A2 => n2821, B1 => 
                           n2820, B2 => n1930, ZN => n2822);
   ashr_130_cell_849348 : AOI22_X1 port map( A1 => n2841, A2 => n2816, B1 => 
                           n2815, B2 => n1930, ZN => n2817);
   ashr_130_cell_849350 : AOI22_X1 port map( A1 => n1915, A2 => n2812, B1 => 
                           n2811, B2 => n2127, ZN => n2814);
   ashr_130_cell_849351 : AOI22_X1 port map( A1 => n2842, A2 => n2810, B1 => 
                           n2809, B2 => n1930, ZN => n2811);
   ashr_130_cell_849356 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => 
                           n2804, B1 => n2803, B2 => n1916, ZN => n2825);
   ashr_130_cell_849357 : NOR2_X1 port map( A1 => lt_x_134_B_4_port, A2 => 
                           n2802, ZN => DataP_ALU_C_shifter_N81);
   ashr_130_cell_849358 : NOR2_X1 port map( A1 => lt_x_134_B_4_port, A2 => 
                           n2801, ZN => DataP_ALU_C_shifter_N80);
   ashr_130_cell_849361 : AOI22_X1 port map( A1 => n2842, A2 => n2820, B1 => 
                           n2797, B2 => n1930, ZN => n2798);
   ashr_130_cell_849362 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => 
                           n2796, B1 => n2795, B2 => n1916, ZN => n2797);
   ashr_130_cell_849363 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => 
                           n2794, B1 => n2793, B2 => n1916, ZN => n2820);
   ashr_130_cell_849364 : AND2_X1 port map( A1 => n2792, A2 => n2847, ZN => 
                           DataP_ALU_C_shifter_N79);
   ashr_130_cell_849365 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => 
                           n2791, ZN => DataP_ALU_C_shifter_N78);
   ashr_130_cell_849366 : AND2_X1 port map( A1 => n2790, A2 => n2847, ZN => 
                           DataP_ALU_C_shifter_N77);
   ashr_130_cell_849367 : AND2_X1 port map( A1 => n2789, A2 => n2065, ZN => 
                           DataP_ALU_C_shifter_N76);
   ashr_130_cell_849368 : AND2_X1 port map( A1 => n2836, A2 => n2847, ZN => 
                           DataP_ALU_C_shifter_N75);
   ashr_130_cell_849419 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => 
                           n2747, B1 => n2746, B2 => n1916, ZN => n2763);
   ashr_130_cell_849420 : AOI22_X1 port map( A1 => n1915, A2 => n2779, B1 => 
                           n2818, B2 => n2845, ZN => n2748);
   ashr_130_cell_849421 : AOI22_X1 port map( A1 => n2842, A2 => n2764, B1 => 
                           n2771, B2 => n1930, ZN => n2818);
   ashr_130_cell_849422 : AOI22_X1 port map( A1 => n2839, A2 => n2745, B1 => 
                           n2744, B2 => n1916, ZN => n2771);
   ashr_130_cell_849423 : AOI22_X1 port map( A1 => n2839, A2 => n2743, B1 => 
                           n2742, B2 => n1916, ZN => n2764);
   ashr_130_cell_849424 : AOI22_X1 port map( A1 => n2842, A2 => n2762, B1 => 
                           n2765, B2 => n1930, ZN => n2779);
   ashr_130_cell_849425 : AOI22_X1 port map( A1 => n2839, A2 => n2741, B1 => 
                           n2740, B2 => n1916, ZN => n2765);
   ashr_130_cell_849426 : AOI22_X1 port map( A1 => n2839, A2 => n2739, B1 => 
                           n2738, B2 => n1916, ZN => n2762);
   ashr_130_cell_849427 : OAI21_X1 port map( B1 => n2847, B2 => n2791, A => 
                           n2737, ZN => DataP_ALU_C_shifter_N62);
   ashr_130_cell_849428 : NAND2_X1 port map( A1 => n2065, A2 => n2736, ZN => 
                           n2737);
   ashr_130_cell_849429 : AOI22_X1 port map( A1 => n1915, A2 => n2777, B1 => 
                           n2812, B2 => n2845, ZN => n2736);
   ashr_130_cell_849430 : AOI22_X1 port map( A1 => n2842, A2 => n2735, B1 => 
                           n2734, B2 => n1930, ZN => n2812);
   ashr_130_cell_849431 : AOI22_X1 port map( A1 => n2842, A2 => n2733, B1 => 
                           n2732, B2 => n1930, ZN => n2777);
   ashr_130_cell_849432 : NAND3_X1 port map( A1 => n2064, A2 => n1930, A3 => 
                           n2776, ZN => n2791);
   ashr_130_cell_849434 : MUX2_X1 port map( A => n2731, B => n2790, S => 
                           lt_x_135_B_4_port, Z => DataP_ALU_C_shifter_N61);
   ashr_130_cell_849435 : NOR2_X1 port map( A1 => n1915, A2 => n2769, ZN => 
                           n2790);
   ashr_130_cell_849436 : AOI22_X1 port map( A1 => n2842, A2 => n2784, B1 => 
                           n2756, B2 => n2844, ZN => n2769);
   ashr_130_cell_849437 : AOI22_X1 port map( A1 => n2839, A2 => n2746, B1 => 
                           n2739, B2 => n1916, ZN => n2756);
   ashr_130_cell_849438 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_28_port, B1 => DataP_alu_a_in_27_port
                           , B2 => n1931, ZN => n2739);
   ashr_130_cell_849439 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_30_port, B1 => DataP_alu_a_in_29_port
                           , B2 => n1931, ZN => n2746);
   ashr_130_cell_849440 : NOR2_X1 port map( A1 => n2840, A2 => n2747, ZN => 
                           n2784);
   ashr_130_cell_849441 : NAND2_X1 port map( A1 => DataP_alu_a_in_31_port, A2 
                           => n1931, ZN => n2747);
   ashr_130_cell_849442 : AOI22_X1 port map( A1 => n1915, A2 => n2768, B1 => 
                           n2807, B2 => n2845, ZN => n2731);
   ashr_130_cell_849443 : AOI22_X1 port map( A1 => n2842, A2 => n2757, B1 => 
                           n2826, B2 => n1930, ZN => n2807);
   ashr_130_cell_849444 : AOI22_X1 port map( A1 => n2839, A2 => n2744, B1 => 
                           n2770, B2 => n1916, ZN => n2826);
   ashr_130_cell_849445 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_12_port, B1 => DataP_alu_a_in_11_port
                           , B2 => n1931, ZN => n2770);
   ashr_130_cell_849446 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_14_port, B1 => DataP_alu_a_in_13_port
                           , B2 => n1931, ZN => n2744);
   ashr_130_cell_849447 : AOI22_X1 port map( A1 => n2839, A2 => n2742, B1 => 
                           n2745, B2 => n1916, ZN => n2757);
   ashr_130_cell_849448 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_16_port, B1 => n1841, B2 => n1931, ZN
                           => n2745);
   ashr_130_cell_849449 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_18_port, B1 => DataP_alu_a_in_17_port
                           , B2 => n1931, ZN => n2742);
   ashr_130_cell_849450 : AOI22_X1 port map( A1 => n2842, A2 => n2755, B1 => 
                           n2758, B2 => n2844, ZN => n2768);
   ashr_130_cell_849451 : AOI22_X1 port map( A1 => n2839, A2 => n2740, B1 => 
                           n2743, B2 => n1916, ZN => n2758);
   ashr_130_cell_849452 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_20_port, B1 => n1553, B2 => n1931, ZN
                           => n2743);
   ashr_130_cell_849453 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_22_port, B1 => DataP_alu_a_in_21_port
                           , B2 => n1931, ZN => n2740);
   ashr_130_cell_849454 : AOI22_X1 port map( A1 => n2839, A2 => n2738, B1 => 
                           n2741, B2 => n1916, ZN => n2755);
   ashr_130_cell_849455 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_24_port, B1 => DataP_alu_a_in_23_port
                           , B2 => n1931, ZN => n2741);
   ashr_130_cell_849456 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_26_port, B1 => DataP_alu_a_in_25_port
                           , B2 => n1931, ZN => n2738);
   ashr_130_cell_849457 : MUX2_X1 port map( A => n2730, B => n2789, S => 
                           lt_x_135_B_4_port, Z => DataP_ALU_C_shifter_N60);
   ashr_130_cell_849458 : NOR2_X1 port map( A1 => n1915, A2 => n2767, ZN => 
                           n2789);
   ashr_130_cell_849459 : AOI22_X1 port map( A1 => n2842, A2 => n2781, B1 => 
                           n2750, B2 => n2844, ZN => n2767);
   ashr_130_cell_849460 : AOI22_X1 port map( A1 => n2839, A2 => n2729, B1 => 
                           n2728, B2 => n1916, ZN => n2750);
   ashr_130_cell_849461 : NOR2_X1 port map( A1 => n2840, A2 => n2727, ZN => 
                           n2781);
   ashr_130_cell_849462 : AOI22_X1 port map( A1 => n1915, A2 => n2766, B1 => 
                           n2799, B2 => n2845, ZN => n2730);
   ashr_130_cell_849463 : AOI22_X1 port map( A1 => n2842, A2 => n2751, B1 => 
                           n2821, B2 => n2844, ZN => n2799);
   ashr_130_cell_849464 : AOI22_X1 port map( A1 => n2840, A2 => n2726, B1 => 
                           n2725, B2 => n1916, ZN => n2821);
   ashr_130_cell_849465 : AOI22_X1 port map( A1 => n2839, A2 => n2724, B1 => 
                           n2723, B2 => n1916, ZN => n2751);
   ashr_130_cell_849466 : AOI22_X1 port map( A1 => n2843, A2 => n2749, B1 => 
                           n2752, B2 => n2844, ZN => n2766);
   ashr_130_cell_849467 : AOI22_X1 port map( A1 => n2840, A2 => n2722, B1 => 
                           n2721, B2 => n1916, ZN => n2752);
   ashr_130_cell_849468 : AOI22_X1 port map( A1 => n2840, A2 => n2720, B1 => 
                           n2719, B2 => n1916, ZN => n2749);
   ashr_130_cell_849469 : MUX2_X1 port map( A => n2718, B => n2761, S => 
                           lt_x_135_B_4_port, Z => DataP_ALU_C_shifter_N50);
   ashr_130_cell_849470 : AOI22_X1 port map( A1 => n1915, A2 => n2787, B1 => 
                           n2831, B2 => n2845, ZN => n2761);
   ashr_130_cell_849471 : AOI22_X1 port map( A1 => n2843, A2 => n2732, B1 => 
                           n2735, B2 => n2844, ZN => n2831);
   ashr_130_cell_849472 : AOI22_X1 port map( A1 => n2840, A2 => n2721, B1 => 
                           n2724, B2 => n1916, ZN => n2735);
   ashr_130_cell_849473 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_17_port, B1 => DataP_alu_a_in_16_port
                           , B2 => n1931, ZN => n2724);
   ashr_130_cell_849474 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_19_port, B1 => DataP_alu_a_in_18_port
                           , B2 => n1931, ZN => n2721);
   ashr_130_cell_849475 : AOI22_X1 port map( A1 => n2840, A2 => n2719, B1 => 
                           n2722, B2 => n1916, ZN => n2732);
   ashr_130_cell_849476 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_21_port, B1 => DataP_alu_a_in_20_port
                           , B2 => n1931, ZN => n2722);
   ashr_130_cell_849477 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_23_port, B1 => DataP_alu_a_in_22_port
                           , B2 => n1931, ZN => n2719);
   ashr_130_cell_849478 : AOI22_X1 port map( A1 => n2843, A2 => n2776, B1 => 
                           n2733, B2 => n2844, ZN => n2787);
   ashr_130_cell_849479 : AOI22_X1 port map( A1 => n2840, A2 => n2728, B1 => 
                           n2720, B2 => n1916, ZN => n2733);
   ashr_130_cell_849480 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_25_port, B1 => DataP_alu_a_in_24_port
                           , B2 => n1931, ZN => n2720);
   ashr_130_cell_849481 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_27_port, B1 => DataP_alu_a_in_26_port
                           , B2 => n1931, ZN => n2728);
   ashr_130_cell_849482 : AOI22_X1 port map( A1 => n2840, A2 => n2727, B1 => 
                           n2729, B2 => n1916, ZN => n2776);
   ashr_130_cell_849483 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_29_port, B1 => DataP_alu_a_in_28_port
                           , B2 => n1931, ZN => n2729);
   ashr_130_cell_849484 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_31_port, B1 => DataP_alu_a_in_30_port
                           , B2 => n1931, ZN => n2727);
   ashr_130_cell_849485 : AOI22_X1 port map( A1 => n2846, A2 => n2830, B1 => 
                           n2717, B2 => n2064, ZN => n2718);
   ashr_130_cell_849487 : AOI21_X1 port map( B1 => n2841, B2 => n2809, A => 
                           n2716, ZN => n2717);
   ashr_130_cell_849488 : AOI221_X1 port map( B1 => n2795, B2 => n2839, C1 => 
                           n2715, C2 => n1916, A => n2841, ZN => n2716);
   ashr_130_cell_849489 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_1_port, B1 => n1605, B2 => n1931, ZN 
                           => n2715);
   ashr_130_cell_849490 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_3_port, B1 => DataP_alu_a_in_2_port, 
                           B2 => n1931, ZN => n2795);
   ashr_130_cell_849491 : AOI22_X1 port map( A1 => n2840, A2 => n2793, B1 => 
                           n2796, B2 => n1916, ZN => n2809);
   ashr_130_cell_849492 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_5_port, B1 => DataP_alu_a_in_4_port, 
                           B2 => n1931, ZN => n2796);
   ashr_130_cell_849493 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_7_port, B1 => DataP_alu_a_in_6_port, 
                           B2 => n1931, ZN => n2793);
   ashr_130_cell_849494 : AOI22_X1 port map( A1 => n2842, A2 => n2734, B1 => 
                           n2810, B2 => n1930, ZN => n2830);
   ashr_130_cell_849496 : AOI22_X1 port map( A1 => n2840, A2 => n2725, B1 => 
                           n2794, B2 => n1916, ZN => n2810);
   ashr_130_cell_849497 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_9_port, B1 => DataP_alu_a_in_8_port, 
                           B2 => n1931, ZN => n2794);
   ashr_130_cell_849498 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_11_port, B1 => DataP_alu_a_in_10_port
                           , B2 => n1931, ZN => n2725);
   ashr_130_cell_849499 : AOI22_X1 port map( A1 => n2839, A2 => n2723, B1 => 
                           n2726, B2 => n1916, ZN => n2734);
   ashr_130_cell_849501 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_13_port, B1 => DataP_alu_a_in_12_port
                           , B2 => n1931, ZN => n2726);
   ashr_130_cell_849502 : AOI22_X1 port map( A1 => n1914, A2 => 
                           DataP_alu_a_in_15_port, B1 => DataP_alu_a_in_14_port
                           , B2 => n1931, ZN => n2723);
   ash_129_cell_849520 : MUX2_X1 port map( A => n2689, B => n2688, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N49);
   ash_129_cell_849521 : AOI22_X1 port map( A1 => n2846, A2 => n2687, B1 => 
                           n2686, B2 => n2064, ZN => n2689);
   ash_129_cell_849522 : AOI22_X1 port map( A1 => n2714, A2 => n2685, B1 => 
                           n2684, B2 => n1930, ZN => n2686);
   ash_129_cell_849523 : AOI22_X1 port map( A1 => n2713, A2 => n2683, B1 => 
                           n2682, B2 => n1916, ZN => n2684);
   ash_129_cell_849524 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_30_port, B1 => DataP_alu_a_in_31_port
                           , B2 => n2711, ZN => n2682);
   ash_129_cell_849525 : MUX2_X1 port map( A => n2681, B => n2680, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N48);
   ash_129_cell_849526 : AOI22_X1 port map( A1 => n1915, A2 => n2679, B1 => 
                           n2678, B2 => n2845, ZN => n2681);
   ash_129_cell_849527 : AOI22_X1 port map( A1 => n2714, A2 => n2677, B1 => 
                           n2676, B2 => n2989, ZN => n2678);
   ash_129_cell_849528 : AOI22_X1 port map( A1 => n2713, A2 => n2675, B1 => 
                           n2674, B2 => n1916, ZN => n2676);
   ash_129_cell_849529 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_29_port, B1 => DataP_alu_a_in_30_port
                           , B2 => n2710, ZN => n2674);
   ash_129_cell_849532 : MUX2_X1 port map( A => n2672, B => n2671, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N47);
   ash_129_cell_849533 : AOI22_X1 port map( A1 => n1915, A2 => n2670, B1 => 
                           n2669, B2 => n2064, ZN => n2672);
   ash_129_cell_849534 : AOI22_X1 port map( A1 => n2714, A2 => n2668, B1 => 
                           n2667, B2 => n1913, ZN => n2669);
   ash_129_cell_849535 : AOI22_X1 port map( A1 => n2713, A2 => n2666, B1 => 
                           n2683, B2 => n1916, ZN => n2667);
   ash_129_cell_849536 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_28_port, B1 => DataP_alu_a_in_29_port
                           , B2 => n2711, ZN => n2683);
   ash_129_cell_849537 : MUX2_X1 port map( A => n2665, B => n2664, S => 
                           lt_x_135_B_4_port, Z => DataP_ALU_C_shifter_N46);
   ash_129_cell_849538 : AOI22_X1 port map( A1 => n1915, A2 => n2663, B1 => 
                           n2662, B2 => n2064, ZN => n2665);
   ash_129_cell_849539 : AOI22_X1 port map( A1 => n2714, A2 => n2661, B1 => 
                           n2660, B2 => n1930, ZN => n2662);
   ash_129_cell_849540 : AOI22_X1 port map( A1 => n2713, A2 => n2659, B1 => 
                           n2675, B2 => n1916, ZN => n2660);
   ash_129_cell_849541 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_27_port, B1 => DataP_alu_a_in_28_port
                           , B2 => n2711, ZN => n2675);
   ash_129_cell_849545 : AOI22_X1 port map( A1 => n2713, A2 => n2655, B1 => 
                           n2666, B2 => n1916, ZN => n2685);
   ash_129_cell_849546 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_26_port, B1 => DataP_alu_a_in_27_port
                           , B2 => n2711, ZN => n2666);
   ash_129_cell_849550 : AOI22_X1 port map( A1 => n2713, A2 => n2651, B1 => 
                           n2659, B2 => n1916, ZN => n2677);
   ash_129_cell_849551 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_25_port, B1 => DataP_alu_a_in_26_port
                           , B2 => n2711, ZN => n2659);
   ash_129_cell_849552 : MUX2_X1 port map( A => n2650, B => n2696, S => 
                           lt_x_135_B_4_port, Z => DataP_ALU_C_shifter_N43);
   ash_129_cell_849553 : AOI22_X1 port map( A1 => n1915, A2 => n2649, B1 => 
                           n2648, B2 => n2845, ZN => n2696);
   ash_129_cell_849554 : AOI22_X1 port map( A1 => n1915, A2 => n2647, B1 => 
                           n2646, B2 => n2845, ZN => n2650);
   ash_129_cell_849555 : AOI22_X1 port map( A1 => n2842, A2 => n2645, B1 => 
                           n2668, B2 => n1913, ZN => n2646);
   ash_129_cell_849556 : AOI22_X1 port map( A1 => n2713, A2 => n2644, B1 => 
                           n2655, B2 => n1916, ZN => n2668);
   ash_129_cell_849557 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_24_port, B1 => DataP_alu_a_in_25_port
                           , B2 => n2710, ZN => n2655);
   ash_129_cell_849558 : MUX2_X1 port map( A => n2643, B => n2695, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N42);
   ash_129_cell_849559 : AOI22_X1 port map( A1 => n1915, A2 => n2642, B1 => 
                           n2641, B2 => n2127, ZN => n2695);
   ash_129_cell_849560 : AOI22_X1 port map( A1 => n1915, A2 => n2640, B1 => 
                           n2639, B2 => n2845, ZN => n2643);
   ash_129_cell_849561 : AOI22_X1 port map( A1 => n2842, A2 => n2638, B1 => 
                           n2661, B2 => n1913, ZN => n2639);
   ash_129_cell_849562 : AOI22_X1 port map( A1 => n2713, A2 => n2637, B1 => 
                           n2651, B2 => n1916, ZN => n2661);
   ash_129_cell_849563 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_23_port, B1 => DataP_alu_a_in_24_port
                           , B2 => n2710, ZN => n2651);
   ash_129_cell_849565 : NOR2_X1 port map( A1 => n1915, A2 => n2636, ZN => 
                           n2694);
   ash_129_cell_849567 : AOI22_X1 port map( A1 => n2842, A2 => n2634, B1 => 
                           n2656, B2 => n1913, ZN => n2687);
   ash_129_cell_849568 : AOI22_X1 port map( A1 => n2713, A2 => n2633, B1 => 
                           n2644, B2 => n1916, ZN => n2656);
   ash_129_cell_849569 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_22_port, B1 => DataP_alu_a_in_23_port
                           , B2 => n2711, ZN => n2644);
   ash_129_cell_849570 : MUX2_X1 port map( A => n2632, B => n2693, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N40);
   ash_129_cell_849571 : NOR2_X1 port map( A1 => n1915, A2 => n2631, ZN => 
                           n2693);
   ash_129_cell_849572 : AOI22_X1 port map( A1 => n1915, A2 => n2630, B1 => 
                           n2679, B2 => n2127, ZN => n2632);
   ash_129_cell_849573 : AOI22_X1 port map( A1 => n2842, A2 => n2629, B1 => 
                           n2652, B2 => n1913, ZN => n2679);
   ash_129_cell_849574 : AOI22_X1 port map( A1 => n2839, A2 => n2628, B1 => 
                           n2637, B2 => n1916, ZN => n2652);
   ash_129_cell_849575 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_21_port, B1 => DataP_alu_a_in_22_port
                           , B2 => n2710, ZN => n2637);
   ash_129_cell_849577 : NOR2_X1 port map( A1 => n1915, A2 => n2627, ZN => 
                           n2692);
   ash_129_cell_849579 : AOI22_X1 port map( A1 => n2842, A2 => n2625, B1 => 
                           n2645, B2 => n1913, ZN => n2670);
   ash_129_cell_849580 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => 
                           n2624, B1 => n2633, B2 => n1916, ZN => n2645);
   ash_129_cell_849581 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_20_port, B1 => DataP_alu_a_in_21_port
                           , B2 => n2710, ZN => n2633);
   ash_129_cell_849582 : MUX2_X1 port map( A => n2623, B => n2691, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N38);
   ash_129_cell_849583 : NOR2_X1 port map( A1 => n1915, A2 => n2622, ZN => 
                           n2691);
   ash_129_cell_849584 : AOI22_X1 port map( A1 => n1915, A2 => n2621, B1 => 
                           n2663, B2 => n2330, ZN => n2623);
   ash_129_cell_849585 : AOI22_X1 port map( A1 => n2842, A2 => n2620, B1 => 
                           n2638, B2 => n1913, ZN => n2663);
   ash_129_cell_849586 : AOI22_X1 port map( A1 => n2839, A2 => n2619, B1 => 
                           n2628, B2 => n1916, ZN => n2638);
   ash_129_cell_849587 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_19_port, B1 => DataP_alu_a_in_20_port
                           , B2 => n2710, ZN => n2628);
   ash_129_cell_849588 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2703
                           , ZN => DataP_ALU_C_shifter_N19);
   ash_129_cell_849590 : MUX2_X1 port map( A => n2617, B => n2690, S => 
                           lt_x_134_B_4_port, Z => DataP_ALU_C_shifter_N37);
   ash_129_cell_849591 : NOR2_X1 port map( A1 => n1915, A2 => n2616, ZN => 
                           n2690);
   ash_129_cell_849592 : AOI22_X1 port map( A1 => n1915, A2 => n2615, B1 => 
                           n2657, B2 => n2845, ZN => n2617);
   ash_129_cell_849593 : AOI22_X1 port map( A1 => n2842, A2 => n2614, B1 => 
                           n2634, B2 => n1913, ZN => n2657);
   ash_129_cell_849594 : AOI22_X1 port map( A1 => n2840, A2 => n2613, B1 => 
                           n2624, B2 => n1916, ZN => n2634);
   ash_129_cell_849595 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_18_port, B1 => DataP_alu_a_in_19_port
                           , B2 => n2710, ZN => n2624);
   ash_129_cell_849597 : NOR2_X1 port map( A1 => n2846, A2 => n2612, ZN => 
                           n2673);
   ash_129_cell_849599 : AOI22_X1 port map( A1 => n2842, A2 => n2610, B1 => 
                           n2629, B2 => n1913, ZN => n2653);
   ash_129_cell_849600 : AOI22_X1 port map( A1 => n2839, A2 => n2609, B1 => 
                           n2619, B2 => n1916, ZN => n2629);
   ash_129_cell_849601 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_17_port, B1 => DataP_alu_a_in_18_port
                           , B2 => n2710, ZN => n2619);
   ash_129_cell_849603 : NOR2_X1 port map( A1 => n2846, A2 => n2649, ZN => 
                           n2618);
   ash_129_cell_849604 : NAND2_X1 port map( A1 => n2608, A2 => n1913, ZN => 
                           n2649);
   ash_129_cell_849606 : AOI22_X1 port map( A1 => n2842, A2 => n2607, B1 => 
                           n2625, B2 => n1913, ZN => n2647);
   ash_129_cell_849607 : AOI22_X1 port map( A1 => n2840, A2 => n2606, B1 => 
                           n2613, B2 => n1916, ZN => n2625);
   ash_129_cell_849608 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_16_port, B1 => DataP_alu_a_in_17_port
                           , B2 => n2710, ZN => n2613);
   ash_129_cell_849609 : AOI22_X1 port map( A1 => n2842, A2 => n2605, B1 => 
                           n2604, B2 => n1913, ZN => n2648);
   ash_129_cell_849610 : MUX2_X1 port map( A => n2603, B => n2602, S => 
                           lt_x_135_B_4_port, Z => DataP_ALU_C_shifter_N34);
   ash_129_cell_849611 : AOI22_X1 port map( A1 => n1915, A2 => n2641, B1 => 
                           n2640, B2 => n2845, ZN => n2603);
   ash_129_cell_849612 : AOI22_X1 port map( A1 => n2842, A2 => n2601, B1 => 
                           n2620, B2 => n1913, ZN => n2640);
   ash_129_cell_849613 : AOI22_X1 port map( A1 => n2840, A2 => n2600, B1 => 
                           n2609, B2 => n1916, ZN => n2620);
   ash_129_cell_849614 : AOI22_X1 port map( A1 => n2709, A2 => n1841, B1 => 
                           DataP_alu_a_in_16_port, B2 => n2710, ZN => n2609);
   ash_129_cell_849615 : AOI22_X1 port map( A1 => n2842, A2 => n2599, B1 => 
                           n2598, B2 => n1913, ZN => n2641);
   ash_129_cell_849616 : NOR2_X1 port map( A1 => lt_x_134_B_4_port, A2 => n2702
                           , ZN => DataP_ALU_C_shifter_N33);
   ash_129_cell_849618 : AOI22_X1 port map( A1 => n2846, A2 => n2636, B1 => 
                           n2635, B2 => n2127, ZN => n2688);
   ash_129_cell_849619 : AOI22_X1 port map( A1 => n2841, A2 => n2597, B1 => 
                           n2614, B2 => n1913, ZN => n2635);
   ash_129_cell_849620 : AOI22_X1 port map( A1 => n2839, A2 => n2596, B1 => 
                           n2606, B2 => n1916, ZN => n2614);
   ash_129_cell_849621 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_14_port, B1 => DataP_alu_a_in_15_port
                           , B2 => n2710, ZN => n2606);
   ash_129_cell_849622 : AOI22_X1 port map( A1 => n2841, A2 => n2595, B1 => 
                           n2594, B2 => n1913, ZN => n2636);
   ash_129_cell_849623 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2701
                           , ZN => DataP_ALU_C_shifter_N32);
   ash_129_cell_849625 : AOI22_X1 port map( A1 => n1915, A2 => n2631, B1 => 
                           n2630, B2 => n2845, ZN => n2680);
   ash_129_cell_849626 : AOI22_X1 port map( A1 => n2841, A2 => n2593, B1 => 
                           n2610, B2 => n2989, ZN => n2630);
   ash_129_cell_849627 : AOI22_X1 port map( A1 => n2839, A2 => n2592, B1 => 
                           n2600, B2 => n1916, ZN => n2610);
   ash_129_cell_849628 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_13_port, B1 => DataP_alu_a_in_14_port
                           , B2 => n2710, ZN => n2600);
   ash_129_cell_849629 : AOI22_X1 port map( A1 => n2841, A2 => n2591, B1 => 
                           n2590, B2 => n1913, ZN => n2631);
   ash_129_cell_849630 : NOR2_X1 port map( A1 => lt_x_134_B_4_port, A2 => n2700
                           , ZN => DataP_ALU_C_shifter_N31);
   ash_129_cell_849632 : AOI22_X1 port map( A1 => n2846, A2 => n2627, B1 => 
                           n2626, B2 => n2127, ZN => n2671);
   ash_129_cell_849633 : AOI22_X1 port map( A1 => n2841, A2 => n2604, B1 => 
                           n2607, B2 => n1913, ZN => n2626);
   ash_129_cell_849634 : AOI22_X1 port map( A1 => n2839, A2 => n2589, B1 => 
                           n2596, B2 => n1916, ZN => n2607);
   ash_129_cell_849635 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_12_port, B1 => DataP_alu_a_in_13_port
                           , B2 => n2710, ZN => n2596);
   ash_129_cell_849636 : AOI22_X1 port map( A1 => n2839, A2 => n2588, B1 => 
                           n2587, B2 => n1916, ZN => n2604);
   ash_129_cell_849637 : AOI22_X1 port map( A1 => n2841, A2 => n2608, B1 => 
                           n2605, B2 => n1913, ZN => n2627);
   ash_129_cell_849638 : AOI22_X1 port map( A1 => n2713, A2 => n2586, B1 => 
                           n2585, B2 => n1916, ZN => n2605);
   ash_129_cell_849639 : NOR2_X1 port map( A1 => n2713, A2 => n2584, ZN => 
                           n2608);
   ash_129_cell_849640 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2699
                           , ZN => DataP_ALU_C_shifter_N30);
   ash_129_cell_849642 : AOI22_X1 port map( A1 => n2846, A2 => n2622, B1 => 
                           n2621, B2 => n2064, ZN => n2664);
   ash_129_cell_849643 : AOI22_X1 port map( A1 => n2841, A2 => n2598, B1 => 
                           n2601, B2 => n1913, ZN => n2621);
   ash_129_cell_849644 : AOI22_X1 port map( A1 => n2713, A2 => n2583, B1 => 
                           n2592, B2 => n1916, ZN => n2601);
   ash_129_cell_849645 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_11_port, B1 => DataP_alu_a_in_12_port
                           , B2 => n2710, ZN => n2592);
   ash_129_cell_849646 : AOI22_X1 port map( A1 => n2713, A2 => n2582, B1 => 
                           n2581, B2 => n1916, ZN => n2598);
   ash_129_cell_849648 : AOI22_X1 port map( A1 => n2713, A2 => n2580, B1 => 
                           n2579, B2 => n1916, ZN => n2599);
   ash_129_cell_849650 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2698
                           , ZN => DataP_ALU_C_shifter_N29);
   ash_129_cell_849652 : AOI22_X1 port map( A1 => n2846, A2 => n2616, B1 => 
                           n2615, B2 => n2127, ZN => n2658);
   ash_129_cell_849653 : AOI22_X1 port map( A1 => n2842, A2 => n2594, B1 => 
                           n2597, B2 => n1913, ZN => n2615);
   ash_129_cell_849654 : AOI22_X1 port map( A1 => n2713, A2 => n2587, B1 => 
                           n2589, B2 => n1916, ZN => n2597);
   ash_129_cell_849655 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_10_port, B1 => DataP_alu_a_in_11_port
                           , B2 => n2710, ZN => n2589);
   ash_129_cell_849656 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_8_port, B1 => DataP_alu_a_in_9_port, 
                           B2 => n2711, ZN => n2587);
   ash_129_cell_849657 : AOI22_X1 port map( A1 => n2713, A2 => n2585, B1 => 
                           n2588, B2 => n1916, ZN => n2594);
   ash_129_cell_849658 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_6_port, B1 => DataP_alu_a_in_7_port, 
                           B2 => n2711, ZN => n2588);
   ash_129_cell_849659 : AOI22_X1 port map( A1 => n2709, A2 => 
                           DataP_alu_a_in_4_port, B1 => DataP_alu_a_in_5_port, 
                           B2 => n2711, ZN => n2585);
   DataP_MEM_WB_s_OPCODE_OUT_reg_5_inst : DFFS_X1 port map( D => n2161, CK => 
                           Clk, SN => Rst, Q => n3049, QN => 
                           DataP_opcode_W_5_port);
   DataP_ID_EXs_RS2_OUT_reg_1_inst : DFFS_X1 port map( D => n2559, CK => Clk, 
                           SN => Rst, Q => n_1372, QN => DataP_Rs2_1_port);
   DataP_ID_EXs_RS2_OUT_reg_0_inst : DFFS_X1 port map( D => n2558, CK => Clk, 
                           SN => Rst, Q => n1885, QN => DataP_Rs2_0_port);
   DataP_ID_EXs_RS2_OUT_reg_3_inst : DFFS_X1 port map( D => n2557, CK => Clk, 
                           SN => Rst, Q => n_1373, QN => DataP_Rs2_3_port);
   DataP_MEM_WB_s_RD_OUT_reg_1_inst : DFFS_X1 port map( D => n529, CK => Clk, 
                           SN => Rst, Q => n1891, QN => DataP_add_D_1_port);
   DataP_MEM_WB_s_RD_OUT_reg_3_inst : DFFS_X1 port map( D => n2570, CK => Clk, 
                           SN => Rst, Q => n2568, QN => DataP_add_D_3_port);
   DataP_IF_IDs_IR_OUT_reg_28_inst : DFFS_X2 port map( D => IRAM_DATA_OUT(28), 
                           CK => Clk, SN => n164, Q => IR_CU_28, QN => n510);
   DataP_IF_IDs_IR_OUT_reg_30_inst : DFFS_X1 port map( D => IRAM_DATA_OUT(30), 
                           CK => Clk, SN => n164, Q => n2129, QN => n515);
   DataP_PC_reg_O_reg_29_inst : DFF_X2 port map( D => DataP_PC_reg_N31, CK => 
                           Clk, Q => DataP_pc_out_29_port, QN => n_1374);
   lt_x_134_cell_849092 : AOI21_X1 port map( B1 => DataP_alu_a_in_4_port, B2 =>
                           n2847, A => n2023, ZN => n2024);
   lt_x_134_cell_849116 : NOR2_X1 port map( A1 => n1572, A2 => n1863, ZN => 
                           n2028);
   lt_x_134_cell_849143 : NAND2_X1 port map( A1 => DataP_alu_b_in_31_port, A2 
                           => n1923, ZN => n2013);
   DataP_PC_reg_O_reg_30_inst : DFF_X2 port map( D => DataP_PC_reg_N32, CK => 
                           Clk, Q => DataP_pc_out_30_port, QN => n_1375);
   DataP_EX_MEM_s_ALU_OUT_reg_26_inst : DFFS_X2 port map( D => n1599, CK => Clk
                           , SN => Rst, Q => n2169, QN => 
                           DataP_alu_out_M_26_port);
   DataP_EX_MEM_s_ALU_OUT_reg_31_inst : DFFS_X1 port map( D => n297, CK => Clk,
                           SN => Rst, Q => n2185, QN => DataP_alu_out_M_31_port
                           );
   DataP_EX_MEM_s_RD_OUT_reg_0_inst : DFFR_X1 port map( D => n1956, CK => Clk, 
                           RN => Rst, Q => DataP_dest_M_0_port, QN => n528);
   DataP_MEM_WB_s_RD_OUT_reg_2_inst : DFFR_X1 port map( D => 
                           DataP_dest_M_2_port, CK => Clk, RN => Rst, Q => 
                           DataP_add_D_2_port, QN => n538);
   DataP_PC_reg_O_reg_31_inst : DFF_X1 port map( D => DataP_PC_reg_N33, CK => 
                           Clk, Q => DataP_pc_out_31_port, QN => n_1376);
   CU_I_cw1_reg_4_inst : DFFR_X1 port map( D => CU_I_cw_4_port, CK => Clk, RN 
                           => Rst, Q => n_1377, QN => n132);
   CU_I_cw1_reg_6_inst : DFFR_X1 port map( D => CU_I_cw_6_port, CK => Clk, RN 
                           => Rst, Q => n_1378, QN => n130);
   CU_I_cw1_reg_3_inst : DFFR_X1 port map( D => CU_I_cw_3_port, CK => Clk, RN 
                           => Rst, Q => n_1379, QN => n131);
   CU_I_cw1_reg_7_inst : DFFR_X1 port map( D => CU_I_cw_7_port, CK => Clk, RN 
                           => Rst, Q => n_1380, QN => n143);
   CU_I_cw1_reg_1_inst : DFFR_X1 port map( D => CU_I_cw_1_port, CK => Clk, RN 
                           => Rst, Q => n_1381, QN => n129);
   CU_I_cw1_reg_0_inst : DFFR_X1 port map( D => CU_I_cw_0_port, CK => Clk, RN 
                           => Rst, Q => n_1382, QN => n136);
   DataP_ID_EXs_RD_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_dest_D_4_port,
                           CK => Clk, RN => Rst, Q => n_1383, QN => n142);
   DataP_ID_EXs_RD_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_dest_D_3_port,
                           CK => Clk, RN => Rst, Q => n_1384, QN => n141);
   DataP_ID_EXs_RD_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_dest_D_2_port,
                           CK => Clk, RN => Rst, Q => n_1385, QN => n140);
   DataP_ID_EXs_RD_OUT_reg_1_inst : DFFR_X1 port map( D => DataP_dest_D_1_port,
                           CK => Clk, RN => Rst, Q => n_1386, QN => n139);
   DataP_ID_EXs_RD_OUT_reg_0_inst : DFFR_X1 port map( D => DataP_dest_D_0_port,
                           CK => Clk, RN => Rst, Q => n1956, QN => n_1387);
   DataP_IF_IDs_PR_OUT_reg : DFFR_X1 port map( D => DataP_prediction, CK => 
                           DataP_IF_IDs_net834167, RN => Rst, Q => n_1388, QN 
                           => n258);
   DataP_ID_EXs_RS1_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_IR1_24_port, 
                           CK => Clk, RN => Rst, Q => n_1389, QN => n523);
   DataP_PC_reg_O_reg_13_inst : DFFRS_X1 port map( D => DataP_PC_reg_N15, CK =>
                           Clk, RN => n1874, SN => n1874, Q => 
                           DataP_pc_out_13_port, QN => n_1390);
   DataP_EX_MEM_s_ALU_OUT_reg_17_inst : DFFS_X2 port map( D => n1604, CK => Clk
                           , SN => Rst, Q => n2170, QN => 
                           DataP_alu_out_M_17_port);
   DataP_ID_EXs_RS2_OUT_reg_4_inst : DFFS_X1 port map( D => n1872, CK => Clk, 
                           SN => Rst, Q => n_1391, QN => DataP_Rs2_4_port);
   DataP_ID_EXs_RS1_OUT_reg_1_inst : DFFS_X1 port map( D => n153, CK => Clk, SN
                           => Rst, Q => n2160, QN => DataP_Rs1_1_port);
   DataP_ID_EXs_OPCODE_OUT_reg_0_inst : DFFS_X1 port map( D => n497, CK => Clk,
                           SN => Rst, Q => n151, QN => DataP_opcode_E_0_port);
   DataP_EX_MEM_s_ALU_OUT_reg_19_inst : DFFS_X1 port map( D => n319, CK => Clk,
                           SN => Rst, Q => n2174, QN => DataP_alu_out_M_19_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_15_inst : DFFS_X1 port map( D => n330, CK => Clk,
                           SN => Rst, Q => n2166, QN => DataP_alu_out_M_15_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_30_inst : DFFS_X1 port map( D => n2567, CK => Clk
                           , SN => Rst, Q => n2187, QN => 
                           DataP_alu_out_M_30_port);
   DataP_ID_EXs_OPCODE_OUT_reg_1_inst : DFFS_X1 port map( D => n504, CK => Clk,
                           SN => Rst, Q => n520, QN => n2573);
   DataP_EX_MEM_s_OPCODE_OUT_reg_4_inst : DFFS_X1 port map( D => n147, CK => 
                           Clk, SN => Rst, Q => n146, QN => 
                           DataP_opcode_M_4_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_0_inst : DFFS_X1 port map( D => n151, CK => 
                           Clk, SN => Rst, Q => n150, QN => 
                           DataP_opcode_M_0_port);
   DataP_ID_EXs_RS1_OUT_reg_0_inst : DFFR_X1 port map( D => DataP_IR1_21_port, 
                           CK => Clk, RN => Rst, Q => n_1392, QN => n2154);
   DataP_PC_reg_O_reg_15_inst : DFF_X2 port map( D => DataP_PC_reg_N17, CK => 
                           Clk, Q => DataP_pc_out_15_port, QN => n_1393);
   DataP_PC_reg_O_reg_19_inst : DFF_X1 port map( D => DataP_PC_reg_N21, CK => 
                           Clk, Q => DataP_pc_out_19_port, QN => n_1394);
   DataP_EX_MEM_s_ALU_OUT_reg_23_inst : DFFS_X2 port map( D => n1549, CK => Clk
                           , SN => Rst, Q => n2168, QN => 
                           DataP_alu_out_M_23_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_2_inst : DFFS_X1 port map( D => n1543, CK => 
                           Clk, SN => Rst, Q => n1545, QN => 
                           DataP_opcode_W_2_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_2_inst : DFFR_X1 port map( D => n2574, CK => 
                           Clk, RN => Rst, Q => n1895, QN => n1894);
   DataP_PC_reg_O_reg_28_inst : DFF_X1 port map( D => DataP_PC_reg_N30, CK => 
                           Clk, Q => DataP_pc_out_28_port, QN => n_1395);
   DataP_EX_MEM_s_ALU_OUT_reg_28_inst : DFFS_X2 port map( D => n1540, CK => Clk
                           , SN => Rst, Q => n2178, QN => 
                           DataP_alu_out_M_28_port);
   DataP_PC_reg_O_reg_26_inst : DFF_X2 port map( D => DataP_PC_reg_N28, CK => 
                           Clk, Q => DataP_pc_out_26_port, QN => n_1396);
   DataP_MEM_WB_s_OPCODE_OUT_reg_1_inst : DFFS_X1 port map( D => n2576, CK => 
                           Clk, SN => Rst, Q => n2571, QN => 
                           DataP_opcode_W_1_port);
   DataP_PC_reg_O_reg_22_inst : DFFRS_X2 port map( D => DataP_PC_reg_N24, CK =>
                           Clk, RN => n1873, SN => n1873, Q => 
                           DataP_pc_out_22_port, QN => n_1397);
   DataP_EX_MEM_s_ALU_OUT_reg_22_inst : DFFS_X2 port map( D => n1519, CK => Clk
                           , SN => Rst, Q => n2180, QN => 
                           DataP_alu_out_M_22_port);
   U1451 : BUF_X1 port map( A => n2564, Z => n1515);
   U1452 : AND2_X2 port map( A1 => DataP_alu_a_in_0_port, A2 => n1537, ZN => 
                           n3361);
   U1453 : AND3_X2 port map( A1 => n3329, A2 => n3046, A3 => n2189, ZN => n3328
                           );
   U1454 : INV_X4 port map( A => n2712, ZN => n2710);
   U1455 : INV_X1 port map( A => n3496, ZN => n1516);
   U1456 : BUF_X1 port map( A => n1886, Z => n1517);
   U1457 : AND3_X2 port map( A1 => n3329, A2 => n3046, A3 => n399, ZN => n1518)
                           ;
   U1458 : AND3_X1 port map( A1 => n3329, A2 => n3046, A3 => n399, ZN => n3327)
                           ;
   U1459 : BUF_X1 port map( A => n311, Z => n1519);
   U1460 : NAND2_X1 port map( A1 => n3458, A2 => n2299, ZN => n1520);
   U1461 : AND2_X1 port map( A1 => n1669, A2 => n1594, ZN => n1521);
   U1462 : AND4_X1 port map( A1 => n1586, A2 => n1521, A3 => n3281, A4 => n3291
                           , ZN => n1522);
   U1463 : OR2_X1 port map( A1 => n3910, A2 => n3990, ZN => n1523);
   U1464 : INV_X2 port map( A => n3689, ZN => n3510);
   U1465 : AND4_X1 port map( A1 => n3095, A2 => n3093, A3 => n3092, A4 => n3094
                           , ZN => n1524);
   U1466 : AND2_X1 port map( A1 => n3105, A2 => n3106, ZN => n1525);
   U1467 : AND2_X1 port map( A1 => n3307, A2 => n3308, ZN => n1526);
   U1468 : OR2_X1 port map( A1 => n3194, A2 => n2213, ZN => n1527);
   U1469 : INV_X2 port map( A => n1561, ZN => DataP_alu_a_in_2_port);
   U1470 : AND3_X2 port map( A1 => n1868, A2 => n3111, A3 => n1527, ZN => n1561
                           );
   U1471 : BUF_X1 port map( A => n2403, Z => n1528);
   U1472 : BUF_X2 port map( A => n3330, Z => n3005);
   U1473 : OAI211_X1 port map( C1 => n1636, C2 => n2185, A => n3306, B => n1809
                           , ZN => DataP_alu_b_in_31_port);
   U1474 : AOI211_X1 port map( C1 => n2055, C2 => n1772, A => n1773, B => n1774
                           , ZN => n2119);
   U1475 : BUF_X1 port map( A => n2542, Z => n1529);
   U1476 : BUF_X1 port map( A => n3330, Z => n3004);
   U1477 : AOI21_X1 port map( B1 => n3001, B2 => DataP_B_s_14_port, A => n1671,
                           ZN => n1530);
   U1478 : AND2_X1 port map( A1 => n2296, A2 => DataP_alu_a_in_18_port, ZN => 
                           n1531);
   U1479 : INV_X1 port map( A => n1863, ZN => DataP_alu_a_in_11_port);
   U1480 : OR2_X4 port map( A1 => n3143, A2 => n3142, ZN => 
                           DataP_alu_a_in_27_port);
   U1481 : INV_X2 port map( A => n1603, ZN => DataP_alu_b_in_6_port);
   U1482 : INV_X1 port map( A => n2571, ZN => n1532);
   U1483 : INV_X2 port map( A => n2712, ZN => n2711);
   U1484 : BUF_X2 port map( A => n2004, Z => n2712);
   U1485 : AND2_X1 port map( A1 => n3578, A2 => n3580, ZN => n1533);
   U1486 : NAND3_X1 port map( A1 => n3310, A2 => n3309, A3 => n1526, ZN => 
                           DataP_alu_b_in_13_port);
   U1487 : AND2_X1 port map( A1 => n1615, A2 => n149, ZN => n1616);
   U1488 : XOR2_X1 port map( A => DataP_Rs2_4_port, B => n2569, Z => n1534);
   U1489 : AND2_X1 port map( A1 => n147, A2 => n145, ZN => n1618);
   U1490 : AND2_X2 port map( A1 => n151, A2 => n521, ZN => n1619);
   U1491 : NAND4_X1 port map( A1 => n1616, A2 => n1534, A3 => n1618, A4 => 
                           n1619, ZN => n1535);
   U1492 : NOR2_X1 port map( A1 => n2157, A2 => n1535, ZN => n1617);
   U1493 : INV_X1 port map( A => n1619, ZN => n3031);
   U1494 : NAND2_X1 port map( A1 => n3381, A2 => n3377, ZN => n1536);
   U1495 : AOI21_X1 port map( B1 => n3205, B2 => n3676, A => n1536, ZN => n1886
                           );
   U1496 : OAI211_X1 port map( C1 => n1886, C2 => n3212, A => n3211, B => n3387
                           , ZN => n3269);
   U1497 : NAND4_X1 port map( A1 => n1542, A2 => n3089, A3 => n3091, A4 => 
                           n3088, ZN => n1537);
   U1498 : NAND2_X1 port map( A1 => n1538, A2 => n1553, ZN => n1552);
   U1499 : OR2_X1 port map( A1 => n1538, A2 => DataP_alu_a_in_19_port, ZN => 
                           n2378);
   U1500 : NAND2_X1 port map( A1 => n1699, A2 => n1700, ZN => n1538);
   U1501 : NAND4_X1 port map( A1 => n2332, A2 => n1584, A3 => n2336, A4 => 
                           n1585, ZN => DataP_alu_b_in_8_port);
   U1502 : BUF_X2 port map( A => n2560, Z => n1539);
   U1503 : BUF_X1 port map( A => n2560, Z => n2562);
   U1504 : BUF_X1 port map( A => n300, Z => n1540);
   U1505 : BUF_X1 port map( A => n3455, Z => n1541);
   U1506 : BUF_X1 port map( A => n3090, Z => n1542);
   U1507 : BUF_X1 port map( A => n1894, Z => n1543);
   U1508 : BUF_X1 port map( A => n2008, Z => n1544);
   U1509 : INV_X1 port map( A => n1545, ZN => n1546);
   U1510 : INV_X1 port map( A => n2467, ZN => n1547);
   U1511 : BUF_X1 port map( A => n3506, Z => n1548);
   U1512 : OAI211_X1 port map( C1 => n2566, C2 => n2175, A => n3306, B => n1721
                           , ZN => DataP_alu_b_in_25_port);
   U1513 : AOI21_X1 port map( B1 => n1541, B2 => n3691, A => n3454, ZN => n1549
                           );
   U1514 : AND4_X2 port map( A1 => n3322, A2 => n3321, A3 => n3320, A4 => n3319
                           , ZN => n1550);
   U1515 : INV_X4 port map( A => n1550, ZN => DataP_alu_b_in_24_port);
   U1516 : NAND2_X1 port map( A1 => n3427, A2 => n3510, ZN => n1551);
   U1517 : INV_X2 port map( A => n1945, ZN => n1553);
   U1518 : AND3_X1 port map( A1 => n1620, A2 => n2314, A3 => n1617, ZN => n1554
                           );
   U1519 : AND4_X1 port map( A1 => n3063, A2 => n3062, A3 => n3027, A4 => n3028
                           , ZN => n1555);
   U1520 : AND4_X1 port map( A1 => n3063, A2 => n3062, A3 => n3027, A4 => n3028
                           , ZN => n3029);
   U1521 : AND4_X1 port map( A1 => n3288, A2 => n3287, A3 => n3286, A4 => n3285
                           , ZN => n1556);
   U1522 : INV_X2 port map( A => n1556, ZN => DataP_alu_b_in_20_port);
   U1523 : AND3_X1 port map( A1 => n1620, A2 => n2314, A3 => n1617, ZN => n2313
                           );
   U1524 : NAND2_X1 port map( A1 => n1551, A2 => n1558, ZN => n1557);
   U1525 : AND2_X1 port map( A1 => n1884, A2 => n2297, ZN => n1558);
   U1526 : AND2_X1 port map( A1 => n2378, A2 => n1552, ZN => n1559);
   U1527 : AND2_X1 port map( A1 => n2378, A2 => n1552, ZN => n1877);
   U1528 : AND2_X2 port map( A1 => n3424, A2 => n3425, ZN => n2245);
   U1529 : NAND2_X1 port map( A1 => n2007, A2 => DataP_alu_a_in_20_port, ZN => 
                           n1560);
   U1530 : OAI21_X1 port map( B1 => n1567, B2 => n121, A => n3115, ZN => n1562)
                           ;
   U1531 : OR2_X2 port map( A1 => n1562, A2 => n3116, ZN => 
                           DataP_alu_a_in_1_port);
   U1532 : AND2_X2 port map( A1 => n3420, A2 => n3421, ZN => n1563);
   U1533 : AND4_X1 port map( A1 => n3305, A2 => n2519, A3 => n3303, A4 => n3304
                           , ZN => n1580);
   U1534 : OR2_X2 port map( A1 => n3184, A2 => n3183, ZN => 
                           DataP_alu_a_in_13_port);
   U1535 : INV_X2 port map( A => n2005, ZN => n3002);
   U1536 : AND2_X2 port map( A1 => n2315, A2 => n1554, ZN => n2005);
   U1537 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_0_port, ZN => n1564)
                           ;
   U1538 : NAND4_X1 port map( A1 => n1861, A2 => n3030, A3 => n2472, A4 => 
                           n2471, ZN => n1565);
   U1539 : NAND4_X1 port map( A1 => n1861, A2 => n3030, A3 => n2472, A4 => 
                           n2471, ZN => n3046);
   U1540 : NAND3_X1 port map( A1 => n3029, A2 => n2472, A3 => n3030, ZN => 
                           n1566);
   U1541 : NOR2_X2 port map( A1 => n1596, A2 => n1595, ZN => n3030);
   U1542 : NAND3_X1 port map( A1 => n1568, A2 => n2998, A3 => n2155, ZN => 
                           n1567);
   U1543 : INV_X1 port map( A => n3191, ZN => n1568);
   U1544 : AND3_X2 port map( A1 => n3104, A2 => n1525, A3 => n3107, ZN => n1569
                           );
   U1545 : INV_X2 port map( A => DataP_alu_b_in_8_port, ZN => n3663);
   U1546 : NAND2_X2 port map( A1 => n1570, A2 => n1571, ZN => n1572);
   U1547 : AND2_X1 port map( A1 => n3244, A2 => n3245, ZN => n1570);
   U1548 : AND2_X1 port map( A1 => n3246, A2 => n3247, ZN => n1571);
   U1549 : OR2_X2 port map( A1 => n3155, A2 => n3154, ZN => 
                           DataP_alu_a_in_23_port);
   U1550 : AOI211_X1 port map( C1 => DataP_alu_a_in_28_port, C2 => n1917, A => 
                           n2067, B => n2048, ZN => n1573);
   U1551 : INV_X1 port map( A => n1575, ZN => n3104);
   U1552 : AND2_X1 port map( A1 => n3004, A2 => DataP_alu_out_W_5_port, ZN => 
                           n1575);
   U1553 : AOI21_X1 port map( B1 => n2325, B2 => n2130, A => n1948, ZN => n1574
                           );
   U1554 : CLKBUF_X3 port map( A => DataP_alu_b_in_5_port, Z => 
                           lt_x_134_B_5_port);
   U1555 : AOI211_X4 port map( C1 => n2047, C2 => n2107, A => n2105, B => n1810
                           , ZN => n2057);
   U1556 : NAND2_X1 port map( A1 => n1576, A2 => n3048, ZN => n2389);
   U1557 : AND2_X1 port map( A1 => n3047, A2 => n2391, ZN => n1576);
   U1558 : AND2_X2 port map( A1 => n1900, A2 => n1637, ZN => n1577);
   U1559 : AND2_X2 port map( A1 => n1578, A2 => n1579, ZN => n3417);
   U1560 : AND3_X1 port map( A1 => n3301, A2 => n3300, A3 => n3302, ZN => n1578
                           );
   U1561 : NAND2_X1 port map( A1 => n1839, A2 => DataP_B_s_15_port, ZN => n1579
                           );
   U1562 : NAND4_X1 port map( A1 => n3095, A2 => n3093, A3 => n3092, A4 => 
                           n3094, ZN => n1581);
   U1563 : NAND2_X1 port map( A1 => n1584, A2 => n1583, ZN => n1582);
   U1564 : AND2_X1 port map( A1 => n1585, A2 => n2332, ZN => n1583);
   U1565 : NAND2_X1 port map( A1 => n2331, A2 => DRAM_ADDRESS_8_port, ZN => 
                           n1584);
   U1566 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_8_port, ZN => n1585)
                           ;
   U1567 : BUF_X4 port map( A => n2712, Z => n2709);
   U1568 : NAND2_X2 port map( A1 => n3224, A2 => n3343, ZN => n3689);
   U1569 : NOR2_X2 port map( A1 => ALU_OPCODE_i_3_port, A2 => 
                           ALU_OPCODE_i_0_port, ZN => n3343);
   U1570 : AND3_X2 port map( A1 => n2442, A2 => n1994, A3 => n2010, ZN => n3421
                           );
   U1571 : OR2_X2 port map( A1 => n3164, A2 => n3163, ZN => 
                           DataP_alu_a_in_20_port);
   U1572 : AND3_X2 port map( A1 => n1998, A2 => n3460, A3 => n3457, ZN => n3494
                           );
   U1573 : INV_X1 port map( A => n2145, ZN => n1586);
   U1574 : NAND2_X1 port map( A1 => n1993, A2 => n3678, ZN => n1587);
   U1575 : OR2_X2 port map( A1 => n3149, A2 => n3148, ZN => 
                           DataP_alu_a_in_25_port);
   U1576 : OR2_X2 port map( A1 => n3003, A2 => n2234, ZN => n3089);
   U1577 : AND2_X1 port map( A1 => n3021, A2 => n3022, ZN => n1588);
   U1578 : NOR2_X1 port map( A1 => n3161, A2 => n3160, ZN => n1589);
   U1579 : AND4_X1 port map( A1 => n3087, A2 => n3085, A3 => n3086, A4 => n3084
                           , ZN => n1907);
   U1580 : NAND3_X1 port map( A1 => n3101, A2 => n3100, A3 => n3102, ZN => 
                           n1625);
   U1581 : OR2_X1 port map( A1 => n2389, A2 => n1846, ZN => 
                           DataP_alu_b_in_9_port);
   U1582 : XOR2_X1 port map( A => n3011, B => n3203, Z => n1957);
   U1583 : BUF_X1 port map( A => n3532, Z => n1590);
   U1584 : BUF_X1 port map( A => n1531, Z => n1591);
   U1585 : NOR3_X1 port map( A1 => n1582, A2 => n2389, A3 => n2333, ZN => n1592
                           );
   U1586 : AND2_X2 port map( A1 => n1569, A2 => n1843, ZN => n1994);
   U1587 : NAND2_X2 port map( A1 => n3464, A2 => DataP_alu_a_in_23_port, ZN => 
                           n3497);
   U1588 : BUF_X2 port map( A => DataP_alu_b_in_12_port, Z => n1880);
   U1589 : NOR2_X2 port map( A1 => n3639, A2 => n1962, ZN => n2225);
   U1590 : OAI21_X1 port map( B1 => n309, B2 => n3911, A => n1593, ZN => 
                           DataP_PC_reg_N25);
   U1591 : OR2_X1 port map( A1 => n3910, A2 => n4013, ZN => n1593);
   U1592 : OAI21_X2 port map( B1 => n2434, B2 => n3911, A => n1523, ZN => n2346
                           );
   U1593 : BUF_X2 port map( A => n3327, Z => n1839);
   U1594 : NAND3_X1 port map( A1 => n1555, A2 => n2472, A3 => n3030, ZN => 
                           n2315);
   U1595 : NOR2_X1 port map( A1 => n3024, A2 => n3025, ZN => n3028);
   U1596 : NAND3_X1 port map( A1 => n1994, A2 => n2442, A3 => n1903, ZN => 
                           n2440);
   U1597 : AND3_X1 port map( A1 => n3067, A2 => n3066, A3 => n432, ZN => n2143)
                           ;
   U1598 : AND4_X2 port map( A1 => n1577, A2 => n2501, A3 => n1569, A4 => n1624
                           , ZN => n3207);
   U1599 : NAND2_X1 port map( A1 => n2331, A2 => DataP_alu_out_M_18_port, ZN =>
                           n1594);
   U1600 : NAND2_X1 port map( A1 => n3020, A2 => n3019, ZN => n1595);
   U1601 : AOI21_X1 port map( B1 => n1597, B2 => n3017, A => n3049, ZN => n1596
                           );
   U1602 : NAND2_X1 port map( A1 => n1953, A2 => DataP_opcode_W_5_port, ZN => 
                           n3017);
   U1603 : AND2_X1 port map( A1 => n3016, A2 => DataP_opcode_W_3_port, ZN => 
                           n1597);
   U1604 : OAI211_X1 port map( C1 => DataP_opcode_W_4_port, C2 => 
                           DataP_opcode_W_0_port, A => DataP_opcode_W_2_port, B
                           => DataP_opcode_W_1_port, ZN => n3016);
   U1605 : OR2_X4 port map( A1 => n3110, A2 => n3109, ZN => 
                           DataP_alu_a_in_3_port);
   U1606 : OR2_X2 port map( A1 => n3181, A2 => n3180, ZN => 
                           DataP_alu_a_in_14_port);
   U1607 : AND4_X1 port map( A1 => n3262, A2 => n2390, A3 => n3419, A4 => n3263
                           , ZN => n1598);
   U1608 : AND4_X1 port map( A1 => n3262, A2 => n3419, A3 => n2390, A4 => n1896
                           , ZN => n3420);
   U1609 : AOI21_X1 port map( B1 => n3542, B2 => n3691, A => n3541, ZN => n1599
                           );
   U1610 : XNOR2_X1 port map( A => n1959, B => n1600, ZN => n3621);
   U1611 : AND2_X2 port map( A1 => n3611, A2 => n1757, ZN => n1600);
   U1612 : OR2_X1 port map( A1 => n1997, A2 => n2244, ZN => n1601);
   U1613 : OR2_X1 port map( A1 => n1997, A2 => n2244, ZN => n3641);
   U1614 : BUF_X1 port map( A => n1983, Z => n1602);
   U1615 : NOR2_X1 port map( A1 => n1911, A2 => n1965, ZN => n1603);
   U1616 : AOI21_X1 port map( B1 => n3621, B2 => n3691, A => n3620, ZN => n1604
                           );
   U1617 : BUF_X2 port map( A => DataP_alu_a_in_0_port, Z => n1605);
   U1618 : NAND2_X1 port map( A1 => n2425, A2 => n2540, ZN => n1606);
   U1619 : OAI21_X1 port map( B1 => n1957, B2 => n1918, A => n2366, ZN => n1607
                           );
   U1620 : OR2_X2 port map( A1 => n3050, A2 => n1865, ZN => n2472);
   U1621 : AND4_X2 port map( A1 => n1847, A2 => n3028, A3 => n3027, A4 => n3062
                           , ZN => n1861);
   U1622 : NOR2_X1 port map( A1 => DataP_alu_b_in_3_port, A2 => 
                           DataP_alu_b_in_2_port, ZN => n1608);
   U1623 : OR2_X1 port map( A1 => n3692, A2 => n3674, ZN => n1609);
   U1624 : INV_X1 port map( A => n1530, ZN => n1932);
   U1625 : NOR2_X2 port map( A1 => n2555, A2 => n2554, ZN => n2552);
   U1626 : BUF_X1 port map( A => n1552, Z => n1610);
   U1627 : NAND4_X2 port map( A1 => n3334, A2 => n3333, A3 => n3332, A4 => 
                           n3331, ZN => DataP_alu_b_in_21_port);
   U1628 : INV_X1 port map( A => DataP_alu_b_in_6_port, ZN => n1611);
   U1629 : NOR2_X1 port map( A1 => n1911, A2 => n1965, ZN => n2362);
   U1630 : INV_X1 port map( A => n1907, ZN => n1612);
   U1631 : NAND2_X1 port map( A1 => n3677, A2 => n3678, ZN => n3676);
   U1632 : NAND2_X1 port map( A1 => n1613, A2 => n3370, ZN => n3677);
   U1633 : NAND2_X1 port map( A1 => n3372, A2 => n3371, ZN => n1613);
   U1634 : NAND2_X1 port map( A1 => n1561, A2 => n2419, ZN => n3371);
   U1635 : NAND2_X1 port map( A1 => n1816, A2 => n3359, ZN => n3372);
   U1636 : NAND2_X1 port map( A1 => n1619, A2 => n1614, ZN => n3065);
   U1637 : AND2_X1 port map( A1 => n1618, A2 => n1616, ZN => n1614);
   U1638 : NOR2_X1 port map( A1 => n2573, A2 => n2468, ZN => n1615);
   U1639 : NAND2_X1 port map( A1 => n3038, A2 => n3039, ZN => n1620);
   U1640 : OAI211_X1 port map( C1 => n3033, C2 => DataP_opcode_M_4_port, A => 
                           n1622, B => n1621, ZN => n3039);
   U1641 : AOI21_X1 port map( B1 => n1543, B2 => DataP_opcode_M_4_port, A => 
                           DataP_opcode_M_5_port, ZN => n1621);
   U1642 : INV_X1 port map( A => n3032, ZN => n1622);
   U1643 : NAND2_X1 port map( A1 => n1623, A2 => DataP_opcode_M_3_port, ZN => 
                           n3038);
   U1644 : OAI21_X1 port map( B1 => n3036, B2 => n146, A => n3035, ZN => n1623)
                           ;
   U1645 : NOR2_X1 port map( A1 => n1626, A2 => n1625, ZN => n1624);
   U1646 : INV_X1 port map( A => n3103, ZN => n1626);
   U1647 : OAI21_X1 port map( B1 => n150, B2 => DataP_opcode_M_1_port, A => 
                           n1627, ZN => n3032);
   U1648 : NAND2_X1 port map( A1 => DataP_opcode_M_1_port, A2 => 
                           DataP_opcode_M_3_port, ZN => n1627);
   U1649 : INV_X1 port map( A => n2243, ZN => n1632);
   U1650 : OAI211_X1 port map( C1 => n1544, C2 => n1633, A => n1629, B => n1628
                           , ZN => n2418);
   U1651 : NAND3_X1 port map( A1 => n2008, A2 => n2430, A3 => n1632, ZN => 
                           n1628);
   U1652 : INV_X1 port map( A => n1630, ZN => n1629);
   U1653 : OAI21_X1 port map( B1 => n2430, B2 => n1633, A => n1631, ZN => n1630
                           );
   U1654 : NAND2_X2 port map( A1 => n1632, A2 => n2426, ZN => n1631);
   U1655 : NAND2_X2 port map( A1 => n2515, A2 => n2243, ZN => n1633);
   U1656 : NAND2_X1 port map( A1 => n1634, A2 => n1980, ZN => DataP_PC_reg_N31)
                           ;
   U1657 : NAND2_X1 port map( A1 => n2418, A2 => n1982, ZN => n1634);
   U1658 : NAND4_X1 port map( A1 => n3095, A2 => n3093, A3 => n3092, A4 => 
                           n3094, ZN => DataP_alu_b_in_3_port);
   U1659 : BUF_X1 port map( A => n3327, Z => n1635);
   U1660 : INV_X1 port map( A => n2331, ZN => n1636);
   U1661 : AND3_X1 port map( A1 => n3087, A2 => n3090, A3 => n3089, ZN => n1637
                           );
   U1662 : OAI21_X1 port map( B1 => n2380, B2 => n2577, A => n2379, ZN => n1638
                           );
   U1663 : BUF_X1 port map( A => n3565, Z => n1639);
   U1664 : INV_X1 port map( A => n2130, ZN => sra_131_SH_4_port);
   U1665 : AND4_X1 port map( A1 => n3673, A2 => n3681, A3 => n3380, A4 => n3316
                           , ZN => n1856);
   U1666 : OR2_X1 port map( A1 => n3003, A2 => n2233, ZN => n3085);
   U1667 : BUF_X2 port map( A => n1887, Z => n1837);
   U1668 : BUF_X1 port map( A => n3612, Z => n1959);
   U1669 : OR2_X1 port map( A1 => n3512, A2 => n2539, ZN => n2226);
   U1670 : INV_X1 port map( A => n2450, ZN => n1976);
   U1671 : INV_X2 port map( A => n2845, ZN => n2846);
   U1672 : INV_X1 port map( A => n2048, ZN => n1640);
   U1673 : OAI22_X1 port map( A1 => DataP_alu_b_in_31_port, A2 => n1923, B1 => 
                           DataP_alu_a_in_30_port, B2 => n2053, ZN => n1641);
   U1674 : AOI211_X1 port map( C1 => n2055, C2 => n1640, A => n2054, B => n1641
                           , ZN => n2056);
   U1675 : INV_X1 port map( A => lt_x_135_B_4_port, ZN => n1642);
   U1676 : OAI21_X1 port map( B1 => n3671, B2 => n1642, A => n3694, ZN => n1643
                           );
   U1677 : AOI22_X1 port map( A1 => DataP_alu_a_in_4_port, A2 => n1643, B1 => 
                           lt_x_134_B_4_port, B2 => n3697, ZN => n3672);
   U1678 : OAI21_X1 port map( B1 => n2065, B2 => n2984, A => n2980, ZN => n1644
                           );
   U1679 : INV_X1 port map( A => lt_x_134_B_4_port, ZN => n1645);
   U1680 : INV_X1 port map( A => lt_x_135_B_4_port, ZN => n1646);
   U1681 : OAI221_X1 port map( B1 => lt_x_135_B_4_port, B2 => n2837, C1 => 
                           n1646, C2 => n2836, A => n3006, ZN => n1647);
   U1682 : NAND2_X1 port map( A1 => n1645, A2 => n3007, ZN => n1648);
   U1683 : OAI21_X1 port map( B1 => n2708, B2 => n1648, A => n1647, ZN => n1649
                           );
   U1684 : AOI21_X1 port map( B1 => n3659, B2 => n3656, A => n3217, ZN => n1650
                           );
   U1685 : NAND2_X1 port map( A1 => n3232, A2 => n3266, ZN => n1651);
   U1686 : AOI21_X1 port map( B1 => n1650, B2 => n1651, A => n3674, ZN => n1652
                           );
   U1687 : OAI21_X1 port map( B1 => n1650, B2 => n1651, A => n1652, ZN => n1653
                           );
   U1688 : OAI211_X1 port map( C1 => n3700, C2 => n3282, A => n3228, B => n1653
                           , ZN => n1654);
   U1689 : AOI211_X1 port map( C1 => n3675, C2 => n1644, A => n1649, B => n1654
                           , ZN => n341);
   U1690 : NAND4_X1 port map( A1 => n2467, A2 => n1550, A3 => n2503, A4 => 
                           n2133, ZN => n1655);
   U1691 : OAI211_X1 port map( C1 => n2467, C2 => n2133, A => n2367, B => n1655
                           , ZN => n1656);
   U1692 : NAND2_X1 port map( A1 => n1547, A2 => n2321, ZN => n1657);
   U1693 : OAI21_X1 port map( B1 => n2368, B2 => n1656, A => n1657, ZN => n3470
                           );
   U1694 : OAI21_X1 port map( B1 => n2847, B2 => n2983, A => n2977, ZN => n1658
                           );
   U1695 : OAI22_X1 port map( A1 => n3663, A2 => n3664, B1 => n1921, B2 => 
                           n3662, ZN => n1659);
   U1696 : INV_X1 port map( A => lt_x_134_B_4_port, ZN => n1660);
   U1697 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2833, C1 => 
                           n1660, C2 => n2832, A => n3703, ZN => n1661);
   U1698 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2707, ZN => n1662)
                           ;
   U1699 : XNOR2_X1 port map( A => DataP_alu_a_in_8_port, B => n3658, ZN => 
                           n1663);
   U1700 : AOI21_X1 port map( B1 => n3657, B2 => n3656, A => n3659, ZN => n1664
                           );
   U1701 : AOI211_X1 port map( C1 => n3659, C2 => n1663, A => n1664, B => n3674
                           , ZN => n1665);
   U1702 : AOI21_X1 port map( B1 => n3706, B2 => n1662, A => n1665, ZN => n1666
                           );
   U1703 : NAND2_X1 port map( A1 => n1661, A2 => n1666, ZN => n1667);
   U1704 : AOI211_X1 port map( C1 => n3675, C2 => n1658, A => n1659, B => n1667
                           , ZN => n345);
   U1705 : NAND3_X1 port map( A1 => n3488, A2 => n3509, A3 => n1917, ZN => 
                           n1668);
   U1706 : XOR2_X1 port map( A => DataP_alu_b_in_29_port, B => n1668, Z => 
                           n2371);
   U1707 : NAND2_X1 port map( A1 => n2565, A2 => DataP_IMM_s_18_port, ZN => 
                           n1669);
   U1708 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_14_port, ZN => 
                           n1670);
   U1709 : NAND3_X1 port map( A1 => n1670, A2 => n3312, A3 => n3311, ZN => 
                           n1671);
   U1710 : AOI21_X1 port map( B1 => n3001, B2 => DataP_B_s_14_port, A => n1671,
                           ZN => n3418);
   U1711 : XOR2_X1 port map( A => n3665, B => n1851, Z => n1672);
   U1712 : AOI22_X1 port map( A1 => n1915, A2 => n2823, B1 => n2064, B2 => 
                           n2822, ZN => n1673);
   U1713 : INV_X1 port map( A => lt_x_135_B_4_port, ZN => n1674);
   U1714 : OAI221_X1 port map( B1 => lt_x_135_B_4_port, B2 => n1673, C1 => 
                           n1674, C2 => n2824, A => n3703, ZN => n1675);
   U1715 : INV_X1 port map( A => n2968, ZN => n1676);
   U1716 : INV_X1 port map( A => n2065, ZN => n1677);
   U1717 : OAI221_X1 port map( B1 => n2065, B2 => n1676, C1 => n1677, C2 => 
                           n2967, A => n3675, ZN => n1678);
   U1718 : OAI211_X1 port map( C1 => n1672, C2 => n3674, A => n1675, B => n1678
                           , ZN => n1679);
   U1719 : AOI21_X1 port map( B1 => n3667, B2 => n3694, A => n2363, ZN => n1680
                           );
   U1720 : AOI21_X1 port map( B1 => n3697, B2 => DataP_alu_a_in_6_port, A => 
                           n1680, ZN => n1681);
   U1721 : NAND3_X1 port map( A1 => n3007, A2 => n2693, A3 => n1674, ZN => 
                           n1682);
   U1722 : OAI211_X1 port map( C1 => n3700, C2 => n3668, A => n1681, B => n1682
                           , ZN => n1683);
   U1723 : NOR2_X1 port map( A1 => n1679, A2 => n1683, ZN => n353);
   U1724 : AOI22_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_26_port, B1 =>
                           n3001, B2 => DataP_B_s_26_port, ZN => n1684);
   U1725 : OAI211_X1 port map( C1 => n1636, C2 => n2169, A => n3306, B => n1684
                           , ZN => DataP_alu_b_in_26_port);
   U1726 : AOI22_X1 port map( A1 => DataP_alu_a_in_5_port, A2 => n3379, B1 => 
                           lt_x_134_B_5_port, B2 => n3697, ZN => n1685);
   U1727 : INV_X1 port map( A => lt_x_134_B_4_port, ZN => n1686);
   U1728 : NAND3_X1 port map( A1 => n3007, A2 => n2692, A3 => n1686, ZN => 
                           n1687);
   U1729 : OAI211_X1 port map( C1 => n3380, C2 => n3700, A => n1685, B => n1687
                           , ZN => n1688);
   U1730 : NAND2_X1 port map( A1 => n1899, A2 => n3382, ZN => n1689);
   U1731 : XNOR2_X1 port map( A => n1689, B => n3383, ZN => n1690);
   U1732 : AOI22_X1 port map( A1 => n2064, A2 => n2817, B1 => n1915, B2 => 
                           n2818, ZN => n1691);
   U1733 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n1691, C1 => 
                           n1686, C2 => n2819, A => n3006, ZN => n1692);
   U1734 : OAI21_X1 port map( B1 => n2065, B2 => n2963, A => n2962, ZN => n1693
                           );
   U1735 : NAND2_X1 port map( A1 => n1693, A2 => n3675, ZN => n1694);
   U1736 : OAI211_X1 port map( C1 => n3674, C2 => n1690, A => n1692, B => n1694
                           , ZN => n1695);
   U1737 : NOR2_X1 port map( A1 => n1688, A2 => n1695, ZN => n354);
   U1738 : INV_X1 port map( A => n3392, ZN => n1696);
   U1739 : NAND3_X1 port map( A1 => n3510, A2 => n1841, A3 => n1696, ZN => 
                           n3416);
   U1740 : AOI22_X1 port map( A1 => n2846, A2 => n2635, B1 => n2127, B2 => 
                           n2687, ZN => n1697);
   U1741 : INV_X1 port map( A => lt_x_135_B_4_port, ZN => n1698);
   U1742 : OAI221_X1 port map( B1 => lt_x_135_B_4_port, B2 => n1697, C1 => 
                           n1698, C2 => n2694, A => n3706, ZN => n3451);
   U1743 : AND3_X2 port map( A1 => n2245, A2 => n2306, A3 => n1522, ZN => n2136
                           );
   U1744 : AOI21_X1 port map( B1 => n2301, B2 => n2300, A => n2183, ZN => n1699
                           );
   U1745 : OAI211_X1 port map( C1 => n1946, C2 => DataP_alu_b_in_18_port, A => 
                           n3426, B => n2496, ZN => n1700);
   U1746 : NAND2_X1 port map( A1 => n1932, A2 => n2478, ZN => n1701);
   U1747 : NAND2_X1 port map( A1 => n3510, A2 => n2377, ZN => n1702);
   U1748 : NAND2_X1 port map( A1 => n3400, A2 => n2372, ZN => n1703);
   U1749 : OAI211_X1 port map( C1 => n1702, C2 => n3400, A => n1703, B => n1701
                           , ZN => n3401);
   U1750 : AOI22_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_30_port, B1 =>
                           DataP_B_s_30_port, B2 => n1859, ZN => n1704);
   U1751 : OAI211_X1 port map( C1 => n2566, C2 => n2187, A => n3306, B => n1704
                           , ZN => DataP_alu_b_in_30_port);
   U1752 : NOR2_X1 port map( A1 => lt_x_134_B_4_port, A2 => n2705, ZN => n1705)
                           ;
   U1753 : XNOR2_X1 port map( A => DataP_alu_a_in_4_port, B => n3670, ZN => 
                           n1706);
   U1754 : XNOR2_X1 port map( A => n1706, B => n1961, ZN => n1707);
   U1755 : OAI21_X1 port map( B1 => n2847, B2 => n2956, A => n2955, ZN => n1708
                           );
   U1756 : NAND2_X1 port map( A1 => n1708, A2 => n3675, ZN => n1709);
   U1757 : OAI21_X1 port map( B1 => n3674, B2 => n1707, A => n1709, ZN => n1710
                           );
   U1758 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2814, C1 => 
                           n1645, C2 => n2813, A => n3703, ZN => n1711);
   U1759 : OAI211_X1 port map( C1 => n3673, C2 => n3700, A => n3672, B => n1711
                           , ZN => n1712);
   U1760 : AOI211_X1 port map( C1 => n3007, C2 => n1705, A => n1710, B => n1712
                           , ZN => n355);
   U1761 : AOI21_X1 port map( B1 => n2478, B2 => n2407, A => 
                           DataP_alu_a_in_29_port, ZN => n2279);
   U1762 : XNOR2_X1 port map( A => DataP_alu_a_in_8_port, B => n3663, ZN => 
                           n1713);
   U1763 : AOI211_X1 port map( C1 => n3335, C2 => n3317, A => n3402, B => n1713
                           , ZN => n1714);
   U1764 : AND3_X1 port map( A1 => n2452, A2 => n1714, A3 => n3668, ZN => n1853
                           );
   U1765 : OAI21_X1 port map( B1 => n2573, B2 => n151, A => 
                           DataP_opcode_E_4_port, ZN => n1715);
   U1766 : AND2_X1 port map( A1 => DataP_opcode_E_3_port, A2 => n2573, ZN => 
                           n1716);
   U1767 : OAI33_X1 port map( A1 => n1715, A2 => n2575, A3 => n1716, B1 => 
                           DataP_opcode_E_4_port, B2 => DataP_opcode_E_0_port, 
                           B3 => n149, ZN => n1717);
   U1768 : AOI21_X1 port map( B1 => n3060, B2 => DataP_opcode_E_4_port, A => 
                           n145, ZN => n1718);
   U1769 : OAI21_X1 port map( B1 => n521, B2 => n520, A => 
                           DataP_opcode_E_3_port, ZN => n1719);
   U1770 : NOR2_X1 port map( A1 => n1718, A2 => n1719, ZN => n1720);
   U1771 : AOI21_X1 port map( B1 => n145, B2 => n1717, A => n1720, ZN => n3073)
                           ;
   U1772 : AOI22_X1 port map( A1 => n3001, A2 => DataP_B_s_25_port, B1 => n3005
                           , B2 => DataP_alu_out_W_25_port, ZN => n1721);
   U1773 : NAND4_X1 port map( A1 => n1882, A2 => n3458, A3 => n2526, A4 => 
                           n2540, ZN => n2424);
   U1774 : AOI22_X1 port map( A1 => n2843, A2 => n2826, B1 => n2844, B2 => 
                           n2825, ZN => n1722);
   U1775 : AOI22_X1 port map( A1 => n1915, A2 => n2827, B1 => n2845, B2 => 
                           n1722, ZN => n2829);
   U1776 : NOR2_X1 port map( A1 => n3510, A2 => n2279, ZN => n1723);
   U1777 : NAND2_X1 port map( A1 => n2281, A2 => n2279, ZN => n1724);
   U1778 : OAI211_X1 port map( C1 => n2371, C2 => n1723, A => n2280, B => n1724
                           , ZN => n2513);
   U1779 : NOR2_X1 port map( A1 => n2177, A2 => n2566, ZN => n1725);
   U1780 : AOI21_X1 port map( B1 => n1515, B2 => DataP_ir_E_12_port, A => n1725
                           , ZN => n1726);
   U1781 : NAND3_X1 port map( A1 => n1726, A2 => n3261, A3 => n2387, ZN => 
                           DataP_alu_b_in_12_port);
   U1782 : NOR2_X1 port map( A1 => n3249, A2 => n1879, ZN => n1727);
   U1783 : XNOR2_X1 port map( A => n1727, B => n1572, ZN => n3251);
   U1784 : OAI221_X1 port map( B1 => n2122, B2 => n2120, C1 => n2122, C2 => 
                           n2121, A => n2119, ZN => n1728);
   U1785 : MUX2_X1 port map( A => n1983, B => n1728, S => ALU_OPCODE_i_2_port, 
                           Z => n3346);
   U1786 : NOR2_X1 port map( A1 => n2713, A2 => n2578, ZN => n1729);
   U1787 : AOI22_X1 port map( A1 => n2599, A2 => n1930, B1 => n2842, B2 => 
                           n1729, ZN => n2622);
   U1788 : AOI22_X1 port map( A1 => n3423, A2 => n1520, B1 => n2002, B2 => 
                           n1840, ZN => n1730);
   U1789 : OAI21_X1 port map( B1 => n1591, B2 => n1730, A => n1960, ZN => n3428
                           );
   U1790 : OAI21_X1 port map( B1 => DataP_alu_a_in_25_port, B2 => n1547, A => 
                           n3697, ZN => n1731);
   U1791 : NAND3_X1 port map( A1 => DataP_alu_a_in_25_port, A2 => n1547, A3 => 
                           n3693, ZN => n1732);
   U1792 : OAI211_X1 port map( C1 => n3547, C2 => n3700, A => n1731, B => n1732
                           , ZN => n3548);
   U1793 : AOI22_X1 port map( A1 => n2508, A2 => n2003, B1 => n3689, B2 => 
                           n3663, ZN => n1733);
   U1794 : NAND3_X1 port map( A1 => n2509, A2 => n2507, A3 => n1733, ZN => 
                           n3658);
   U1795 : OAI21_X1 port map( B1 => n2065, B2 => n2949, A => n2948, ZN => n1734
                           );
   U1796 : AOI22_X1 port map( A1 => n1916, A2 => n2805, B1 => n2840, B2 => 
                           n2806, ZN => n1735);
   U1797 : AOI22_X1 port map( A1 => n2842, A2 => n2825, B1 => n1930, B2 => 
                           n1735, ZN => n1736);
   U1798 : AOI22_X1 port map( A1 => n2330, A2 => n1736, B1 => n2846, B2 => 
                           n2807, ZN => n1737);
   U1799 : INV_X1 port map( A => lt_x_135_B_4_port, ZN => n1738);
   U1800 : OAI221_X1 port map( B1 => lt_x_135_B_4_port, B2 => n1737, C1 => 
                           n1738, C2 => n2808, A => n3006, ZN => n1739);
   U1801 : INV_X1 port map( A => n2690, ZN => n1740);
   U1802 : AOI22_X1 port map( A1 => DataP_alu_a_in_3_port, A2 => n3680, B1 => 
                           n1963, B2 => n3697, ZN => n1741);
   U1803 : OAI211_X1 port map( C1 => n3678, C2 => n1993, A => n2001, B => n3691
                           , ZN => n1742);
   U1804 : OAI211_X1 port map( C1 => n3700, C2 => n3681, A => n1741, B => n1742
                           , ZN => n1743);
   U1805 : NOR2_X1 port map( A1 => n1740, A2 => lt_x_134_B_4_port, ZN => n1744)
                           ;
   U1806 : AOI21_X1 port map( B1 => n1744, B2 => n3706, A => n1743, ZN => n1745
                           );
   U1807 : NAND2_X1 port map( A1 => n1745, A2 => n1739, ZN => n1746);
   U1808 : AOI21_X1 port map( B1 => n3675, B2 => n1734, A => n1746, ZN => n356)
                           ;
   U1809 : OAI21_X1 port map( B1 => n1589, B2 => DataP_alu_b_in_21_port, A => 
                           DataP_alu_b_in_20_port, ZN => n1747);
   U1810 : OAI22_X1 port map( A1 => DataP_alu_a_in_20_port, A2 => n1747, B1 => 
                           DataP_alu_a_in_21_port, B2 => n1952, ZN => n2107);
   U1811 : INV_X1 port map( A => n1838, ZN => n1748);
   U1812 : NAND2_X1 port map( A1 => n2493, A2 => n3510, ZN => n1749);
   U1813 : AOI21_X1 port map( B1 => n2538, B2 => n1749, A => n1748, ZN => n2491
                           );
   U1814 : NAND2_X1 port map( A1 => n1947, A2 => n1881, ZN => n1750);
   U1815 : NAND2_X1 port map( A1 => n1932, A2 => n1750, ZN => n2377);
   U1816 : INV_X1 port map( A => n1605, ZN => n1751);
   U1817 : NAND2_X1 port map( A1 => n2985, A2 => n1751, ZN => n3335);
   U1818 : AND4_X1 port map( A1 => n2476, A2 => n3058, A3 => n2477, A4 => n2163
                           , ZN => n1752);
   U1819 : NAND4_X1 port map( A1 => n3062, A2 => n3064, A3 => n1752, A4 => 
                           n1883, ZN => n3069);
   U1820 : AOI22_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_29_port, B1 =>
                           n1859, B2 => DataP_B_s_29_port, ZN => n1753);
   U1821 : NAND2_X1 port map( A1 => n2331, A2 => DataP_alu_out_M_29_port, ZN =>
                           n1754);
   U1822 : NAND3_X1 port map( A1 => n1754, A2 => n1753, A3 => n3306, ZN => 
                           DataP_alu_b_in_29_port);
   U1823 : NAND3_X1 port map( A1 => n3510, A2 => DataP_alu_a_in_11_port, A3 => 
                           n3251, ZN => n3272);
   U1824 : INV_X1 port map( A => n3202, ZN => n1755);
   U1825 : NAND2_X1 port map( A1 => DataP_alu_a_in_3_port, A2 => n1755, ZN => 
                           n3375);
   U1826 : OAI21_X1 port map( B1 => DataP_alu_b_in_22_port, B2 => n3510, A => 
                           DataP_alu_a_in_22_port, ZN => n1756);
   U1827 : AOI21_X1 port map( B1 => n3446, B2 => n3510, A => n1756, ZN => n2312
                           );
   U1828 : NAND2_X1 port map( A1 => n1986, A2 => n1878, ZN => n1757);
   U1829 : OAI22_X1 port map( A1 => n2989, A2 => n3694, B1 => n1561, B2 => 
                           n3373, ZN => n1758);
   U1830 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2704, ZN => n1759)
                           ;
   U1831 : NAND2_X1 port map( A1 => n3370, A2 => n3371, ZN => n1760);
   U1832 : XNOR2_X1 port map( A => n1760, B => n3372, ZN => n1761);
   U1833 : AOI22_X1 port map( A1 => n1759, A2 => n3706, B1 => n1761, B2 => 
                           n3691, ZN => n1762);
   U1834 : INV_X1 port map( A => n2937, ZN => n1763);
   U1835 : INV_X1 port map( A => n2065, ZN => n1764);
   U1836 : AOI22_X1 port map( A1 => n2841, A2 => n2964, B1 => n2935, B2 => 
                           n2989, ZN => n1765);
   U1837 : AOI22_X1 port map( A1 => n2846, A2 => n2936, B1 => n2845, B2 => 
                           n1765, ZN => n1766);
   U1838 : OAI221_X1 port map( B1 => n2065, B2 => n1763, C1 => n1764, C2 => 
                           n1766, A => n3675, ZN => n1767);
   U1839 : AOI22_X1 port map( A1 => n2846, A2 => n2799, B1 => n2845, B2 => 
                           n2798, ZN => n1768);
   U1840 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n1768, C1 => 
                           n1660, C2 => n2800, A => n3703, ZN => n1769);
   U1841 : NAND3_X1 port map( A1 => n1762, A2 => n1767, A3 => n1769, ZN => 
                           n1770);
   U1842 : AOI211_X1 port map( C1 => n3374, C2 => n1939, A => n1758, B => n1770
                           , ZN => n357);
   U1843 : XNOR2_X1 port map( A => n1946, B => DataP_alu_b_in_18_port, ZN => 
                           n2300);
   U1844 : AOI22_X1 port map( A1 => n2997, A2 => DataP_alu_out_M_17_port, B1 =>
                           DataP_alu_out_W_17_port, B2 => n2992, ZN => n1771);
   U1845 : OAI21_X1 port map( B1 => n57, B2 => n2999, A => n1771, ZN => n3172);
   U1846 : INV_X1 port map( A => n2109, ZN => n1772);
   U1847 : AOI221_X1 port map( B1 => n2123, B2 => n2117, C1 => n2116, C2 => 
                           n2117, A => n2124, ZN => n1773);
   U1848 : OAI22_X1 port map( A1 => DataP_alu_a_in_31_port, A2 => n1935, B1 => 
                           DataP_alu_a_in_30_port, B2 => n2118, ZN => n1774);
   U1849 : INV_X1 port map( A => n3490, ZN => n1775);
   U1850 : NAND2_X1 port map( A1 => n3510, A2 => n1775, ZN => n1776);
   U1851 : XNOR2_X1 port map( A => n1917, B => n1776, ZN => n3523);
   U1852 : OAI221_X1 port map( B1 => n3510, B2 => n2358, C1 => n2383, C2 => 
                           n3233, A => n3236, ZN => n3268);
   U1853 : AOI21_X1 port map( B1 => n2383, B2 => n2382, A => 
                           DataP_alu_a_in_21_port, ZN => n2379);
   U1854 : AOI21_X1 port map( B1 => n3465, B2 => n2131, A => n2421, ZN => n1777
                           );
   U1855 : NAND2_X1 port map( A1 => n2422, A2 => n1777, ZN => n3533);
   U1856 : AOI211_X1 port map( C1 => n3353, C2 => n3352, A => n2132, B => 
                           ALU_OPCODE_i_0_port, ZN => n1778);
   U1857 : AOI211_X1 port map( C1 => n3353, C2 => DataP_ALU_C_comp_N24, A => 
                           ALU_OPCODE_i_1_port, B => n2150, ZN => n1779);
   U1858 : OR2_X1 port map( A1 => n1778, A2 => n1779, ZN => n3354);
   U1859 : OAI221_X1 port map( B1 => n1520, B2 => n3456, C1 => n1520, C2 => 
                           n2002, A => n3423, ZN => n1987);
   U1860 : AND4_X1 port map( A1 => n2477, A2 => n2476, A3 => n3058, A4 => n2163
                           , ZN => n1780);
   U1861 : AND3_X1 port map( A1 => n3062, A2 => Rst, A3 => n1780, ZN => n2475);
   U1862 : INV_X1 port map( A => n1899, ZN => n1781);
   U1863 : AOI21_X1 port map( B1 => n3382, B2 => n3383, A => n1781, ZN => n3665
                           );
   U1864 : NOR2_X1 port map( A1 => DataP_alu_b_in_19_port, A2 => n1938, ZN => 
                           n2496);
   U1865 : NAND2_X1 port map( A1 => DataP_alu_a_in_26_port, A2 => n1936, ZN => 
                           n1782);
   U1866 : OAI21_X1 port map( B1 => n1912, B2 => DataP_alu_b_in_27_port, A => 
                           n1782, ZN => n2060);
   U1867 : AOI21_X1 port map( B1 => n2478, B2 => n2512, A => 
                           DataP_alu_a_in_16_port, ZN => n1979);
   U1868 : NOR2_X1 port map( A1 => n3554, A2 => n2556, ZN => n2131);
   U1869 : AOI22_X1 port map( A1 => n3001, A2 => DataP_B_s_23_port, B1 => n2565
                           , B2 => DataP_IMM_s_23_port, ZN => n1783);
   U1870 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_23_port, ZN =>
                           n1784);
   U1871 : OAI211_X1 port map( C1 => n1636, C2 => n2168, A => n1783, B => n1784
                           , ZN => DataP_alu_b_in_23_port);
   U1872 : AOI22_X1 port map( A1 => n2846, A2 => n2648, B1 => n2127, B2 => 
                           n2647, ZN => n1785);
   U1873 : INV_X1 port map( A => lt_x_135_B_4_port, ZN => n1786);
   U1874 : OAI221_X1 port map( B1 => lt_x_135_B_4_port, B2 => n1785, C1 => 
                           n1786, C2 => n2618, A => n3007, ZN => n3617);
   U1875 : AOI22_X1 port map( A1 => n2842, A2 => n2652, B1 => n1913, B2 => 
                           n2677, ZN => n1787);
   U1876 : AOI22_X1 port map( A1 => n2127, A2 => n1787, B1 => n2653, B2 => 
                           n1915, ZN => n1788);
   U1877 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n1788, C1 => 
                           n1686, C2 => n2654, A => n3007, ZN => n3540);
   U1878 : OAI211_X1 port map( C1 => n2321, C2 => n2365, A => n2364, B => n1944
                           , ZN => n3580);
   U1879 : INV_X1 port map( A => n1960, ZN => n1789);
   U1880 : NOR2_X1 port map( A1 => n1591, A2 => n1789, ZN => n2572);
   U1881 : NAND3_X1 port map( A1 => DataP_alu_a_in_14_port, A2 => n1932, A3 => 
                           n3693, ZN => n1790);
   U1882 : OAI21_X1 port map( B1 => DataP_alu_a_in_14_port, B2 => n1932, A => 
                           n3697, ZN => n1791);
   U1883 : OAI211_X1 port map( C1 => n3633, C2 => n3700, A => n1790, B => n1791
                           , ZN => n3634);
   U1884 : NAND2_X1 port map( A1 => n3657, A2 => n3266, ZN => n1792);
   U1885 : INV_X1 port map( A => n3659, ZN => n1793);
   U1886 : NAND2_X1 port map( A1 => n3232, A2 => n1792, ZN => n1794);
   U1887 : OAI21_X1 port map( B1 => n1793, B2 => n3267, A => n1794, ZN => n3248
                           );
   U1888 : AOI22_X1 port map( A1 => n2127, A2 => n2978, B1 => n1915, B2 => 
                           n2979, ZN => n1795);
   U1889 : NAND2_X1 port map( A1 => n2065, A2 => n1795, ZN => n2980);
   U1890 : AOI22_X1 port map( A1 => n2064, A2 => n2975, B1 => n1915, B2 => 
                           n2976, ZN => n1796);
   U1891 : NAND2_X1 port map( A1 => n2065, A2 => n1796, ZN => n2977);
   U1892 : AOI22_X1 port map( A1 => n1914, A2 => DataP_alu_a_in_2_port, B1 => 
                           n1931, B2 => DataP_alu_a_in_1_port, ZN => n1797);
   U1893 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2805, B1 => n1916
                           , B2 => n1797, ZN => n2772);
   U1894 : AOI21_X1 port map( B1 => n3050, B2 => n3049, A => n1865, ZN => n1798
                           );
   U1895 : INV_X1 port map( A => n1798, ZN => n3064);
   U1896 : INV_X1 port map( A => n3983, ZN => n1799);
   U1897 : AOI221_X1 port map( B1 => n3984, B2 => n3983, C1 => n3709, C2 => 
                           n1799, A => n3982, ZN => DataP_wrong_br);
   U1898 : NOR2_X1 port map( A1 => lt_x_134_B_4_port, A2 => n2706, ZN => n1800)
                           ;
   U1899 : OAI21_X1 port map( B1 => n3665, B2 => n3386, A => n3385, ZN => n1801
                           );
   U1900 : XOR2_X1 port map( A => DataP_alu_a_in_7_port, B => n3213, Z => n1802
                           );
   U1901 : XNOR2_X1 port map( A => n1801, B => n1802, ZN => n1803);
   U1902 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N89, A2 => n3675, ZN =>
                           n1804);
   U1903 : OAI21_X1 port map( B1 => n3674, B2 => n1803, A => n1804, ZN => n1805
                           );
   U1904 : INV_X1 port map( A => lt_x_134_B_4_port, ZN => n1806);
   U1905 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2829, C1 => 
                           n1806, C2 => n2828, A => n3006, ZN => n1807);
   U1906 : OAI211_X1 port map( C1 => n3700, C2 => n3390, A => n3389, B => n1807
                           , ZN => n1808);
   U1907 : AOI211_X1 port map( C1 => n3007, C2 => n1800, A => n1805, B => n1808
                           , ZN => n350);
   U1908 : AOI22_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_31_port, B1 =>
                           DataP_B_s_31_port, B2 => n1859, ZN => n1809);
   U1909 : AOI221_X1 port map( B1 => n3709, B2 => n3983, C1 => n3984, C2 => 
                           n1799, A => n3982, ZN => DataP_right_br);
   U1910 : AOI221_X1 port map( B1 => n2061, B2 => n2103, C1 => n2102, C2 => 
                           n2103, A => n2046, ZN => n1810);
   U1911 : INV_X1 port map( A => DataP_alu_a_in_28_port, ZN => n1811);
   U1912 : NAND2_X1 port map( A1 => n3523, A2 => n1811, ZN => n2515);
   U1913 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_10_port, ZN =>
                           n2388);
   U1914 : OR2_X1 port map( A1 => sra_131_SH_4_port, A2 => n3510, ZN => n2461);
   U1915 : INV_X1 port map( A => n3470, ZN => n1812);
   U1916 : NAND2_X1 port map( A1 => n1929, A2 => n1812, ZN => n3543);
   U1917 : INV_X1 port map( A => n3493, ZN => n1813);
   U1918 : NAND2_X1 port map( A1 => DataP_alu_a_in_30_port, A2 => n1813, ZN => 
                           n3683);
   U1919 : OR2_X1 port map( A1 => n3401, A2 => DataP_alu_a_in_14_port, ZN => 
                           n3410);
   U1920 : AOI21_X1 port map( B1 => n2543, B2 => n2547, A => 
                           DataP_alu_a_in_12_port, ZN => n2542);
   U1921 : NAND2_X1 port map( A1 => n3203, A2 => n3011, ZN => n1814);
   U1922 : NAND2_X1 port map( A1 => n1814, A2 => n3510, ZN => n1815);
   U1923 : XNOR2_X1 port map( A => n1815, B => n2330, ZN => n3202);
   U1924 : NAND2_X1 port map( A1 => n3358, A2 => n3361, ZN => n1816);
   U1925 : NAND3_X1 port map( A1 => n3007, A2 => n2602, A3 => n1806, ZN => 
                           n3339);
   U1926 : OAI221_X1 port map( B1 => n2981, B2 => n2924, C1 => n2981, C2 => 
                           n2065, A => n3675, ZN => n3538);
   U1927 : AOI21_X1 port map( B1 => n3466, B2 => n3467, A => n3465, ZN => n1817
                           );
   U1928 : INV_X1 port map( A => n1817, ZN => n2423);
   U1929 : AOI22_X1 port map( A1 => n2127, A2 => n2670, B1 => n2846, B2 => 
                           n2626, ZN => n1818);
   U1930 : MUX2_X1 port map( A => n1818, B => n2692, S => lt_x_135_B_4_port, Z 
                           => DataP_ALU_C_shifter_N39);
   U1931 : AOI22_X1 port map( A1 => n2064, A2 => n2653, B1 => n2846, B2 => 
                           n2611, ZN => n1819);
   U1932 : MUX2_X1 port map( A => n1819, B => n2673, S => lt_x_134_B_4_port, Z 
                           => DataP_ALU_C_shifter_N36);
   U1933 : INV_X1 port map( A => n3658, ZN => n1820);
   U1934 : NAND2_X1 port map( A1 => DataP_alu_a_in_8_port, A2 => n1820, ZN => 
                           n3657);
   U1935 : AOI22_X1 port map( A1 => n2841, A2 => n2965, B1 => n2989, B2 => 
                           n2964, ZN => n1821);
   U1936 : AOI22_X1 port map( A1 => n1915, A2 => n2966, B1 => n2845, B2 => 
                           n1821, ZN => n2967);
   U1937 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_2_port, B1 => 
                           n2710, B2 => DataP_alu_a_in_1_port, ZN => n1822);
   U1938 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2942, B1 => n2988
                           , B2 => n1822, ZN => n2905);
   U1939 : NOR3_X1 port map( A1 => n3806, A2 => IR_CU_4_port, A3 => 
                           IR_CU_5_port, ZN => n1823);
   U1940 : AOI21_X1 port map( B1 => n3797, B2 => n606, A => n1823, ZN => n1824)
                           ;
   U1941 : OAI221_X1 port map( B1 => n3837, B2 => n3828, C1 => n3837, C2 => 
                           n3817, A => n1824, ZN => n3807);
   U1942 : AOI22_X1 port map( A1 => n2842, A2 => n2656, B1 => n1913, B2 => 
                           n2685, ZN => n1825);
   U1943 : AOI22_X1 port map( A1 => n2127, A2 => n1825, B1 => n2657, B2 => 
                           n1915, ZN => n1826);
   U1944 : OAI221_X1 port map( B1 => lt_x_134_B_4_port, B2 => n1826, C1 => 
                           n1806, C2 => n2658, A => n3007, ZN => n3480);
   U1945 : AND3_X1 port map( A1 => n2475, A2 => n3070, A3 => n3064, ZN => n3710
                           );
   U1946 : NAND2_X1 port map( A1 => n3765, A2 => n3766, ZN => n1827);
   U1947 : NOR3_X1 port map( A1 => n3770, A2 => n3771, A3 => n3772, ZN => n1828
                           );
   U1948 : NAND4_X1 port map( A1 => n3773, A2 => n3774, A3 => n3769, A4 => 
                           n1828, ZN => n1829);
   U1949 : NOR4_X1 port map( A1 => n3767, A2 => n3768, A3 => n1827, A4 => n1829
                           , ZN => n1830);
   U1950 : INV_X1 port map( A => n3757, ZN => n1831);
   U1951 : NAND4_X1 port map( A1 => n3758, A2 => n3759, A3 => n3760, A4 => 
                           n1831, ZN => n1832);
   U1952 : NOR2_X1 port map( A1 => n3755, A2 => n3756, ZN => n1833);
   U1953 : NAND3_X1 port map( A1 => n3754, A2 => n3753, A3 => n1833, ZN => 
                           n1834);
   U1954 : NOR4_X1 port map( A1 => n3761, A2 => n3762, A3 => n1832, A4 => n1834
                           , ZN => n1835);
   U1955 : NAND4_X1 port map( A1 => n3763, A2 => n3764, A3 => n1830, A4 => 
                           n1835, ZN => n1836);
   U1956 : NAND2_X1 port map( A1 => n3775, A2 => n1836, ZN => DataP_NPC_add_N0)
                           ;
   U1957 : CLKBUF_X3 port map( A => n1907, Z => n2988);
   U1958 : NAND4_X1 port map( A1 => n2388, A2 => n3231, A3 => n3230, A4 => 
                           n2335, ZN => n1879);
   U1959 : NOR2_X1 port map( A1 => n3172, A2 => n3171, ZN => n1838);
   U1960 : OR2_X2 port map( A1 => n3131, A2 => n3130, ZN => 
                           DataP_alu_a_in_31_port);
   U1961 : AND2_X1 port map( A1 => n3456, A2 => n3423, ZN => n1840);
   U1962 : BUF_X2 port map( A => n3193, Z => n2999);
   U1963 : INV_X1 port map( A => n1864, ZN => n1841);
   U1964 : INV_X1 port map( A => DataP_alu_a_in_15_port, ZN => n1842);
   U1965 : INV_X1 port map( A => n1864, ZN => DataP_alu_a_in_15_port);
   U1966 : NOR2_X1 port map( A1 => n3178, A2 => n3177, ZN => n1864);
   U1967 : AND4_X1 port map( A1 => n3103, A2 => n3102, A3 => n3101, A4 => n3100
                           , ZN => n1843);
   U1968 : BUF_X4 port map( A => sra_131_SH_4_port, Z => lt_x_134_B_4_port);
   U1969 : NAND2_X1 port map( A1 => n2469, A2 => n2470, ZN => n1844);
   U1970 : NAND2_X1 port map( A1 => n2469, A2 => n2470, ZN => n1845);
   U1971 : NAND2_X1 port map( A1 => n2469, A2 => n2470, ZN => n2998);
   U1972 : OR2_X4 port map( A1 => n3119, A2 => n3118, ZN => 
                           DataP_alu_a_in_4_port);
   U1973 : AND2_X1 port map( A1 => n1518, A2 => DataP_B_s_9_port, ZN => n1846);
   U1974 : NAND4_X1 port map( A1 => n1588, A2 => n2186, A3 => n3023, A4 => 
                           n2140, ZN => n1847);
   U1975 : BUF_X1 port map( A => n3328, Z => n1848);
   U1976 : BUF_X1 port map( A => n3328, Z => n2565);
   U1977 : BUF_X1 port map( A => n3328, Z => n1905);
   U1978 : AOI21_X2 port map( B1 => n3412, B2 => n3411, A => n2541, ZN => n2540
                           );
   U1979 : NAND3_X1 port map( A1 => n1967, A2 => n3494, A3 => n3497, ZN => 
                           n1849);
   U1980 : NAND3_X1 port map( A1 => n3501, A2 => n3499, A3 => n3500, ZN => 
                           n1850);
   U1981 : BUF_X1 port map( A => n3666, Z => n1851);
   U1982 : INV_X1 port map( A => n1862, ZN => n1852);
   U1983 : AND4_X2 port map( A1 => n1853, A2 => n1854, A3 => n1855, A4 => n1856
                           , ZN => n2369);
   U1984 : AND3_X1 port map( A1 => n3484, A2 => n3701, A3 => n3633, ZN => n1854
                           );
   U1985 : AND4_X1 port map( A1 => n3615, A2 => n3624, A3 => n3651, A4 => n3390
                           , ZN => n1855);
   U1986 : AND2_X1 port map( A1 => n3067, A2 => n3066, ZN => n1857);
   U1987 : INV_X1 port map( A => n3001, ZN => n1858);
   U1988 : INV_X1 port map( A => n1858, ZN => n1859);
   U1989 : INV_X1 port map( A => n3396, ZN => n1860);
   U1990 : AND3_X1 port map( A1 => n2442, A2 => n1994, A3 => n2010, ZN => n1889
                           );
   U1991 : INV_X1 port map( A => n1565, ZN => n3330);
   U1992 : BUF_X1 port map( A => n536, Z => n1862);
   U1993 : NOR2_X2 port map( A1 => n3190, A2 => n3189, ZN => n1863);
   U1994 : AND3_X1 port map( A1 => n3016, A2 => n3017, A3 => 
                           DataP_opcode_W_3_port, ZN => n1865);
   U1995 : AND2_X1 port map( A1 => n2322, A2 => n2320, ZN => n1866);
   U1996 : XOR2_X1 port map( A => n2570, B => DataP_add_D_3_port, Z => n2186);
   U1997 : BUF_X1 port map( A => n1548, Z => n1867);
   U1998 : OR2_X1 port map( A1 => n1567, A2 => n117, ZN => n1868);
   U1999 : INV_X1 port map( A => DataP_dest_M_0_port, ZN => n1869);
   U2000 : XNOR2_X1 port map( A => n2576, B => n1894, ZN => n3036);
   U2001 : XNOR2_X1 port map( A => n1870, B => n1933, ZN => n3446);
   U2002 : NOR2_X1 port map( A1 => n3444, A2 => n3445, ZN => n1870);
   U2003 : BUF_X1 port map( A => n538, Z => n1871);
   U2004 : INV_X2 port map( A => n2126, ZN => n2839);
   U2005 : INV_X2 port map( A => n1963, ZN => n2845);
   U2006 : INV_X4 port map( A => n2845, ZN => n1915);
   U2007 : INV_X1 port map( A => n1581, ZN => n2064);
   U2008 : NOR2_X4 port map( A1 => n3013, A2 => n4022, ZN => n164);
   U2009 : INV_X1 port map( A => DataP_add_S2_4_port, ZN => n1872);
   n1873 <= '1';
   n1874 <= '1';
   U2012 : OR2_X2 port map( A1 => n3167, A2 => n3166, ZN => 
                           DataP_alu_a_in_19_port);
   U2013 : AOI211_X2 port map( C1 => n2108, C2 => n2107, A => n2106, B => n2105
                           , ZN => n2120);
   U2014 : NAND3_X1 port map( A1 => n2449, A2 => n2448, A3 => n3270, ZN => 
                           n1875);
   U2015 : OAI221_X1 port map( B1 => n2122, B2 => n2121, C1 => n2122, C2 => 
                           n2120, A => n2119, ZN => n1876);
   U2016 : INV_X2 port map( A => n1844, ZN => n2995);
   U2017 : INV_X1 port map( A => n1893, ZN => n1878);
   U2018 : NAND4_X1 port map( A1 => n2388, A2 => n3231, A3 => n3230, A4 => 
                           n2335, ZN => DataP_alu_b_in_10_port);
   U2019 : BUF_X1 port map( A => n1581, Z => n1963);
   U2020 : OR2_X1 port map( A1 => DataP_alu_b_in_13_port, A2 => 
                           DataP_alu_b_in_12_port, ZN => n1881);
   U2021 : NAND2_X1 port map( A1 => n1875, A2 => n2225, ZN => n1882);
   U2022 : BUF_X1 port map( A => n1847, Z => n1883);
   U2023 : AND2_X1 port map( A1 => n2576, A2 => n1543, ZN => n3033);
   U2024 : INV_X1 port map( A => DataP_alu_a_in_18_port, ZN => n1884);
   U2025 : XNOR2_X1 port map( A => DataP_add_D_0_port, B => n1885, ZN => n3025)
                           ;
   U2026 : NAND3_X1 port map( A1 => n2994, A2 => n2998, A3 => n2155, ZN => 
                           n1887);
   U2027 : NAND3_X1 port map( A1 => n1568, A2 => n2998, A3 => n2155, ZN => 
                           n3193);
   U2028 : BUF_X1 port map( A => n3384, Z => n1888);
   U2029 : MUX2_X2 port map( A => n3690, B => n3701, S => n3689, Z => n3692);
   U2030 : NAND2_X1 port map( A1 => n3545, A2 => n2552, ZN => n1890);
   U2031 : INV_X1 port map( A => n1891, ZN => n1892);
   U2032 : OR2_X2 port map( A1 => n3076, A2 => n3075, ZN => 
                           DataP_alu_a_in_9_port);
   U2033 : AND2_X1 port map( A1 => n1978, A2 => n1979, ZN => n1893);
   U2034 : NOR3_X1 port map( A1 => n1582, A2 => n2389, A3 => n2333, ZN => n1896
                           );
   U2035 : NOR3_X1 port map( A1 => n1582, A2 => n2389, A3 => n2333, ZN => n1897
                           );
   U2036 : NOR3_X1 port map( A1 => n1582, A2 => n2389, A3 => n2333, ZN => n3263
                           );
   U2037 : OR2_X2 port map( A1 => n3079, A2 => n3078, ZN => 
                           DataP_alu_a_in_7_port);
   U2038 : NOR2_X1 port map( A1 => n1572, A2 => DataP_alu_b_in_10_port, ZN => 
                           n1898);
   U2039 : BUF_X1 port map( A => n3381, Z => n1899);
   U2040 : AND4_X1 port map( A1 => n1564, A2 => n2498, A3 => n3086, A4 => n3085
                           , ZN => n1900);
   U2041 : AND2_X1 port map( A1 => n1879, A2 => n2083, ZN => n1901);
   U2042 : AND2_X1 port map( A1 => n1572, A2 => n1863, ZN => n1902);
   U2043 : NOR2_X1 port map( A1 => n1901, A2 => n1902, ZN => n2088);
   U2044 : NOR2_X1 port map( A1 => n1966, A2 => n1910, ZN => n1903);
   U2045 : AOI21_X1 port map( B1 => n3039, B2 => n3038, A => n2157, ZN => n1904
                           );
   U2046 : NOR2_X1 port map( A1 => n1966, A2 => n1910, ZN => n2010);
   U2047 : NAND2_X1 port map( A1 => n3503, A2 => n3502, ZN => n1906);
   U2048 : AOI21_X1 port map( B1 => n1890, B2 => n2224, A => n2427, ZN => n1908
                           );
   U2049 : OR2_X1 port map( A1 => n3685, A2 => n3684, ZN => n1909);
   U2050 : OR2_X1 port map( A1 => n3685, A2 => n3684, ZN => n3708);
   U2051 : NAND4_X2 port map( A1 => n3098, A2 => n3099, A3 => n3096, A4 => 
                           n3097, ZN => n1910);
   U2052 : CLKBUF_X3 port map( A => n3327, Z => n3001);
   U2053 : AND4_X2 port map( A1 => n3103, A2 => n3102, A3 => n3101, A4 => n3100
                           , ZN => n2130);
   U2054 : AND2_X1 port map( A1 => n1635, A2 => DataP_B_s_6_port, ZN => n1911);
   U2055 : OR2_X2 port map( A1 => DataP_alu_b_in_17_port, A2 => n3510, ZN => 
                           n2538);
   U2056 : INV_X2 port map( A => n1580, ZN => DataP_alu_b_in_17_port);
   U2057 : OR2_X2 port map( A1 => n3170, A2 => n3169, ZN => 
                           DataP_alu_a_in_18_port);
   U2058 : NOR2_X2 port map( A1 => n1562, A2 => n3116, ZN => n1996);
   U2059 : NAND4_X1 port map( A1 => n3098, A2 => n3099, A3 => n3096, A4 => 
                           n3097, ZN => DataP_alu_b_in_2_port);
   U2060 : INV_X1 port map( A => DataP_alu_a_in_27_port, ZN => n1912);
   U2061 : OR2_X1 port map( A1 => n3137, A2 => n3136, ZN => 
                           DataP_alu_a_in_29_port);
   U2062 : OR2_X1 port map( A1 => n3161, A2 => n3160, ZN => 
                           DataP_alu_a_in_21_port);
   U2063 : OR2_X1 port map( A1 => n2302, A2 => n2145, ZN => 
                           DataP_alu_b_in_18_port);
   U2064 : OR2_X1 port map( A1 => n3134, A2 => n3133, ZN => 
                           DataP_alu_a_in_30_port);
   U2065 : OR2_X1 port map( A1 => n3128, A2 => n3127, ZN => 
                           DataP_alu_a_in_8_port);
   U2066 : INV_X1 port map( A => n2843, ZN => n1930);
   U2067 : BUF_X2 port map( A => n2990, Z => n2842);
   U2068 : INV_X2 port map( A => n2714, ZN => n1913);
   U2069 : INV_X2 port map( A => n2838, ZN => n1914);
   U2070 : BUF_X4 port map( A => n1907, Z => n1916);
   U2071 : INV_X1 port map( A => DataP_alu_b_in_28_port, ZN => n1917);
   U2072 : INV_X1 port map( A => n3510, ZN => n1918);
   U2073 : INV_X1 port map( A => n3911, ZN => n1919);
   U2074 : INV_X1 port map( A => DataP_alu_a_in_5_port, ZN => n1920);
   U2075 : INV_X1 port map( A => DataP_alu_a_in_8_port, ZN => n1921);
   U2076 : INV_X1 port map( A => DataP_alu_a_in_9_port, ZN => n1922);
   U2077 : INV_X1 port map( A => DataP_alu_a_in_31_port, ZN => n1923);
   U2078 : INV_X1 port map( A => DataP_alu_a_in_30_port, ZN => n1924);
   U2079 : INV_X1 port map( A => DataP_alu_a_in_29_port, ZN => n1925);
   U2080 : INV_X1 port map( A => DataP_alu_a_in_7_port, ZN => n1926);
   U2081 : INV_X1 port map( A => DataP_alu_a_in_13_port, ZN => n1927);
   U2082 : INV_X1 port map( A => DataP_alu_b_in_18_port, ZN => n1928);
   U2083 : INV_X1 port map( A => DataP_alu_a_in_25_port, ZN => n1929);
   U2084 : BUF_X2 port map( A => n2990, Z => n2841);
   U2085 : BUF_X2 port map( A => n2838, Z => n1931);
   U2086 : INV_X1 port map( A => DataP_alu_b_in_22_port, ZN => n1933);
   U2087 : INV_X1 port map( A => DataP_alu_b_in_29_port, ZN => n1934);
   U2088 : INV_X1 port map( A => DataP_alu_b_in_31_port, ZN => n1935);
   U2089 : INV_X1 port map( A => DataP_alu_b_in_26_port, ZN => n1936);
   U2090 : INV_X1 port map( A => DataP_alu_b_in_23_port, ZN => n1937);
   U2091 : INV_X1 port map( A => n3510, ZN => n1938);
   U2092 : INV_X1 port map( A => n3700, ZN => n1939);
   U2093 : AOI21_X1 port map( B1 => n3522, B2 => n1919, A => n1981, ZN => n1980
                           );
   U2094 : NOR2_X1 port map( A1 => n3910, A2 => n4019, ZN => n1981);
   U2095 : AND4_X1 port map( A1 => n2395, A2 => n2393, A3 => n2396, A4 => n2392
                           , ZN => n301);
   U2096 : AND4_X1 port map( A1 => n3260, A2 => n3259, A3 => n3258, A4 => n3257
                           , ZN => n2137);
   U2097 : INV_X2 port map( A => n3010, ZN => n1940);
   U2098 : OAI21_X1 port map( B1 => n3248, B2 => n1976, A => n1985, ZN => n3252
                           );
   U2099 : OR2_X1 port map( A1 => n3515, A2 => n3514, ZN => n2243);
   U2100 : NOR2_X1 port map( A1 => n3234, A2 => n1976, ZN => n3235);
   U2101 : AND2_X1 port map( A1 => n3416, A2 => n3415, ZN => n3456);
   U2102 : XNOR2_X1 port map( A => n3213, B => DataP_alu_a_in_7_port, ZN => 
                           n3387);
   U2103 : AND2_X1 port map( A1 => n3393, A2 => n3416, ZN => n3413);
   U2104 : AND2_X1 port map( A1 => n2282, A2 => n2283, ZN => n1958);
   U2105 : AND2_X1 port map( A1 => DataP_alu_a_in_10_port, A2 => n2357, ZN => 
                           n2356);
   U2106 : INV_X1 port map( A => DataP_alu_a_in_12_port, ZN => n1941);
   U2107 : INV_X1 port map( A => DataP_alu_a_in_3_port, ZN => n1942);
   U2108 : OR2_X1 port map( A1 => n3196, A2 => n3195, ZN => 
                           DataP_alu_a_in_10_port);
   U2109 : INV_X1 port map( A => DataP_alu_a_in_23_port, ZN => n1943);
   U2110 : OR2_X1 port map( A1 => n3158, A2 => n3157, ZN => 
                           DataP_alu_a_in_22_port);
   U2111 : OR2_X1 port map( A1 => n3175, A2 => n3174, ZN => 
                           DataP_alu_a_in_16_port);
   U2112 : INV_X1 port map( A => DataP_alu_a_in_20_port, ZN => n1944);
   U2113 : OR2_X1 port map( A1 => n3152, A2 => n3151, ZN => 
                           DataP_alu_a_in_24_port);
   U2114 : OR2_X1 port map( A1 => n3146, A2 => n3145, ZN => 
                           DataP_alu_a_in_26_port);
   U2115 : INV_X1 port map( A => DataP_alu_a_in_19_port, ZN => n1945);
   U2116 : OR2_X1 port map( A1 => n3140, A2 => n3139, ZN => 
                           DataP_alu_a_in_28_port);
   U2117 : INV_X2 port map( A => n1448, ZN => n4022);
   U2118 : INV_X1 port map( A => DataP_alu_b_in_19_port, ZN => n1946);
   U2119 : AND2_X1 port map( A1 => n3473, A2 => n1550, ZN => n2241);
   U2120 : INV_X1 port map( A => n2985, ZN => n2987);
   U2121 : INV_X1 port map( A => n1916, ZN => sra_131_SH_1_port);
   U2122 : BUF_X1 port map( A => n2990, Z => n2714);
   U2123 : INV_X1 port map( A => n1932, ZN => n1947);
   U2124 : BUF_X1 port map( A => n2990, Z => n2843);
   U2125 : INV_X2 port map( A => n2847, ZN => lt_x_135_B_4_port);
   U2126 : INV_X1 port map( A => DataP_alu_b_in_5_port, ZN => n1948);
   U2127 : INV_X1 port map( A => DataP_alu_b_in_21_port, ZN => n3442);
   U2128 : INV_X1 port map( A => DataP_alu_b_in_15_port, ZN => n1949);
   U2129 : INV_X1 port map( A => DataP_alu_b_in_7_port, ZN => n1950);
   U2130 : INV_X1 port map( A => DataP_alu_b_in_16_port, ZN => n1951);
   U2131 : INV_X2 port map( A => n2004, ZN => n2985);
   U2132 : INV_X1 port map( A => DataP_alu_b_in_21_port, ZN => n1952);
   U2133 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_6_port, ZN => 
                           n2152);
   U2134 : INV_X1 port map( A => n3071, ZN => n2469);
   U2135 : NOR2_X1 port map( A1 => n3674, A2 => n3911, ZN => n1982);
   U2136 : OAI21_X1 port map( B1 => n3948, B2 => n3947, A => Rst, ZN => n3949);
   U2137 : INV_X1 port map( A => n3065, ZN => n2471);
   U2138 : NAND2_X2 port map( A1 => n3229, A2 => Rst, ZN => n3910);
   U2139 : OR2_X2 port map( A1 => n3008, A2 => n3943, ZN => n3946);
   U2140 : INV_X1 port map( A => n3856, ZN => n3837);
   U2141 : AND2_X2 port map( A1 => WB_MUX_SEL_i_1_port, A2 => n294, ZN => n3943
                           );
   U2142 : CLKBUF_X1 port map( A => DataP_add_D_2_port, Z => n1955);
   U2143 : NOR2_X1 port map( A1 => IR_CU_27, A2 => IR_CU_26, ZN => n3856);
   U2144 : AOI21_X1 port map( B1 => n2413, B2 => n3691, A => n2226, ZN => n2567
                           );
   U2145 : AND3_X1 port map( A1 => n3692, A2 => n3705, A3 => n3691, ZN => n2153
                           );
   U2146 : NOR2_X2 port map( A1 => n3345, A2 => n3903, ZN => n3703);
   U2147 : BUF_X2 port map( A => n3706, Z => n3007);
   U2148 : NAND2_X2 port map( A1 => n3223, A2 => n3226, ZN => n3700);
   U2149 : NAND3_X1 port map( A1 => n1606, A2 => n3494, A3 => n3497, ZN => 
                           n3501);
   U2150 : OAI21_X1 port map( B1 => DataP_opcode_W_2_port, B2 => 
                           DataP_opcode_W_1_port, A => DataP_opcode_W_4_port, 
                           ZN => n1953);
   U2151 : AND2_X2 port map( A1 => n1563, A2 => n2136, ZN => n2503);
   U2152 : BUF_X1 port map( A => n3377, Z => n1954);
   U2153 : NAND3_X1 port map( A1 => n2449, A2 => n2448, A3 => n3270, ZN => 
                           n2290);
   U2154 : OAI21_X1 port map( B1 => n1957, B2 => n1918, A => n2366, ZN => n2419
                           );
   U2155 : INV_X1 port map( A => n1607, ZN => n2420);
   U2156 : NAND3_X1 port map( A1 => n3408, A2 => n2284, A3 => n1958, ZN => 
                           n3647);
   U2157 : NAND2_X1 port map( A1 => n3233, A2 => n3510, ZN => n1977);
   U2158 : NAND2_X1 port map( A1 => n1977, A2 => n2356, ZN => n2450);
   U2159 : BUF_X1 port map( A => n1557, Z => n1960);
   U2160 : BUF_X1 port map( A => n3669, Z => n1961);
   U2161 : NAND2_X1 port map( A1 => n3411, A2 => n3409, ZN => n1962);
   U2162 : NOR2_X1 port map( A1 => DataP_alu_b_in_13_port, A2 => 
                           DataP_alu_b_in_12_port, ZN => n3419);
   U2163 : NAND2_X1 port map( A1 => n1964, A2 => n3510, ZN => n2339);
   U2164 : XNOR2_X1 port map( A => n2009, B => DataP_alu_b_in_0_port, ZN => 
                           n1964);
   U2165 : NAND4_X1 port map( A1 => n3090, A2 => n3089, A3 => n3091, A4 => 
                           n3088, ZN => DataP_alu_b_in_0_port);
   U2166 : NAND4_X1 port map( A1 => n1564, A2 => n2498, A3 => n3086, A4 => 
                           n3085, ZN => n2506);
   U2167 : AND3_X2 port map( A1 => n1524, A2 => n1900, A3 => n2362, ZN => n2442
                           );
   U2168 : NAND3_X1 port map( A1 => n2500, A2 => n2499, A3 => n2152, ZN => 
                           n1965);
   U2169 : NAND2_X1 port map( A1 => n1637, A2 => n3214, ZN => n1966);
   U2170 : NAND2_X1 port map( A1 => n2002, A2 => n3494, ZN => n3467);
   U2171 : NAND2_X1 port map( A1 => n2425, A2 => n2540, ZN => n1967);
   U2172 : XNOR2_X1 port map( A => n3202, B => DataP_alu_a_in_3_port, ZN => 
                           n3678);
   U2173 : INV_X1 port map( A => n1968, ZN => n300);
   U2174 : OAI211_X1 port map( C1 => n1975, C2 => n2008, A => n1972, B => n1969
                           , ZN => n1968);
   U2175 : INV_X1 port map( A => n1970, ZN => n1969);
   U2176 : OAI21_X1 port map( B1 => n1975, B2 => n2550, A => n1971, ZN => n1970
                           );
   U2177 : INV_X1 port map( A => n3531, ZN => n1971);
   U2178 : NAND2_X1 port map( A1 => n2008, A2 => n1973, ZN => n1972);
   U2179 : AND2_X1 port map( A1 => n2550, A2 => n1974, ZN => n1973);
   U2180 : NOR2_X1 port map( A1 => n3524, A2 => n3674, ZN => n1974);
   U2181 : NAND2_X1 port map( A1 => n3524, A2 => n3691, ZN => n1975);
   U2182 : NAND2_X1 port map( A1 => n1906, A2 => n2552, ZN => n2008);
   U2183 : NAND2_X1 port map( A1 => n1978, A2 => n1979, ZN => n3458);
   U2184 : NAND2_X1 port map( A1 => n3422, A2 => n2512, ZN => n1978);
   U2185 : AOI21_X1 port map( B1 => n2418, B2 => n3691, A => n3522, ZN => n299)
                           ;
   U2186 : OAI221_X1 port map( B1 => n2059, B2 => n2058, C1 => n2059, C2 => 
                           n2057, A => n2056, ZN => n1983);
   U2187 : AOI21_X1 port map( B1 => n3354, B2 => n2438, A => n2437, ZN => n1984
                           );
   U2188 : AND2_X1 port map( A1 => n3488, A2 => n3509, ZN => n3490);
   U2189 : BUF_X1 port map( A => n3268, Z => n1985);
   U2190 : NAND2_X1 port map( A1 => n2002, A2 => n3456, ZN => n1986);
   U2191 : AOI21_X1 port map( B1 => n2131, B2 => n3465, A => n2421, ZN => n1988
                           );
   U2192 : NAND2_X1 port map( A1 => n2424, A2 => n2523, ZN => n1989);
   U2193 : INV_X1 port map( A => n2535, ZN => n1990);
   U2194 : BUF_X1 port map( A => n1909, Z => n1991);
   U2195 : XNOR2_X1 port map( A => n2293, B => n2292, ZN => n1992);
   U2196 : BUF_X1 port map( A => n3677, Z => n1993);
   U2197 : AND2_X1 port map( A1 => n1569, A2 => n2130, ZN => n1995);
   U2198 : AND2_X1 port map( A1 => n3088, A2 => n3084, ZN => n2498);
   U2199 : AND3_X1 port map( A1 => n2449, A2 => n3270, A3 => n2448, ZN => n1997
                           );
   U2200 : AND3_X2 port map( A1 => n3329, A2 => n1565, A3 => n2189, ZN => n2564
                           );
   U2201 : OAI211_X1 port map( C1 => n3441, C2 => n1531, A => n1559, B => n1960
                           , ZN => n1998);
   U2202 : INV_X1 port map( A => DataP_dest_M_2_port, ZN => n1999);
   U2203 : OAI211_X1 port map( C1 => n2492, C2 => n2494, A => n2489, B => n2491
                           , ZN => n2000);
   U2204 : BUF_X1 port map( A => n1587, Z => n2001);
   U2205 : NAND2_X1 port map( A1 => n1882, A2 => n2540, ZN => n2002);
   U2206 : NAND2_X1 port map( A1 => n1577, A2 => n1608, ZN => n2003);
   U2207 : NAND2_X1 port map( A1 => n1577, A2 => n1608, ZN => n3216);
   U2208 : NAND4_X1 port map( A1 => n1542, A2 => n1564, A3 => n3089, A4 => 
                           n3088, ZN => n2004);
   U2209 : INV_X1 port map( A => n1565, ZN => n2006);
   U2210 : OAI21_X1 port map( B1 => n2365, B2 => n2321, A => n2364, ZN => n2007
                           );
   U2211 : NAND2_X2 port map( A1 => n1845, A2 => n2143, ZN => n2561);
   U2212 : INV_X1 port map( A => n2843, ZN => n2844);
   U2213 : NAND4_X1 port map( A1 => n3087, A2 => n3085, A3 => n3086, A4 => 
                           n3084, ZN => n2009);
   U2214 : OAI21_X1 port map( B1 => n2380, B2 => n2577, A => n2379, ZN => n2011
                           );
   U2215 : OAI21_X1 port map( B1 => n2577, B2 => n2380, A => n2379, ZN => n3577
                           );
   U2216 : OAI211_X1 port map( C1 => n3212, C2 => n1517, A => n3211, B => n3387
                           , ZN => n2012);
   U2217 : OR2_X2 port map( A1 => n3113, A2 => n3114, ZN => 
                           DataP_alu_a_in_0_port);
   U2218 : OAI21_X1 port map( B1 => DataP_alu_b_in_30_port, B2 => n1924, A => 
                           n2013, ZN => n2048);
   U2219 : AOI211_X1 port map( C1 => DataP_alu_a_in_28_port, C2 => n1917, A => 
                           n2067, B => n2048, ZN => n2050);
   U2220 : AOI211_X1 port map( C1 => DataP_alu_a_in_24_port, C2 => n1550, A => 
                           n2113, B => n2060, ZN => n2014);
   U2221 : NAND2_X1 port map( A1 => n1573, A2 => n2014, ZN => n2059);
   U2222 : NOR2_X1 port map( A1 => DataP_alu_b_in_9_port, A2 => n1922, ZN => 
                           n2029);
   U2223 : NAND2_X1 port map( A1 => DataP_alu_a_in_13_port, A2 => n3396, ZN => 
                           n2015);
   U2224 : OAI211_X1 port map( C1 => n1880, C2 => n1941, A => n2035, B => n2015
                           , ZN => n2031);
   U2225 : NOR2_X1 port map( A1 => DataP_alu_b_in_8_port, A2 => n1921, ZN => 
                           n2017);
   U2226 : AOI21_X1 port map( B1 => n2358, B2 => DataP_alu_a_in_10_port, A => 
                           n2028, ZN => n2016);
   U2227 : OR4_X1 port map( A1 => n2029, A2 => n2031, A3 => n2017, A4 => n2063,
                           ZN => n2038);
   U2228 : OAI21_X1 port map( B1 => lt_x_134_B_5_port, B2 => n1920, A => 
                           lt_x_134_B_4_port, ZN => n2018);
   U2229 : OAI22_X1 port map( A1 => DataP_alu_a_in_4_port, A2 => n2018, B1 => 
                           DataP_alu_a_in_5_port, B2 => n1948, ZN => n2026);
   U2230 : AOI21_X1 port map( B1 => DataP_alu_a_in_6_port, B2 => n1611, A => 
                           n2072, ZN => n2025);
   U2231 : OAI21_X1 port map( B1 => n1612, B2 => n1996, A => n1537, ZN => n2019
                           );
   U2232 : OAI22_X1 port map( A1 => n1605, A2 => n2019, B1 => 
                           DataP_alu_a_in_1_port, B2 => n2126, ZN => n2020);
   U2233 : OAI221_X1 port map( B1 => n1963, B2 => n1942, C1 => n1910, C2 => 
                           n1561, A => n2020, ZN => n2021);
   U2234 : OAI221_X1 port map( B1 => DataP_alu_a_in_3_port, B2 => n2064, C1 => 
                           DataP_alu_a_in_2_port, C2 => n2076, A => n2021, ZN 
                           => n2022);
   U2235 : OAI21_X1 port map( B1 => lt_x_134_B_5_port, B2 => n1920, A => n2022,
                           ZN => n2023);
   U2236 : AOI221_X1 port map( B1 => n2026, B2 => n2025, C1 => n2024, C2 => 
                           n2025, A => n2080, ZN => n2037);
   U2237 : OAI21_X1 port map( B1 => n1860, B2 => n1927, A => n1880, ZN => n2027
                           );
   U2238 : AOI22_X1 port map( A1 => n2083, A2 => n1879, B1 => n1572, B2 => 
                           n1863, ZN => n2033);
   U2239 : NOR2_X1 port map( A1 => DataP_alu_a_in_8_port, A2 => n2029, ZN => 
                           n2030);
   U2240 : AOI22_X1 port map( A1 => n2030, A2 => DataP_alu_b_in_8_port, B1 => 
                           DataP_alu_b_in_9_port, B2 => n1922, ZN => n2032);
   U2241 : AOI221_X1 port map( B1 => n2063, B2 => n2033, C1 => n2032, C2 => 
                           n2033, A => n2031, ZN => n2034);
   U2242 : AOI211_X1 port map( C1 => n2035, C2 => n2092, A => n2090, B => n2034
                           , ZN => n2036);
   U2243 : OAI21_X1 port map( B1 => n2037, B2 => n2038, A => n2036, ZN => n2042
                           );
   U2244 : NOR2_X1 port map( A1 => DataP_alu_b_in_23_port, A2 => n1943, ZN => 
                           n2039);
   U2245 : AOI21_X1 port map( B1 => DataP_alu_a_in_22_port, B2 => n1933, A => 
                           n2039, ZN => n2047);
   U2246 : NAND2_X1 port map( A1 => DataP_alu_a_in_21_port, A2 => n1952, ZN => 
                           n2040);
   U2247 : OAI211_X1 port map( C1 => DataP_alu_b_in_20_port, C2 => n1944, A => 
                           n2047, B => n2040, ZN => n2046);
   U2248 : NOR2_X1 port map( A1 => DataP_alu_b_in_19_port, A2 => n1945, ZN => 
                           n2043);
   U2249 : AOI211_X1 port map( C1 => DataP_alu_a_in_16_port, C2 => n1951, A => 
                           n2046, B => n2061, ZN => n2041);
   U2250 : NAND3_X1 port map( A1 => n2042, A2 => n2125, A3 => n2041, ZN => 
                           n2058);
   U2251 : NOR2_X1 port map( A1 => DataP_alu_a_in_18_port, A2 => n2043, ZN => 
                           n2044);
   U2252 : NOR2_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => n2100, ZN => 
                           n2045);
   U2253 : OAI22_X1 port map( A1 => DataP_alu_a_in_28_port, A2 => n2110, B1 => 
                           DataP_alu_a_in_29_port, B2 => n1934, ZN => n2055);
   U2254 : AOI22_X1 port map( A1 => DataP_alu_b_in_26_port, A2 => n2112, B1 => 
                           DataP_alu_b_in_27_port, B2 => n1912, ZN => n2052);
   U2255 : NOR2_X1 port map( A1 => DataP_alu_a_in_24_port, A2 => n2113, ZN => 
                           n2049);
   U2256 : AOI22_X1 port map( A1 => DataP_alu_b_in_24_port, A2 => n2049, B1 => 
                           DataP_alu_b_in_25_port, B2 => n1929, ZN => n2051);
   U2257 : AOI221_X1 port map( B1 => n2060, B2 => n2052, C1 => n2051, C2 => 
                           n2052, A => n2062, ZN => n2054);
   U2258 : OAI21_X1 port map( B1 => DataP_alu_a_in_31_port, B2 => n1935, A => 
                           DataP_alu_b_in_30_port, ZN => n2053);
   U2259 : OAI221_X1 port map( B1 => n2059, B2 => n2058, C1 => n2059, C2 => 
                           n2057, A => n2056, ZN => DataP_ALU_C_comp_N24);
   U2260 : INV_X1 port map( A => lt_x_134_B_4_port, ZN => n2065);
   U2261 : AOI22_X1 port map( A1 => DataP_alu_a_in_15_port, A2 => n1949, B1 => 
                           DataP_alu_a_in_14_port, B2 => n1947, ZN => n2035);
   U2262 : INV_X1 port map( A => n2016, ZN => n2063);
   U2263 : INV_X1 port map( A => n2097, ZN => n2061);
   U2264 : INV_X1 port map( A => n2050, ZN => n2062);
   U2265 : NOR2_X1 port map( A1 => DataP_alu_b_in_29_port, A2 => n1925, ZN => 
                           n2067);
   U2266 : NAND2_X1 port map( A1 => DataP_alu_a_in_31_port, A2 => n1935, ZN => 
                           n2066);
   U2267 : OAI21_X1 port map( B1 => DataP_alu_b_in_30_port, B2 => n1924, A => 
                           n2066, ZN => n2109);
   U2268 : AOI211_X1 port map( C1 => DataP_alu_a_in_28_port, C2 => n1917, A => 
                           n2067, B => n2109, ZN => n2115);
   U2269 : NOR2_X1 port map( A1 => DataP_alu_b_in_25_port, A2 => n1929, ZN => 
                           n2113);
   U2270 : NOR2_X1 port map( A1 => n1912, A2 => DataP_alu_b_in_27_port, ZN => 
                           n2111);
   U2271 : AOI21_X1 port map( B1 => n1936, B2 => DataP_alu_a_in_26_port, A => 
                           n2111, ZN => n2068);
   U2272 : AOI211_X1 port map( C1 => DataP_alu_a_in_24_port, C2 => n1550, A => 
                           n2113, B => n2123, ZN => n2069);
   U2273 : NAND2_X1 port map( A1 => n2115, A2 => n2069, ZN => n2122);
   U2274 : NOR2_X1 port map( A1 => DataP_alu_b_in_9_port, A2 => n1922, ZN => 
                           n2084);
   U2275 : NOR2_X1 port map( A1 => DataP_alu_b_in_15_port, A2 => n1864, ZN => 
                           n2070);
   U2276 : AOI21_X1 port map( B1 => DataP_alu_a_in_14_port, B2 => n1947, A => 
                           n2070, ZN => n2093);
   U2277 : OAI211_X1 port map( C1 => n1880, C2 => n1941, A => n2093, B => n2015
                           , ZN => n2086);
   U2278 : OR4_X1 port map( A1 => n2084, A2 => n2086, A3 => n2017, A4 => n2063,
                           ZN => n2096);
   U2279 : OAI21_X1 port map( B1 => lt_x_134_B_5_port, B2 => n1920, A => 
                           lt_x_134_B_4_port, ZN => n2071);
   U2280 : OAI22_X1 port map( A1 => DataP_alu_a_in_4_port, A2 => n2071, B1 => 
                           DataP_alu_a_in_5_port, B2 => n1948, ZN => n2082);
   U2281 : NOR2_X1 port map( A1 => DataP_alu_b_in_7_port, A2 => n1926, ZN => 
                           n2072);
   U2282 : OAI21_X1 port map( B1 => n1963, B2 => n1942, A => n1910, ZN => n2076
                           );
   U2283 : OAI21_X1 port map( B1 => n1612, B2 => n1996, A => n2004, ZN => n2073
                           );
   U2284 : OAI22_X1 port map( A1 => n1605, A2 => n2073, B1 => 
                           DataP_alu_a_in_1_port, B2 => n2126, ZN => n2074);
   U2285 : OAI221_X1 port map( B1 => n1963, B2 => n1942, C1 => n1910, C2 => 
                           n1561, A => n2074, ZN => n2075);
   U2286 : OAI221_X1 port map( B1 => DataP_alu_a_in_3_port, B2 => n2127, C1 => 
                           DataP_alu_a_in_2_port, C2 => n2076, A => n2075, ZN 
                           => n2077);
   U2287 : OAI21_X1 port map( B1 => lt_x_134_B_5_port, B2 => n1920, A => n2077,
                           ZN => n2078);
   U2288 : AOI21_X1 port map( B1 => DataP_alu_a_in_4_port, B2 => n2847, A => 
                           n2078, ZN => n2081);
   U2289 : OAI21_X1 port map( B1 => DataP_alu_b_in_7_port, B2 => n1926, A => 
                           DataP_alu_b_in_6_port, ZN => n2079);
   U2290 : OAI22_X1 port map( A1 => DataP_alu_a_in_6_port, A2 => n2079, B1 => 
                           DataP_alu_a_in_7_port, B2 => n1950, ZN => n2080);
   U2291 : AOI221_X1 port map( B1 => n2082, B2 => n2025, C1 => n2081, C2 => 
                           n2025, A => n2080, ZN => n2095);
   U2292 : OAI22_X1 port map( A1 => DataP_alu_a_in_12_port, A2 => n2027, B1 => 
                           DataP_alu_a_in_13_port, B2 => n3396, ZN => n2092);
   U2293 : NOR2_X1 port map( A1 => DataP_alu_a_in_10_port, A2 => n2028, ZN => 
                           n2083);
   U2294 : NOR2_X1 port map( A1 => DataP_alu_a_in_8_port, A2 => n2084, ZN => 
                           n2085);
   U2295 : AOI22_X1 port map( A1 => DataP_alu_b_in_8_port, A2 => n2085, B1 => 
                           DataP_alu_b_in_9_port, B2 => n1922, ZN => n2087);
   U2296 : AOI221_X1 port map( B1 => n2063, B2 => n2088, C1 => n2087, C2 => 
                           n2088, A => n2086, ZN => n2091);
   U2297 : OAI21_X1 port map( B1 => DataP_alu_b_in_15_port, B2 => n1842, A => 
                           n1932, ZN => n2089);
   U2298 : OAI22_X1 port map( A1 => DataP_alu_a_in_14_port, A2 => n2089, B1 => 
                           n1841, B2 => n1949, ZN => n2090);
   U2299 : AOI211_X1 port map( C1 => n2093, C2 => n2092, A => n2090, B => n2091
                           , ZN => n2094);
   U2300 : OAI21_X1 port map( B1 => n2096, B2 => n2095, A => n2094, ZN => n2099
                           );
   U2301 : NOR2_X1 port map( A1 => DataP_alu_b_in_17_port, A2 => n1838, ZN => 
                           n2100);
   U2302 : AOI21_X1 port map( B1 => DataP_alu_a_in_22_port, B2 => n1933, A => 
                           n2039, ZN => n2108);
   U2303 : OAI211_X1 port map( C1 => DataP_alu_b_in_20_port, C2 => n1944, A => 
                           n2108, B => n2040, ZN => n2101);
   U2304 : AOI21_X1 port map( B1 => n1928, B2 => DataP_alu_a_in_18_port, A => 
                           n2043, ZN => n2097);
   U2305 : AOI211_X1 port map( C1 => DataP_alu_a_in_16_port, C2 => n1951, A => 
                           n2101, B => n2061, ZN => n2098);
   U2306 : NAND3_X1 port map( A1 => n2099, A2 => n2125, A3 => n2098, ZN => 
                           n2121);
   U2307 : AOI22_X1 port map( A1 => DataP_alu_b_in_18_port, A2 => n2044, B1 => 
                           DataP_alu_b_in_19_port, B2 => n1945, ZN => n2103);
   U2308 : AOI22_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n2045, B1 => 
                           DataP_alu_b_in_17_port, B2 => n1838, ZN => n2102);
   U2309 : AOI221_X1 port map( B1 => n2061, B2 => n2103, C1 => n2102, C2 => 
                           n2103, A => n2101, ZN => n2106);
   U2310 : OAI21_X1 port map( B1 => DataP_alu_b_in_23_port, B2 => n1943, A => 
                           DataP_alu_b_in_22_port, ZN => n2104);
   U2311 : OAI22_X1 port map( A1 => DataP_alu_a_in_22_port, A2 => n2104, B1 => 
                           DataP_alu_a_in_23_port, B2 => n1937, ZN => n2105);
   U2312 : OAI21_X1 port map( B1 => DataP_alu_b_in_29_port, B2 => n1925, A => 
                           DataP_alu_b_in_28_port, ZN => n2110);
   U2313 : NOR2_X1 port map( A1 => DataP_alu_a_in_26_port, A2 => n2111, ZN => 
                           n2112);
   U2314 : AOI22_X1 port map( A1 => DataP_alu_b_in_26_port, A2 => n2112, B1 => 
                           DataP_alu_b_in_27_port, B2 => n1912, ZN => n2117);
   U2315 : NOR2_X1 port map( A1 => DataP_alu_a_in_24_port, A2 => n2113, ZN => 
                           n2114);
   U2316 : AOI22_X1 port map( A1 => DataP_alu_b_in_24_port, A2 => n2114, B1 => 
                           DataP_alu_b_in_25_port, B2 => n1929, ZN => n2116);
   U2317 : OAI21_X1 port map( B1 => DataP_alu_b_in_31_port, B2 => n1923, A => 
                           DataP_alu_b_in_30_port, ZN => n2118);
   U2318 : INV_X1 port map( A => n1612, ZN => n2126);
   U2319 : INV_X1 port map( A => DataP_alu_b_in_3_port, ZN => n2127);
   U2320 : INV_X1 port map( A => n2068, ZN => n2123);
   U2321 : INV_X1 port map( A => n2100, ZN => n2125);
   U2322 : INV_X1 port map( A => n2115, ZN => n2124);
   U2323 : NAND2_X1 port map( A1 => n1566, A2 => n2313, ZN => n3329);
   U2324 : AND2_X1 port map( A1 => n3021, A2 => n3022, ZN => n2480);
   U2325 : NAND4_X1 port map( A1 => n3107, A2 => n3106, A3 => n3105, A4 => 
                           n3104, ZN => DataP_alu_b_in_5_port);
   U2326 : OR2_X1 port map( A1 => n2231, A2 => n3003, ZN => n3093);
   U2327 : OR2_X1 port map( A1 => n3003, A2 => n2227, ZN => n3105);
   U2328 : INV_X1 port map( A => n1844, ZN => n2996);
   U2329 : OR2_X1 port map( A1 => n3070, A2 => n3012, ZN => n3071);
   U2330 : AND3_X1 port map( A1 => n3655, A2 => n3654, A3 => n3653, ZN => n333)
                           ;
   U2331 : INV_X1 port map( A => sra_131_SH_4_port, ZN => n2847);
   U2332 : OR2_X1 port map( A1 => n3172, A2 => n3171, ZN => 
                           DataP_alu_a_in_17_port);
   U2333 : OR2_X1 port map( A1 => n3953, A2 => CU_I_cw_7_port, ZN => n3947);
   U2334 : NOR3_X1 port map( A1 => n3795, A2 => n3955, A3 => n3837, ZN => n3953
                           );
   U2335 : BUF_X1 port map( A => n1910, Z => n2990);
   U2336 : INV_X1 port map( A => n3425, ZN => DataP_alu_b_in_16_port);
   U2337 : INV_X1 port map( A => n2005, ZN => n3003);
   U2338 : OR2_X1 port map( A1 => n3026, A2 => n1892, ZN => n3062);
   U2339 : INV_X1 port map( A => n3987, ZN => n492);
   U2340 : INV_X1 port map( A => n3988, ZN => n491);
   U2341 : NOR2_X1 port map( A1 => n3853, A2 => n3852, ZN => CU_I_cw_7_port);
   U2342 : INV_X1 port map( A => n3951, ZN => n3853);
   U2343 : INV_X1 port map( A => n3956, ZN => n3948);
   U2344 : INV_X1 port map( A => n3695, ZN => n3675);
   U2345 : INV_X1 port map( A => n3674, ZN => n3691);
   U2346 : AND3_X1 port map( A1 => n3201, A2 => n3689, A3 => n3200, ZN => n3674
                           );
   U2347 : OR2_X1 port map( A1 => n3002, A2 => n2229, ZN => n3101);
   U2348 : INV_X1 port map( A => n3985, ZN => n494);
   U2349 : INV_X1 port map( A => n3989, ZN => n490);
   U2350 : INV_X1 port map( A => n3986, ZN => n493);
   U2351 : NOR2_X1 port map( A1 => n487, A2 => n3949, ZN => DataP_add_S2_2_port
                           );
   U2352 : NOR2_X1 port map( A1 => n486, A2 => n3949, ZN => DataP_add_S2_1_port
                           );
   U2353 : INV_X1 port map( A => n2923, ZN => n2981);
   U2354 : BUF_X1 port map( A => n3703, Z => n3006);
   U2355 : AND4_X1 port map( A1 => n3037, A2 => n1869, A3 => n1999, A4 => n529,
                           ZN => n2157);
   U2356 : NOR2_X1 port map( A1 => n489, A2 => n3949, ZN => DataP_add_S2_4_port
                           );
   U2357 : NOR2_X1 port map( A1 => n485, A2 => n3949, ZN => DataP_add_S2_0_port
                           );
   U2358 : NOR2_X1 port map( A1 => n488, A2 => n3949, ZN => DataP_add_S2_3_port
                           );
   U2359 : NAND2_X1 port map( A1 => n516, A2 => n510, ZN => n3795);
   U2360 : NOR2_X1 port map( A1 => n504, A2 => n497, ZN => n3966);
   U2361 : AND3_X2 port map( A1 => n2453, A2 => n3272, A3 => n2451, ZN => n3270
                           );
   U2362 : OR2_X1 port map( A1 => n2232, A2 => n3003, ZN => n3097);
   U2363 : NOR2_X1 port map( A1 => n3795, A2 => n2141, ZN => n144);
   U2364 : AND2_X1 port map( A1 => BR_EN_i, A2 => n3901, ZN => n3711);
   U2365 : NAND2_X1 port map( A1 => n514, A2 => n515, ZN => n3955);
   U2366 : NAND3_X1 port map( A1 => n3966, A2 => n144, A3 => n2129, ZN => n3956
                           );
   U2367 : NAND2_X2 port map( A1 => n3711, A2 => Rst, ZN => n3911);
   U2368 : NOR2_X1 port map( A1 => n3221, A2 => n3903, ZN => n3706);
   U2369 : OR2_X2 port map( A1 => n3474, A2 => DataP_alu_a_in_26_port, ZN => 
                           n3504);
   U2370 : AND3_X2 port map( A1 => n3468, A2 => n1933, A3 => n1937, ZN => n2133
                           );
   U2371 : AND4_X2 port map( A1 => n3081, A2 => n3083, A3 => n3080, A4 => n3082
                           , ZN => n3214);
   U2372 : AND2_X1 port map( A1 => n3198, A2 => ALU_OPCODE_i_1_port, ZN => 
                           n3224);
   U2373 : BUF_X1 port map( A => n4021, Z => n3009);
   U2374 : NOR2_X1 port map( A1 => n1448, A2 => n3013, ZN => n4021);
   U2375 : INV_X1 port map( A => Rst, ZN => n3014);
   U2376 : INV_X1 port map( A => Rst, ZN => n3013);
   U2377 : INV_X1 port map( A => DataP_npc_mux_sel, ZN => n3010);
   U2378 : BUF_X1 port map( A => n3944, Z => n3008);
   U2379 : NOR2_X1 port map( A1 => WB_MUX_SEL_i_1_port, A2 => n294, ZN => n3944
                           );
   U2380 : INV_X1 port map( A => n3965, ZN => n3981);
   U2381 : NOR2_X1 port map( A1 => n3711, A2 => DataP_wrong_br, ZN => n1448);
   U2382 : AND2_X2 port map( A1 => n2503, A2 => n2133, ZN => n3488);
   U2383 : AND4_X2 port map( A1 => n3315, A2 => n2520, A3 => n3313, A4 => n3314
                           , ZN => n3425);
   U2384 : AND4_X2 port map( A1 => n3305, A2 => n2519, A3 => n3303, A4 => n3304
                           , ZN => n3424);
   U2385 : AND2_X2 port map( A1 => n3420, A2 => n3421, ZN => n3437);
   U2386 : OR2_X2 port map( A1 => n3187, A2 => n3186, ZN => 
                           DataP_alu_a_in_12_port);
   U2387 : OR2_X2 port map( A1 => n3122, A2 => n3121, ZN => 
                           DataP_alu_a_in_5_port);
   U2388 : INV_X2 port map( A => n3694, ZN => n3697);
   U2389 : INV_X2 port map( A => n1857, ZN => n2991);
   U2390 : BUF_X2 port map( A => n3194, Z => n2563);
   U2391 : OR2_X2 port map( A1 => n3125, A2 => n3124, ZN => 
                           DataP_alu_a_in_6_port);
   U2392 : INV_X2 port map( A => n1857, ZN => n2992);
   U2393 : BUF_X2 port map( A => n1887, Z => n3000);
   U2394 : NOR4_X1 port map( A1 => n443, A2 => ALU_OPCODE_i_3_port, A3 => 
                           ALU_OPCODE_i_2_port, A4 => ALU_OPCODE_i_1_port, ZN 
                           => n3901);
   U2395 : NAND2_X1 port map( A1 => n3226, A2 => ALU_OPCODE_i_0_port, ZN => 
                           n3709);
   U2396 : AOI211_X1 port map( C1 => n3675, C2 => DataP_ALU_C_shifter_N83, A =>
                           n3369, B => n3368, ZN => n358);
   U2397 : AND2_X1 port map( A1 => DataP_ALU_C_shifter_N51, A2 => n3006, ZN => 
                           n3368);
   U2398 : OAI211_X1 port map( C1 => n3674, C2 => n3367, A => n3366, B => n3365
                           , ZN => n3369);
   U2399 : AOI21_X1 port map( B1 => n1939, B2 => n3364, A => n3363, ZN => n3365
                           );
   U2400 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N19, A2 => n3007, ZN =>
                           n3366);
   U2401 : INV_X1 port map( A => n2618, ZN => n2703);
   U2402 : NAND2_X1 port map( A1 => n3359, A2 => n3358, ZN => n3360);
   U2403 : INV_X1 port map( A => DataP_add_S2_1_port, ZN => n2559);
   U2404 : AOI21_X1 port map( B1 => n2990, B2 => n3693, A => n3697, ZN => n3373
                           );
   U2405 : INV_X1 port map( A => n2673, ZN => n2704);
   U2406 : OAI22_X1 port map( A1 => n355, A2 => n3911, B1 => n3994, B2 => n3910
                           , ZN => DataP_PC_reg_N6);
   U2407 : INV_X1 port map( A => n2691, ZN => n2705);
   U2408 : OAI22_X1 port map( A1 => n356, A2 => n3911, B1 => n3993, B2 => n3910
                           , ZN => DataP_PC_reg_N5);
   U2409 : AOI21_X1 port map( B1 => n2330, B2 => n3694, A => n3679, ZN => n3680
                           );
   U2410 : INV_X1 port map( A => DataP_add_S2_3_port, ZN => n2557);
   U2411 : INV_X1 port map( A => DataP_add_S2_0_port, ZN => n2558);
   U2412 : OAI22_X1 port map( A1 => n353, A2 => n3911, B1 => n3996, B2 => n3910
                           , ZN => DataP_PC_reg_N8);
   U2413 : NAND2_X1 port map( A1 => DataP_alu_b_in_6_port, A2 => n3660, ZN => 
                           n2363);
   U2414 : AOI22_X1 port map( A1 => n3388, A2 => DataP_alu_b_in_7_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_7_port, ZN => n3389);
   U2415 : OAI21_X1 port map( B1 => n1926, B2 => n3671, A => n3694, ZN => n3388
                           );
   U2416 : INV_X1 port map( A => n2694, ZN => n2706);
   U2417 : INV_X1 port map( A => n1888, ZN => n3386);
   U2418 : OAI21_X1 port map( B1 => n3670, B2 => n3378, A => n1954, ZN => n3383
                           );
   U2419 : INV_X1 port map( A => n3376, ZN => n3378);
   U2420 : NAND2_X1 port map( A1 => n2001, A2 => n3375, ZN => n3670);
   U2421 : OAI22_X1 port map( A1 => n345, A2 => n3911, B1 => n3998, B2 => n3910
                           , ZN => DataP_PC_reg_N10);
   U2422 : AOI21_X1 port map( B1 => n3663, B2 => n1939, A => n3697, ZN => n3662
                           );
   U2423 : NOR2_X1 port map( A1 => n1939, A2 => n3697, ZN => n3661);
   U2424 : INV_X1 port map( A => n2695, ZN => n2707);
   U2425 : AOI22_X1 port map( A1 => n3227, A2 => DataP_alu_b_in_9_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_9_port, ZN => n3228);
   U2426 : OAI21_X1 port map( B1 => n1922, B2 => n3671, A => n3694, ZN => n3227
                           );
   U2427 : INV_X1 port map( A => n2696, ZN => n2708);
   U2428 : INV_X1 port map( A => n3657, ZN => n3217);
   U2429 : NOR2_X1 port map( A1 => n3911, A2 => n443, ZN => n2347);
   U2430 : INV_X1 port map( A => n3243, ZN => n340);
   U2431 : OAI211_X1 port map( C1 => n3674, C2 => n3242, A => n3241, B => n3240
                           , ZN => n3243);
   U2432 : AOI22_X1 port map( A1 => n3006, A2 => DataP_ALU_C_shifter_N60, B1 =>
                           DataP_ALU_C_shifter_N92, B2 => n3675, ZN => n3240);
   U2433 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N28, B2 => n3007, A => 
                           n3239, ZN => n3241);
   U2434 : OAI21_X1 port map( B1 => n3700, B2 => n3283, A => n3238, ZN => n3239
                           );
   U2435 : AOI22_X1 port map( A1 => n3237, A2 => n1879, B1 => n3697, B2 => 
                           DataP_alu_a_in_10_port, ZN => n3238);
   U2436 : OAI21_X1 port map( B1 => n3236, B2 => n3671, A => n3694, ZN => n3237
                           );
   U2437 : INV_X1 port map( A => n2654, ZN => n2697);
   U2438 : XNOR2_X1 port map( A => n3248, B => n3235, ZN => n3242);
   U2439 : INV_X1 port map( A => n1985, ZN => n3234);
   U2440 : NAND2_X1 port map( A1 => n2343, A2 => n2342, ZN => n296);
   U2441 : INV_X1 port map( A => DataP_ALU_C_comp_N24, ZN => n3352);
   U2442 : NAND2_X1 port map( A1 => n2345, A2 => n2344, ZN => n2343);
   U2443 : NOR3_X1 port map( A1 => n2431, A2 => n2349, A3 => n443, ZN => n2344)
                           ;
   U2444 : NAND4_X1 port map( A1 => n3340, A2 => n3339, A3 => n3338, A4 => 
                           n3337, ZN => n3357);
   U2445 : OAI21_X1 port map( B1 => n3336, B2 => n3697, A => n3335, ZN => n3337
                           );
   U2446 : AOI21_X1 port map( B1 => n3674, B2 => n3700, A => n3361, ZN => n3336
                           );
   U2447 : NAND2_X1 port map( A1 => n3361, A2 => n3693, ZN => n3338);
   U2448 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N50, A2 => n3006, ZN =>
                           n3340);
   U2449 : OAI21_X1 port map( B1 => n3350, B2 => n3356, A => n3349, ZN => n3351
                           );
   U2450 : INV_X1 port map( A => n3355, ZN => n3349);
   U2451 : INV_X1 port map( A => n1876, ZN => n3350);
   U2452 : AND2_X1 port map( A1 => n3353, A2 => n3223, ZN => n3341);
   U2453 : NAND2_X1 port map( A1 => n2516, A2 => n2369, ZN => n3353);
   U2454 : INV_X1 port map( A => n3374, ZN => n3316);
   U2455 : XNOR2_X1 port map( A => DataP_alu_a_in_2_port, B => n2844, ZN => 
                           n3374);
   U2456 : XNOR2_X1 port map( A => DataP_alu_a_in_4_port, B => 
                           lt_x_134_B_4_port, ZN => n3673);
   U2457 : XNOR2_X1 port map( A => DataP_alu_a_in_7_port, B => 
                           DataP_alu_b_in_7_port, ZN => n3390);
   U2458 : XNOR2_X1 port map( A => DataP_alu_a_in_6_port, B => 
                           DataP_alu_b_in_6_port, ZN => n3668);
   U2459 : INV_X1 port map( A => n3361, ZN => n3317);
   U2460 : AND2_X1 port map( A1 => n2517, A2 => n3904, ZN => n2516);
   U2461 : NOR3_X1 port map( A1 => n3299, A2 => n3364, A3 => n3298, ZN => n3904
                           );
   U2462 : NAND4_X1 port map( A1 => n3518, A2 => n3527, A3 => n3477, A4 => 
                           n3536, ZN => n3298);
   U2463 : INV_X1 port map( A => n3547, ZN => n3299);
   U2464 : NOR2_X1 port map( A1 => n3905, A2 => n2518, ZN => n2517);
   U2465 : NAND4_X1 port map( A1 => n3586, A2 => n3908, A3 => n3909, A4 => 
                           n3570, ZN => n2518);
   U2466 : AND4_X1 port map( A1 => n3605, A2 => n3284, A3 => n3283, A4 => n3282
                           , ZN => n2222);
   U2467 : XNOR2_X1 port map( A => DataP_alu_a_in_9_port, B => 
                           DataP_alu_b_in_9_port, ZN => n3282);
   U2468 : XNOR2_X1 port map( A => DataP_alu_a_in_10_port, B => n1879, ZN => 
                           n3283);
   U2469 : OAI21_X1 port map( B1 => n3346, B2 => n3345, A => n3344, ZN => n3347
                           );
   U2470 : OAI22_X1 port map( A1 => n317, A2 => n3911, B1 => n3910, B2 => n4010
                           , ZN => DataP_PC_reg_N22);
   U2471 : INV_X1 port map( A => DataP_npc_20_port, ZN => n4010);
   U2472 : AOI21_X1 port map( B1 => n3601, B2 => n3691, A => n3600, ZN => n317)
                           ;
   U2473 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N38, A2 => n3007, ZN =>
                           n3597);
   U2474 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N70, B2 => n3703, A => 
                           n3596, ZN => n3598);
   U2475 : OAI211_X1 port map( C1 => n3907, C2 => n3700, A => n3595, B => n3594
                           , ZN => n3596);
   U2476 : NAND2_X1 port map( A1 => DataP_alu_a_in_20_port, A2 => n3697, ZN => 
                           n3594);
   U2477 : OAI211_X1 port map( C1 => DataP_alu_a_in_20_port, C2 => n3697, A => 
                           DataP_alu_b_in_20_port, B => n3660, ZN => n3595);
   U2478 : XNOR2_X1 port map( A => DataP_alu_a_in_20_port, B => 
                           DataP_alu_b_in_20_port, ZN => n3907);
   U2479 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N102, A2 => n3675, ZN 
                           => n3599);
   U2480 : OAI22_X1 port map( A1 => n326, A2 => n3911, B1 => n3910, B2 => n4006
                           , ZN => DataP_PC_reg_N18);
   U2481 : INV_X1 port map( A => DataP_npc_16_port, ZN => n4006);
   U2482 : AOI21_X1 port map( B1 => n3630, B2 => n3691, A => n3629, ZN => n326)
                           ;
   U2483 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N34, A2 => n3007, ZN =>
                           n3626);
   U2484 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N98, A2 => n3675, ZN =>
                           n3627);
   U2485 : INV_X1 port map( A => n2894, ZN => DataP_ALU_C_shifter_N98);
   U2486 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N66, B2 => n3703, A => 
                           n3625, ZN => n3628);
   U2487 : OAI211_X1 port map( C1 => n3624, C2 => n3700, A => n3623, B => n3622
                           , ZN => n3625);
   U2488 : OAI21_X1 port map( B1 => DataP_alu_a_in_16_port, B2 => 
                           DataP_alu_b_in_16_port, A => n3697, ZN => n3622);
   U2489 : XNOR2_X1 port map( A => DataP_alu_a_in_16_port, B => 
                           DataP_alu_b_in_16_port, ZN => n3624);
   U2490 : INV_X1 port map( A => n3280, ZN => n337);
   U2491 : OAI211_X1 port map( C1 => n3279, C2 => n3674, A => n3278, B => n3277
                           , ZN => n3280);
   U2492 : AOI22_X1 port map( A1 => DataP_ALU_C_shifter_N30, A2 => n3007, B1 =>
                           n3675, B2 => DataP_ALU_C_shifter_N94, ZN => n3277);
   U2493 : INV_X1 port map( A => n2664, ZN => n2699);
   U2494 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N62, B2 => n3006, A => 
                           n3276, ZN => n3278);
   U2495 : OAI211_X1 port map( C1 => n3284, C2 => n3700, A => n3275, B => n3274
                           , ZN => n3276);
   U2496 : OAI21_X1 port map( B1 => DataP_alu_a_in_12_port, B2 => n1880, A => 
                           n3697, ZN => n3275);
   U2497 : XNOR2_X1 port map( A => DataP_alu_a_in_12_port, B => n1880, ZN => 
                           n3284);
   U2498 : NAND2_X1 port map( A1 => n3642, A2 => n3640, ZN => n3273);
   U2499 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N29, A2 => n3007, ZN =>
                           n3257);
   U2500 : INV_X1 port map( A => n2658, ZN => n2698);
   U2501 : AOI21_X1 port map( B1 => n3318, B2 => n1939, A => n3256, ZN => n3258
                           );
   U2502 : OAI22_X1 port map( A1 => n3255, A2 => n3254, B1 => n1863, B2 => 
                           n3694, ZN => n3256);
   U2503 : AOI21_X1 port map( B1 => DataP_alu_a_in_11_port, B2 => n3693, A => 
                           n3697, ZN => n3255);
   U2504 : AOI22_X1 port map( A1 => n3006, A2 => DataP_ALU_C_shifter_N61, B1 =>
                           DataP_ALU_C_shifter_N93, B2 => n3675, ZN => n3259);
   U2505 : NAND2_X1 port map( A1 => n3253, A2 => n3691, ZN => n3260);
   U2506 : XNOR2_X1 port map( A => n3252, B => n3270, ZN => n3253);
   U2507 : NAND2_X1 port map( A1 => n2012, A2 => n3265, ZN => n3659);
   U2508 : OAI22_X1 port map( A1 => n333, A2 => n3911, B1 => n3910, B2 => n4003
                           , ZN => DataP_PC_reg_N15);
   U2509 : INV_X1 port map( A => DataP_npc_13_port, ZN => n4003);
   U2510 : AOI22_X1 port map( A1 => n3006, A2 => DataP_ALU_C_shifter_N63, B1 =>
                           DataP_ALU_C_shifter_N95, B2 => n3675, ZN => n3653);
   U2511 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N31, B2 => n3007, A => 
                           n3652, ZN => n3654);
   U2512 : OAI211_X1 port map( C1 => n3651, C2 => n3700, A => n3650, B => n3649
                           , ZN => n3652);
   U2513 : INV_X1 port map( A => n2671, ZN => n2700);
   U2514 : OAI211_X1 port map( C1 => n3648, C2 => n3647, A => n3646, B => n3691
                           , ZN => n3655);
   U2515 : OAI211_X1 port map( C1 => n3645, C2 => n3644, A => n3643, B => n3642
                           , ZN => n3646);
   U2516 : NAND2_X1 port map( A1 => n1601, A2 => n3640, ZN => n3643);
   U2517 : NOR2_X1 port map( A1 => n1997, A2 => n3639, ZN => n3648);
   U2518 : OAI22_X1 port map( A1 => n301, A2 => n3911, B1 => n3910, B2 => n4017
                           , ZN => DataP_PC_reg_N29);
   U2519 : INV_X1 port map( A => DataP_npc_27_port, ZN => n4017);
   U2520 : NOR2_X1 port map( A1 => n2397, A2 => n3481, ZN => n2396);
   U2521 : OAI211_X1 port map( C1 => n3695, C2 => n2926, A => n3480, B => n3479
                           , ZN => n3481);
   U2522 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N77, B2 => n3006, A => 
                           n3478, ZN => n3479);
   U2523 : OAI21_X1 port map( B1 => n3700, B2 => n3477, A => n3476, ZN => n3478
                           );
   U2524 : AOI22_X1 port map( A1 => n3475, A2 => DataP_alu_b_in_27_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_27_port, ZN => n3476);
   U2525 : OAI21_X1 port map( B1 => n1912, B2 => n3671, A => n3694, ZN => n3475
                           );
   U2526 : XNOR2_X1 port map( A => DataP_alu_a_in_27_port, B => 
                           DataP_alu_b_in_27_port, ZN => n3477);
   U2527 : NAND2_X1 port map( A1 => n2400, A2 => n2398, ZN => n2397);
   U2528 : NAND2_X1 port map( A1 => n1867, A2 => n2399, ZN => n2398);
   U2529 : NOR2_X1 port map( A1 => n3504, A2 => n3674, ZN => n2399);
   U2530 : NAND2_X1 port map( A1 => n2401, A2 => n2553, ZN => n2400);
   U2531 : OR2_X1 port map( A1 => n2422, A2 => n2394, ZN => n2393);
   U2532 : NOR2_X1 port map( A1 => n1867, A2 => n2402, ZN => n2401);
   U2533 : NAND2_X1 port map( A1 => n3504, A2 => n3691, ZN => n2402);
   U2534 : OAI22_X1 port map( A1 => n313, A2 => n3911, B1 => n3910, B2 => n4011
                           , ZN => DataP_PC_reg_N23);
   U2535 : INV_X1 port map( A => DataP_npc_21_port, ZN => n4011);
   U2536 : AOI21_X1 port map( B1 => n3591, B2 => n3691, A => n3590, ZN => n313)
                           ;
   U2537 : OAI21_X1 port map( B1 => n3695, B2 => n3589, A => n3588, ZN => n3590
                           );
   U2538 : AOI21_X1 port map( B1 => n3007, B2 => DataP_ALU_C_shifter_N39, A => 
                           n3587, ZN => n3588);
   U2539 : OAI211_X1 port map( C1 => n3700, C2 => n3586, A => n3585, B => n3584
                           , ZN => n3587);
   U2540 : AOI22_X1 port map( A1 => n3583, A2 => DataP_alu_b_in_21_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_21_port, ZN => n3584);
   U2541 : OAI21_X1 port map( B1 => n1589, B2 => n3671, A => n3694, ZN => n3583
                           );
   U2542 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N71, A2 => n3006, ZN =>
                           n3585);
   U2543 : XNOR2_X1 port map( A => DataP_alu_a_in_21_port, B => 
                           DataP_alu_b_in_21_port, ZN => n3586);
   U2544 : INV_X1 port map( A => DataP_ALU_C_shifter_N103, ZN => n3589);
   U2545 : AOI21_X1 port map( B1 => n1989, B2 => n3580, A => n3579, ZN => n3581
                           );
   U2546 : INV_X1 port map( A => n1560, ZN => n3579);
   U2547 : OAI22_X1 port map( A1 => n304, A2 => n3911, B1 => n3910, B2 => n4015
                           , ZN => DataP_PC_reg_N27);
   U2548 : INV_X1 port map( A => DataP_npc_25_port, ZN => n4015);
   U2549 : AOI21_X1 port map( B1 => n3553, B2 => n3691, A => n3552, ZN => n304)
                           ;
   U2550 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N75, B2 => n3703, A => 
                           n3548, ZN => n3549);
   U2551 : XNOR2_X1 port map( A => DataP_alu_a_in_25_port, B => 
                           DataP_alu_b_in_25_port, ZN => n3547);
   U2552 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N43, A2 => n3007, ZN =>
                           n3550);
   U2553 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N107, A2 => n3675, ZN 
                           => n3551);
   U2554 : INV_X1 port map( A => n2922, ZN => n2984);
   U2555 : NOR2_X1 port map( A1 => n2556, A2 => n3544, ZN => n3546);
   U2556 : OAI22_X1 port map( A1 => n311, A2 => n3911, B1 => n3910, B2 => n4012
                           , ZN => DataP_PC_reg_N24);
   U2557 : INV_X1 port map( A => DataP_npc_22_port, ZN => n4012);
   U2558 : AOI21_X1 port map( B1 => n3575, B2 => n3691, A => n3574, ZN => n311)
                           ;
   U2559 : OAI21_X1 port map( B1 => n3695, B2 => n3573, A => n3572, ZN => n3574
                           );
   U2560 : AOI21_X1 port map( B1 => n3007, B2 => DataP_ALU_C_shifter_N40, A => 
                           n3571, ZN => n3572);
   U2561 : OAI211_X1 port map( C1 => n3700, C2 => n3570, A => n3569, B => n3568
                           , ZN => n3571);
   U2562 : AOI22_X1 port map( A1 => n3567, A2 => DataP_alu_b_in_22_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_22_port, ZN => n3568);
   U2563 : OAI21_X1 port map( B1 => n3566, B2 => n3671, A => n3694, ZN => n3567
                           );
   U2564 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N72, A2 => n3006, ZN =>
                           n3569);
   U2565 : XNOR2_X1 port map( A => DataP_alu_a_in_22_port, B => 
                           DataP_alu_b_in_22_port, ZN => n3570);
   U2566 : INV_X1 port map( A => DataP_ALU_C_shifter_N104, ZN => n3573);
   U2567 : XNOR2_X1 port map( A => n1639, B => n3564, ZN => n3575);
   U2568 : OAI22_X1 port map( A1 => n308, A2 => n3911, B1 => n3910, B2 => n4014
                           , ZN => DataP_PC_reg_N26);
   U2569 : INV_X1 port map( A => DataP_npc_24_port, ZN => n4014);
   U2570 : AOI21_X1 port map( B1 => n3563, B2 => n3691, A => n3562, ZN => n308)
                           ;
   U2571 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N42, A2 => n3007, ZN =>
                           n3559);
   U2572 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N74, B2 => n3703, A => 
                           n3558, ZN => n3560);
   U2573 : OAI211_X1 port map( C1 => n3909, C2 => n3700, A => n3557, B => n3556
                           , ZN => n3558);
   U2574 : NAND2_X1 port map( A1 => DataP_alu_a_in_24_port, A2 => n3697, ZN => 
                           n3556);
   U2575 : OAI211_X1 port map( C1 => DataP_alu_a_in_24_port, C2 => n3697, A => 
                           DataP_alu_b_in_24_port, B => n3660, ZN => n3557);
   U2576 : XNOR2_X1 port map( A => DataP_alu_a_in_24_port, B => 
                           DataP_alu_b_in_24_port, ZN => n3909);
   U2577 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N106, A2 => n3675, ZN 
                           => n3561);
   U2578 : INV_X1 port map( A => n2919, ZN => n2983);
   U2579 : XNOR2_X1 port map( A => n2423, B => n2158, ZN => n3563);
   U2580 : OAI22_X1 port map( A1 => n323, A2 => n3911, B1 => n3910, B2 => n4007
                           , ZN => DataP_PC_reg_N19);
   U2581 : INV_X1 port map( A => DataP_npc_17_port, ZN => n4007);
   U2582 : AOI21_X1 port map( B1 => n3621, B2 => n3691, A => n3620, ZN => n323)
                           ;
   U2583 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N67, B2 => n3703, A => 
                           n3616, ZN => n3618);
   U2584 : OAI211_X1 port map( C1 => n3615, C2 => n3700, A => n3614, B => n3613
                           , ZN => n3616);
   U2585 : OAI211_X1 port map( C1 => DataP_alu_a_in_17_port, C2 => n3697, A => 
                           DataP_alu_b_in_17_port, B => n3660, ZN => n3613);
   U2586 : NAND2_X1 port map( A1 => DataP_alu_a_in_17_port, A2 => n3697, ZN => 
                           n3614);
   U2587 : XNOR2_X1 port map( A => DataP_alu_a_in_17_port, B => 
                           DataP_alu_b_in_17_port, ZN => n3615);
   U2588 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N99, A2 => n3675, ZN =>
                           n3619);
   U2589 : OAI22_X1 port map( A1 => n303, A2 => n3911, B1 => n3910, B2 => n4016
                           , ZN => DataP_PC_reg_N28);
   U2590 : INV_X1 port map( A => DataP_npc_26_port, ZN => n4016);
   U2591 : AOI21_X1 port map( B1 => n3542, B2 => n3691, A => n3541, ZN => n303)
                           ;
   U2592 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N76, B2 => n3703, A => 
                           n3537, ZN => n3539);
   U2593 : OAI211_X1 port map( C1 => n3536, C2 => n3700, A => n3535, B => n3534
                           , ZN => n3537);
   U2594 : NAND2_X1 port map( A1 => DataP_alu_a_in_26_port, A2 => n3697, ZN => 
                           n3534);
   U2595 : OAI211_X1 port map( C1 => DataP_alu_a_in_26_port, C2 => n3697, A => 
                           DataP_alu_b_in_26_port, B => n3660, ZN => n3535);
   U2596 : XNOR2_X1 port map( A => DataP_alu_a_in_26_port, B => 
                           DataP_alu_b_in_26_port, ZN => n3536);
   U2597 : XNOR2_X1 port map( A => n1590, B => n3533, ZN => n3542);
   U2598 : INV_X1 port map( A => n3472, ZN => n2421);
   U2599 : OAI21_X1 port map( B1 => n3544, B2 => n3555, A => n3543, ZN => n3472
                           );
   U2600 : INV_X1 port map( A => n3502, ZN => n3555);
   U2601 : INV_X1 port map( A => n3497, ZN => n3465);
   U2602 : INV_X1 port map( A => DataP_npc_28_port, ZN => n4018);
   U2603 : OAI211_X1 port map( C1 => n3695, C2 => n2928, A => n3530, B => n3529
                           , ZN => n3531);
   U2604 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N78, B2 => n3703, A => 
                           n3528, ZN => n3529);
   U2605 : OAI21_X1 port map( B1 => n3700, B2 => n3527, A => n3526, ZN => n3528
                           );
   U2606 : AOI22_X1 port map( A1 => n3525, A2 => DataP_alu_b_in_28_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_28_port, ZN => n3526);
   U2607 : OAI21_X1 port map( B1 => n1811, B2 => n3671, A => n3694, ZN => n3525
                           );
   U2608 : XNOR2_X1 port map( A => DataP_alu_a_in_28_port, B => 
                           DataP_alu_b_in_28_port, ZN => n3527);
   U2609 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N46, A2 => n3007, ZN =>
                           n3530);
   U2610 : XNOR2_X1 port map( A => n3523, B => n1811, ZN => n3524);
   U2611 : INV_X1 port map( A => DataP_npc_23_port, ZN => n4013);
   U2612 : AOI21_X1 port map( B1 => n3455, B2 => n3691, A => n3454, ZN => n309)
                           ;
   U2613 : OAI211_X1 port map( C1 => n3453, C2 => n3695, A => n3452, B => n3451
                           , ZN => n3454);
   U2614 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N73, B2 => n3703, A => 
                           n3450, ZN => n3452);
   U2615 : OAI211_X1 port map( C1 => n3908, C2 => n3700, A => n3449, B => n3448
                           , ZN => n3450);
   U2616 : NAND2_X1 port map( A1 => DataP_alu_a_in_23_port, A2 => n3697, ZN => 
                           n3448);
   U2617 : OAI211_X1 port map( C1 => DataP_alu_a_in_23_port, C2 => n3697, A => 
                           DataP_alu_b_in_23_port, B => n3660, ZN => n3449);
   U2618 : XNOR2_X1 port map( A => DataP_alu_a_in_23_port, B => 
                           DataP_alu_b_in_23_port, ZN => n3908);
   U2619 : INV_X1 port map( A => DataP_ALU_C_shifter_N105, ZN => n3453);
   U2620 : INV_X1 port map( A => n2917, ZN => n2982);
   U2621 : AND2_X1 port map( A1 => n2527, A2 => n2524, ZN => n2523);
   U2622 : NAND2_X1 port map( A1 => n2526, A2 => n2525, ZN => n2524);
   U2623 : NOR2_X1 port map( A1 => n3456, A2 => n1893, ZN => n2525);
   U2624 : AND2_X1 port map( A1 => n1998, A2 => n1610, ZN => n2527);
   U2625 : AND3_X1 port map( A1 => n1559, A2 => n1557, A3 => n1959, ZN => n2526
                           );
   U2626 : INV_X1 port map( A => DataP_npc_31_port, ZN => n4023);
   U2627 : OAI22_X1 port map( A1 => n319, A2 => n3911, B1 => n3910, B2 => n4009
                           , ZN => DataP_PC_reg_N21);
   U2628 : INV_X1 port map( A => DataP_npc_19_port, ZN => n4009);
   U2629 : AOI21_X1 port map( B1 => n3436, B2 => n3691, A => n3435, ZN => n319)
                           ;
   U2630 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N37, A2 => n3007, ZN =>
                           n3432);
   U2631 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N69, B2 => n3006, A => 
                           n3431, ZN => n3433);
   U2632 : OAI211_X1 port map( C1 => n3906, C2 => n3700, A => n3430, B => n3429
                           , ZN => n3431);
   U2633 : NAND2_X1 port map( A1 => n1553, A2 => n3697, ZN => n3429);
   U2634 : OAI211_X1 port map( C1 => n1553, C2 => n3697, A => 
                           DataP_alu_b_in_19_port, B => n3660, ZN => n3430);
   U2635 : XNOR2_X1 port map( A => n1553, B => DataP_alu_b_in_19_port, ZN => 
                           n3906);
   U2636 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N101, A2 => n3675, ZN 
                           => n3434);
   U2637 : AOI21_X1 port map( B1 => n2226, B2 => n1919, A => n2223, ZN => n2411
                           );
   U2638 : INV_X1 port map( A => DataP_npc_30_port, ZN => n4020);
   U2639 : NOR2_X1 port map( A1 => n3674, A2 => n3911, ZN => n2412);
   U2640 : OAI22_X1 port map( A1 => n322, A2 => n3911, B1 => n3910, B2 => n4008
                           , ZN => DataP_PC_reg_N20);
   U2641 : INV_X1 port map( A => DataP_npc_18_port, ZN => n4008);
   U2642 : INV_X1 port map( A => n3610, ZN => n322);
   U2643 : OAI211_X1 port map( C1 => n3609, C2 => n3674, A => n3608, B => n3607
                           , ZN => n3610);
   U2644 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N100, A2 => n3675, ZN 
                           => n3607);
   U2645 : AOI21_X1 port map( B1 => n3007, B2 => DataP_ALU_C_shifter_N36, A => 
                           n3606, ZN => n3608);
   U2646 : OAI211_X1 port map( C1 => n3700, C2 => n3605, A => n3604, B => n3603
                           , ZN => n3606);
   U2647 : AOI22_X1 port map( A1 => n3602, A2 => DataP_alu_b_in_18_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_18_port, ZN => n3603);
   U2648 : OAI21_X1 port map( B1 => n1884, B2 => n3671, A => n3694, ZN => n3602
                           );
   U2649 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N68, A2 => n3006, ZN =>
                           n3604);
   U2650 : XNOR2_X1 port map( A => DataP_alu_a_in_18_port, B => 
                           DataP_alu_b_in_18_port, ZN => n3605);
   U2651 : INV_X1 port map( A => n3441, ZN => n3423);
   U2652 : OAI22_X1 port map( A1 => n332, A2 => n3911, B1 => n3910, B2 => n4004
                           , ZN => DataP_PC_reg_N16);
   U2653 : INV_X1 port map( A => DataP_npc_14_port, ZN => n4004);
   U2654 : INV_X1 port map( A => n3638, ZN => n332);
   U2655 : OAI211_X1 port map( C1 => n3637, C2 => n3674, A => n3636, B => n3635
                           , ZN => n3638);
   U2656 : AOI22_X1 port map( A1 => DataP_ALU_C_shifter_N32, A2 => n3706, B1 =>
                           n3675, B2 => DataP_ALU_C_shifter_N96, ZN => n3635);
   U2657 : INV_X1 port map( A => n2680, ZN => n2701);
   U2658 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N64, B2 => n3006, A => 
                           n3634, ZN => n3636);
   U2659 : XNOR2_X1 port map( A => DataP_alu_a_in_14_port, B => n1932, ZN => 
                           n3633);
   U2660 : XNOR2_X1 port map( A => n3632, B => n3631, ZN => n3637);
   U2661 : OAI21_X1 port map( B1 => n2939, B2 => n3695, A => n3486, ZN => n3512
                           );
   U2662 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N80, B2 => n3006, A => 
                           n3485, ZN => n3486);
   U2663 : OAI211_X1 port map( C1 => n3484, C2 => n3700, A => n3483, B => n3482
                           , ZN => n3485);
   U2664 : NAND2_X1 port map( A1 => DataP_alu_a_in_30_port, A2 => n3697, ZN => 
                           n3482);
   U2665 : OAI211_X1 port map( C1 => DataP_alu_a_in_30_port, C2 => n3697, A => 
                           DataP_alu_b_in_30_port, B => n3660, ZN => n3483);
   U2666 : XNOR2_X1 port map( A => DataP_alu_a_in_30_port, B => 
                           DataP_alu_b_in_30_port, ZN => n3484);
   U2667 : NAND2_X1 port map( A1 => n3705, A2 => n3683, ZN => n3511);
   U2668 : OAI22_X1 port map( A1 => n330, A2 => n3911, B1 => n3910, B2 => n4005
                           , ZN => DataP_PC_reg_N17);
   U2669 : INV_X1 port map( A => DataP_npc_15_port, ZN => n4005);
   U2670 : AOI21_X1 port map( B1 => n2385, B2 => n3691, A => n2384, ZN => n330)
                           ;
   U2671 : NAND2_X1 port map( A1 => n3406, A2 => n3407, ZN => n2384);
   U2672 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N65, B2 => n3006, A => 
                           n3405, ZN => n3407);
   U2673 : OAI211_X1 port map( C1 => n1842, C2 => n3694, A => n3404, B => n3403
                           , ZN => n3405);
   U2674 : NAND2_X1 port map( A1 => n3694, A2 => n3671, ZN => n3660);
   U2675 : NAND2_X1 port map( A1 => n3402, A2 => n1939, ZN => n3404);
   U2676 : AOI22_X1 port map( A1 => DataP_ALU_C_shifter_N33, A2 => n3706, B1 =>
                           n3675, B2 => DataP_ALU_C_shifter_N97, ZN => n3406);
   U2677 : INV_X1 port map( A => n2688, ZN => n2702);
   U2678 : XNOR2_X1 port map( A => n2386, B => n3413, ZN => n2385);
   U2679 : OAI21_X1 port map( B1 => n3632, B2 => n3414, A => n3410, ZN => n2386
                           );
   U2680 : AOI21_X1 port map( B1 => n3399, B2 => n3409, A => n3644, ZN => n3632
                           );
   U2681 : INV_X1 port map( A => n3408, ZN => n3644);
   U2682 : OAI21_X1 port map( B1 => n3641, B2 => n3394, A => n3640, ZN => n3399
                           );
   U2683 : OAI21_X1 port map( B1 => n3264, B2 => n2481, A => n1529, ZN => n3640
                           );
   U2684 : INV_X1 port map( A => n3642, ZN => n3394);
   U2685 : NAND2_X1 port map( A1 => n2288, A2 => n2294, ZN => n3642);
   U2686 : NAND2_X1 port map( A1 => n3264, A2 => n3510, ZN => n2288);
   U2687 : INV_X1 port map( A => DataP_npc_29_port, ZN => n4019);
   U2688 : INV_X1 port map( A => n3711, ZN => n3229);
   U2689 : OAI211_X1 port map( C1 => n3695, C2 => n2930, A => n3521, B => n3520
                           , ZN => n3522);
   U2690 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N79, B2 => n3703, A => 
                           n3519, ZN => n3520);
   U2691 : OAI21_X1 port map( B1 => n3700, B2 => n3518, A => n3517, ZN => n3519
                           );
   U2692 : AOI22_X1 port map( A1 => n3516, A2 => DataP_alu_b_in_29_port, B1 => 
                           n3697, B2 => DataP_alu_a_in_29_port, ZN => n3517);
   U2693 : OAI21_X1 port map( B1 => n1925, B2 => n3671, A => n3694, ZN => n3516
                           );
   U2694 : XNOR2_X1 port map( A => DataP_alu_a_in_29_port, B => 
                           DataP_alu_b_in_29_port, ZN => n3518);
   U2695 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N47, A2 => n3007, ZN =>
                           n3521);
   U2696 : INV_X1 port map( A => n2514, ZN => n3514);
   U2697 : INV_X1 port map( A => n3513, ZN => n3515);
   U2698 : OAI21_X1 port map( B1 => n2371, B2 => n2321, A => n2280, ZN => n3513
                           );
   U2699 : INV_X1 port map( A => n2515, ZN => n2426);
   U2700 : AND2_X1 port map( A1 => n2550, A2 => n2147, ZN => n2430);
   U2701 : AOI21_X1 port map( B1 => n2417, B2 => n2416, A => n2414, ZN => n3707
                           );
   U2702 : NAND2_X1 port map( A1 => n2415, A2 => n3704, ZN => n2414);
   U2703 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N81, B2 => n3006, A => 
                           n3702, ZN => n3704);
   U2704 : OAI21_X1 port map( B1 => n3701, B2 => n3700, A => n3699, ZN => n3702
                           );
   U2705 : AOI22_X1 port map( A1 => DataP_alu_a_in_31_port, A2 => n3698, B1 => 
                           n3697, B2 => DataP_alu_b_in_31_port, ZN => n3699);
   U2706 : NAND2_X1 port map( A1 => n3226, A2 => n3343, ZN => n3694);
   U2707 : INV_X1 port map( A => n3903, ZN => n3222);
   U2708 : NAND2_X1 port map( A1 => DataP_alu_b_in_31_port, A2 => n3693, ZN => 
                           n3696);
   U2709 : INV_X1 port map( A => n3671, ZN => n3693);
   U2710 : OR2_X1 port map( A1 => n3225, A2 => n3345, ZN => n3671);
   U2711 : INV_X1 port map( A => n3224, ZN => n3225);
   U2712 : NOR2_X1 port map( A1 => n3015, A2 => ALU_OPCODE_i_1_port, ZN => 
                           n3226);
   U2713 : NAND2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => n443, ZN => 
                           n3015);
   U2714 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N49, A2 => n3007, ZN =>
                           n2415);
   U2715 : INV_X1 port map( A => n3343, ZN => n3221);
   U2716 : NOR2_X1 port map( A1 => n3692, A2 => n3674, ZN => n2416);
   U2717 : INV_X1 port map( A => n3705, ZN => n2417);
   U2718 : XNOR2_X1 port map( A => ALU_OPCODE_i_2_port, B => n3902, ZN => n3199
                           );
   U2719 : NAND2_X1 port map( A1 => n3197, A2 => n3348, ZN => n3201);
   U2720 : NOR2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => 
                           ALU_OPCODE_i_1_port, ZN => n3348);
   U2721 : OAI21_X1 port map( B1 => n443, B2 => ALU_OPCODE_i_3_port, A => n3345
                           , ZN => n3197);
   U2722 : NAND2_X1 port map( A1 => n3493, A2 => n1924, ZN => n3705);
   U2723 : INV_X1 port map( A => n3687, ZN => n3701);
   U2724 : XNOR2_X1 port map( A => n3688, B => n3687, ZN => n3690);
   U2725 : XNOR2_X1 port map( A => DataP_alu_a_in_31_port, B => n1935, ZN => 
                           n3687);
   U2726 : NOR2_X1 port map( A1 => n2562, A2 => n2191, ZN => n3130);
   U2727 : OAI21_X1 port map( B1 => n1837, B2 => n1, A => n3129, ZN => n3131);
   U2728 : OR2_X1 port map( A1 => n3686, A2 => DataP_alu_b_in_30_port, ZN => 
                           n3688);
   U2729 : INV_X1 port map( A => n3683, ZN => n3684);
   U2730 : NOR2_X1 port map( A1 => n2563, A2 => n2192, ZN => n3133);
   U2731 : OAI21_X1 port map( B1 => n2999, B2 => n5, A => n3132, ZN => n3134);
   U2732 : XNOR2_X1 port map( A => n3686, B => DataP_alu_b_in_30_port, ZN => 
                           n3491);
   U2733 : NAND2_X1 port map( A1 => n3490, A2 => n3489, ZN => n3686);
   U2734 : NOR2_X1 port map( A1 => DataP_alu_b_in_29_port, A2 => 
                           DataP_alu_b_in_28_port, ZN => n3489);
   U2735 : INV_X1 port map( A => DataP_alu_b_in_30_port, ZN => n3492);
   U2736 : AND2_X1 port map( A1 => n2429, A2 => n2513, ZN => n2427);
   U2737 : NAND2_X1 port map( A1 => n2515, A2 => n2514, ZN => n2429);
   U2738 : NAND2_X1 port map( A1 => n2278, A2 => n2279, ZN => n2514);
   U2739 : NAND2_X1 port map( A1 => n2371, A2 => n2407, ZN => n2278);
   U2740 : AND2_X1 port map( A1 => n2513, A2 => n2147, ZN => n2428);
   U2741 : NOR2_X1 port map( A1 => n2563, A2 => n2206, ZN => n3139);
   U2742 : OAI21_X1 port map( B1 => n2999, B2 => n13, A => n3138, ZN => n3140);
   U2743 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_28_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_28_port, ZN => n3138);
   U2744 : NOR2_X1 port map( A1 => n1925, A2 => n2281, ZN => n2280);
   U2745 : NOR2_X1 port map( A1 => n2561, A2 => n2199, ZN => n3136);
   U2746 : OAI21_X1 port map( B1 => n2999, B2 => n9, A => n3135, ZN => n3137);
   U2747 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_29_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_29_port, ZN => n3135);
   U2748 : NAND4_X1 port map( A1 => n3306, A2 => n3294, A3 => n3293, A4 => 
                           n3292, ZN => DataP_alu_b_in_28_port);
   U2749 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_28_port, ZN =>
                           n3292);
   U2750 : OR2_X1 port map( A1 => n1636, A2 => n2178, ZN => n3293);
   U2751 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_28_port, ZN => n3294
                           );
   U2752 : NOR2_X1 port map( A1 => n3487, A2 => DataP_alu_b_in_27_port, ZN => 
                           n3509);
   U2753 : NAND2_X1 port map( A1 => n3507, A2 => DataP_alu_a_in_27_port, ZN => 
                           n3508);
   U2754 : NAND2_X1 port map( A1 => n2474, A2 => n2473, ZN => n3507);
   U2755 : INV_X1 port map( A => n1548, ZN => n2554);
   U2756 : NOR2_X1 port map( A1 => n2563, A2 => n2193, ZN => n3142);
   U2757 : OAI21_X1 port map( B1 => n1837, B2 => n17, A => n3141, ZN => n3143);
   U2758 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_27_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_27_port, ZN => n3141);
   U2759 : INV_X1 port map( A => n3487, ZN => n2497);
   U2760 : NAND2_X1 port map( A1 => n2241, A2 => n1936, ZN => n3487);
   U2761 : NAND4_X1 port map( A1 => n3306, A2 => n3297, A3 => n3296, A4 => 
                           n3295, ZN => DataP_alu_b_in_27_port);
   U2762 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_27_port, ZN =>
                           n3295);
   U2763 : OR2_X1 port map( A1 => n2566, A2 => n2165, ZN => n3296);
   U2764 : NAND2_X1 port map( A1 => n1859, A2 => DataP_B_s_27_port, ZN => n3297
                           );
   U2765 : OR2_X1 port map( A1 => n3532, A2 => n2556, ZN => n2555);
   U2766 : NOR2_X1 port map( A1 => n2563, A2 => n2207, ZN => n3148);
   U2767 : OAI21_X1 port map( B1 => n2999, B2 => n25, A => n3147, ZN => n3149);
   U2768 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_25_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_25_port, ZN => n3147);
   U2769 : NOR2_X1 port map( A1 => n2563, A2 => n2200, ZN => n3145);
   U2770 : OAI21_X1 port map( B1 => n3000, B2 => n21, A => n3144, ZN => n3146);
   U2771 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_26_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_26_port, ZN => n3144);
   U2772 : NAND2_X1 port map( A1 => DataP_alu_b_in_26_port, A2 => n1938, ZN => 
                           n2502);
   U2773 : INV_X1 port map( A => DataP_alu_b_in_25_port, ZN => n3473);
   U2774 : NAND2_X1 port map( A1 => n2565, A2 => DataP_IMM_s_31_port, ZN => 
                           n3306);
   U2775 : NAND2_X1 port map( A1 => n3471, A2 => DataP_alu_a_in_24_port, ZN => 
                           n3502);
   U2776 : AND2_X1 port map( A1 => n3497, A2 => n3496, ZN => n2353);
   U2777 : NAND2_X1 port map( A1 => n3496, A2 => n3463, ZN => n3564);
   U2778 : NAND2_X1 port map( A1 => n3447, A2 => n3566, ZN => n3463);
   U2779 : INV_X1 port map( A => DataP_alu_a_in_22_port, ZN => n3566);
   U2780 : AND2_X1 port map( A1 => n3459, A2 => n1533, ZN => n2352);
   U2781 : AND2_X1 port map( A1 => n3578, A2 => n3580, ZN => n3593);
   U2782 : AOI21_X1 port map( B1 => n3495, B2 => n3497, A => n3554, ZN => n3500
                           );
   U2783 : NOR2_X1 port map( A1 => n3471, A2 => DataP_alu_a_in_24_port, ZN => 
                           n3554);
   U2784 : NOR2_X1 port map( A1 => n1539, A2 => n2217, ZN => n3151);
   U2785 : OAI21_X1 port map( B1 => n3000, B2 => n29, A => n3150, ZN => n3152);
   U2786 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_24_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_24_port, ZN => n3150);
   U2787 : XNOR2_X1 port map( A => n3488, B => DataP_alu_b_in_24_port, ZN => 
                           n3469);
   U2788 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_24_port, ZN =>
                           n3319);
   U2789 : OR2_X1 port map( A1 => n1636, A2 => n2179, ZN => n3320);
   U2790 : NAND2_X1 port map( A1 => n1905, A2 => DataP_IMM_s_24_port, ZN => 
                           n3321);
   U2791 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_24_port, ZN => n3322
                           );
   U2792 : XNOR2_X1 port map( A => n3464, B => DataP_alu_a_in_23_port, ZN => 
                           n3495);
   U2793 : NOR2_X1 port map( A1 => n1539, A2 => n2194, ZN => n3154);
   U2794 : OAI21_X1 port map( B1 => n1837, B2 => n33, A => n3153, ZN => n3155);
   U2795 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_23_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_23_port, ZN => n3153);
   U2796 : XNOR2_X1 port map( A => n3439, B => n1937, ZN => n3440);
   U2797 : INV_X1 port map( A => n3444, ZN => n3468);
   U2798 : INV_X1 port map( A => n2382, ZN => n2380);
   U2799 : NAND2_X1 port map( A1 => n1560, A2 => n3576, ZN => n3443);
   U2800 : AND2_X1 port map( A1 => n2382, A2 => DataP_alu_a_in_21_port, ZN => 
                           n2370);
   U2801 : NOR2_X1 port map( A1 => n2563, A2 => n2201, ZN => n3160);
   U2802 : OAI21_X1 port map( B1 => n2999, B2 => n41, A => n3159, ZN => n3161);
   U2803 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_21_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_21_port, ZN => n3159);
   U2804 : NAND2_X1 port map( A1 => n2007, A2 => DataP_alu_a_in_20_port, ZN => 
                           n3578);
   U2805 : NOR2_X1 port map( A1 => n2561, A2 => n2208, ZN => n3163);
   U2806 : OAI21_X1 port map( B1 => n2999, B2 => n45, A => n3162, ZN => n3164);
   U2807 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_20_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_20_port, ZN => n3162);
   U2808 : AND3_X1 port map( A1 => n3496, A2 => n1610, A3 => n3456, ZN => n3457
                           );
   U2809 : NOR2_X1 port map( A1 => n2561, A2 => n2218, ZN => n3157);
   U2810 : OAI21_X1 port map( B1 => n2999, B2 => n37, A => n3156, ZN => n3158);
   U2811 : AOI22_X1 port map( A1 => n2995, A2 => DataP_alu_out_M_22_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_22_port, ZN => n3156);
   U2812 : NAND4_X1 port map( A1 => n3326, A2 => n3325, A3 => n3324, A4 => 
                           n3323, ZN => DataP_alu_b_in_22_port);
   U2813 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_22_port, ZN =>
                           n3323);
   U2814 : OR2_X1 port map( A1 => n3002, A2 => n2180, ZN => n3324);
   U2815 : NAND2_X1 port map( A1 => n1848, A2 => DataP_IMM_s_22_port, ZN => 
                           n3325);
   U2816 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_22_port, ZN => n3326
                           );
   U2817 : NAND2_X1 port map( A1 => n3442, A2 => n1556, ZN => n3444);
   U2818 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_20_port, ZN =>
                           n3285);
   U2819 : OR2_X1 port map( A1 => n1636, A2 => n2173, ZN => n3286);
   U2820 : NAND2_X1 port map( A1 => n1905, A2 => DataP_IMM_s_20_port, ZN => 
                           n3287);
   U2821 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_20_port, ZN => n3288
                           );
   U2822 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_21_port, ZN =>
                           n3331);
   U2823 : OR2_X1 port map( A1 => n3002, A2 => n2172, ZN => n3332);
   U2824 : NAND2_X1 port map( A1 => n1848, A2 => DataP_IMM_s_21_port, ZN => 
                           n3333);
   U2825 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_21_port, ZN => n3334
                           );
   U2826 : OAI211_X1 port map( C1 => n3441, C2 => n1531, A => n1877, B => n1557
                           , ZN => n3462);
   U2827 : NOR2_X1 port map( A1 => n2561, A2 => n2202, ZN => n3166);
   U2828 : OAI21_X1 port map( B1 => n3000, B2 => n49, A => n3165, ZN => n3167);
   U2829 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_19_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_19_port, ZN => n3165);
   U2830 : NAND2_X1 port map( A1 => n2306, A2 => n3291, ZN => 
                           DataP_alu_b_in_19_port);
   U2831 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_19_port, ZN => n3291
                           );
   U2832 : NAND2_X1 port map( A1 => n3289, A2 => n3290, ZN => n2307);
   U2833 : OR2_X1 port map( A1 => n3002, A2 => n2174, ZN => n3289);
   U2834 : NOR2_X1 port map( A1 => n1539, A2 => n2209, ZN => n3169);
   U2835 : OAI21_X1 port map( B1 => n2999, B2 => n53, A => n3168, ZN => n3170);
   U2836 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_18_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_18_port, ZN => n3168);
   U2837 : NAND2_X1 port map( A1 => n3001, A2 => DataP_B_s_18_port, ZN => n3281
                           );
   U2838 : INV_X1 port map( A => n2245, ZN => n2439);
   U2839 : AOI21_X1 port map( B1 => n2354, B2 => n3611, A => n2308, ZN => n3441
                           );
   U2840 : OAI211_X1 port map( C1 => n2494, C2 => n2492, A => n2489, B => n2491
                           , ZN => n2299);
   U2841 : OR2_X1 port map( A1 => n3437, A2 => n2490, ZN => n2489);
   U2842 : NAND2_X1 port map( A1 => n2538, A2 => n3424, ZN => n2490);
   U2843 : INV_X1 port map( A => n2538, ZN => n2492);
   U2844 : OAI21_X1 port map( B1 => n3422, B2 => n2383, A => n2465, ZN => n3611
                           );
   U2845 : NOR2_X1 port map( A1 => n2563, A2 => n2219, ZN => n3174);
   U2846 : OAI21_X1 port map( B1 => n2999, B2 => n61, A => n3173, ZN => n3175);
   U2847 : AOI22_X1 port map( A1 => n2997, A2 => DataP_alu_out_M_16_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_16_port, ZN => n3173);
   U2848 : XNOR2_X1 port map( A => n1563, B => DataP_alu_b_in_16_port, ZN => 
                           n3422);
   U2849 : NOR2_X1 port map( A1 => n1539, A2 => n2195, ZN => n3171);
   U2850 : NAND3_X1 port map( A1 => n2488, A2 => n2494, A3 => n2463, ZN => 
                           n2462);
   U2851 : NAND2_X1 port map( A1 => n1848, A2 => DataP_IMM_s_16_port, ZN => 
                           n3314);
   U2852 : OR2_X1 port map( A1 => n3002, A2 => n2167, ZN => n3313);
   U2853 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_16_port, ZN =>
                           n2520);
   U2854 : NAND2_X1 port map( A1 => n1839, A2 => DataP_B_s_16_port, ZN => n3315
                           );
   U2855 : NAND2_X1 port map( A1 => n1905, A2 => DataP_IMM_s_17_port, ZN => 
                           n3304);
   U2856 : OR2_X1 port map( A1 => n2566, A2 => n2170, ZN => n3303);
   U2857 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_17_port, ZN =>
                           n2519);
   U2858 : NAND2_X1 port map( A1 => n1839, A2 => DataP_B_s_17_port, ZN => n3305
                           );
   U2859 : AND2_X1 port map( A1 => n3417, A2 => n3418, ZN => n2390);
   U2860 : INV_X1 port map( A => n3413, ZN => n2541);
   U2861 : XNOR2_X1 port map( A => DataP_alu_a_in_15_port, B => n3417, ZN => 
                           n3402);
   U2862 : NAND2_X1 port map( A1 => n3392, A2 => n1842, ZN => n3391);
   U2863 : NOR2_X1 port map( A1 => n2561, A2 => n2196, ZN => n3177);
   U2864 : OAI21_X1 port map( B1 => n3000, B2 => n65, A => n3176, ZN => n3178);
   U2865 : AOI22_X1 port map( A1 => n2997, A2 => DataP_alu_out_M_15_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_15_port, ZN => n3176);
   U2866 : INV_X1 port map( A => n1881, ZN => n2482);
   U2867 : INV_X1 port map( A => n3417, ZN => DataP_alu_b_in_15_port);
   U2868 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_15_port, ZN => 
                           n3302);
   U2869 : NAND2_X1 port map( A1 => n3004, A2 => DataP_alu_out_W_15_port, ZN =>
                           n3300);
   U2870 : OR2_X1 port map( A1 => n3002, A2 => n2166, ZN => n3301);
   U2871 : NOR2_X1 port map( A1 => n1881, A2 => n1932, ZN => n2487);
   U2872 : AND2_X1 port map( A1 => n3411, A2 => n3410, ZN => n3631);
   U2873 : INV_X1 port map( A => n3510, ZN => n2543);
   U2874 : NAND2_X1 port map( A1 => n3398, A2 => n1927, ZN => n3408);
   U2875 : AOI21_X1 port map( B1 => n3397, B2 => n3510, A => n2546, ZN => n3398
                           );
   U2876 : INV_X1 port map( A => n3411, ZN => n3414);
   U2877 : NAND2_X1 port map( A1 => n3401, A2 => DataP_alu_a_in_14_port, ZN => 
                           n3411);
   U2878 : NOR2_X1 port map( A1 => n1539, A2 => n2203, ZN => n3180);
   U2879 : OAI21_X1 port map( B1 => n3000, B2 => n69, A => n3179, ZN => n3181);
   U2880 : AOI22_X1 port map( A1 => n2997, A2 => DataP_alu_out_M_14_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_14_port, ZN => n3179);
   U2881 : OAI21_X1 port map( B1 => n2375, B2 => n2376, A => n2373, ZN => n2372
                           );
   U2882 : NAND2_X1 port map( A1 => n1881, A2 => n2374, ZN => n2373);
   U2883 : NOR2_X1 port map( A1 => n1932, A2 => n2375, ZN => n2374);
   U2884 : NAND2_X1 port map( A1 => n2482, A2 => n1932, ZN => n2376);
   U2885 : INV_X1 port map( A => n3510, ZN => n2375);
   U2886 : OR2_X1 port map( A1 => n3002, A2 => n2171, ZN => n3312);
   U2887 : NAND2_X1 port map( A1 => n3004, A2 => DataP_alu_out_W_14_port, ZN =>
                           n3311);
   U2888 : INV_X1 port map( A => n3409, ZN => n3645);
   U2889 : OAI21_X1 port map( B1 => n2546, B2 => n3397, A => n2149, ZN => n3409
                           );
   U2890 : NAND2_X1 port map( A1 => n2548, A2 => n2545, ZN => n2544);
   U2891 : INV_X1 port map( A => n3510, ZN => n2545);
   U2892 : NOR2_X1 port map( A1 => n1539, A2 => n2210, ZN => n3183);
   U2893 : OAI21_X1 port map( B1 => n3000, B2 => n73, A => n3182, ZN => n3184);
   U2894 : AOI22_X1 port map( A1 => n2997, A2 => DataP_alu_out_M_13_port, B1 =>
                           n2991, B2 => DataP_alu_out_W_13_port, ZN => n3182);
   U2895 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_13_port, ZN =>
                           n3307);
   U2896 : OR2_X1 port map( A1 => n2566, A2 => n2176, ZN => n3308);
   U2897 : NAND2_X1 port map( A1 => n1848, A2 => DataP_ir_E_13_port, ZN => 
                           n3309);
   U2898 : NAND2_X1 port map( A1 => n1839, A2 => DataP_B_s_13_port, ZN => n3310
                           );
   U2899 : AND2_X1 port map( A1 => n1903, A2 => n2442, ZN => n2504);
   U2900 : NAND2_X1 port map( A1 => n2294, A2 => n1938, ZN => n2289);
   U2901 : NOR2_X1 port map( A1 => n2561, A2 => n2197, ZN => n3186);
   U2902 : OAI21_X1 port map( B1 => n3000, B2 => n77, A => n3185, ZN => n3187);
   U2903 : AOI22_X1 port map( A1 => n2997, A2 => DataP_alu_out_M_12_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_12_port, ZN => n3185);
   U2904 : NAND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_12_port, ZN =>
                           n3261);
   U2905 : AND2_X1 port map( A1 => n1889, A2 => n2142, ZN => n3400);
   U2906 : INV_X1 port map( A => DataP_alu_a_in_10_port, ZN => n3236);
   U2907 : NAND2_X1 port map( A1 => n3232, A2 => n3656, ZN => n3267);
   U2908 : NAND2_X1 port map( A1 => n3658, A2 => n1921, ZN => n3656);
   U2909 : NAND2_X1 port map( A1 => n3220, A2 => n1922, ZN => n3232);
   U2910 : INV_X1 port map( A => n1572, ZN => n3254);
   U2911 : NOR2_X1 port map( A1 => n2561, A2 => n2204, ZN => n3189);
   U2912 : OAI21_X1 port map( B1 => n1837, B2 => n81, A => n3188, ZN => n3190);
   U2913 : AOI22_X1 port map( A1 => n2997, A2 => DRAM_ADDRESS_11_port, B1 => 
                           n2992, B2 => DataP_alu_out_W_11_port, ZN => n3188);
   U2914 : INV_X1 port map( A => n3251, ZN => n3250);
   U2915 : NAND2_X1 port map( A1 => n3004, A2 => DataP_alu_out_W_11_port, ZN =>
                           n3244);
   U2916 : OR2_X1 port map( A1 => n2566, A2 => n2164, ZN => n3245);
   U2917 : AND4_X1 port map( A1 => n3265, A2 => n2450, A3 => n3266, A4 => n3657
                           , ZN => n2319);
   U2918 : NOR2_X1 port map( A1 => n2999, A2 => n93, ZN => n3127);
   U2919 : OAI21_X1 port map( B1 => n2561, B2 => n2220, A => n3126, ZN => n3128
                           );
   U2920 : NAND2_X1 port map( A1 => n3215, A2 => n2508, ZN => n2509);
   U2921 : AND2_X1 port map( A1 => DataP_alu_b_in_8_port, A2 => n3510, ZN => 
                           n2508);
   U2922 : NAND2_X1 port map( A1 => n3219, A2 => DataP_alu_a_in_9_port, ZN => 
                           n3266);
   U2923 : NOR2_X1 port map( A1 => n2562, A2 => n2190, ZN => n3075);
   U2924 : OAI21_X1 port map( B1 => n1837, B2 => n89, A => n3074, ZN => n3076);
   U2925 : INV_X1 port map( A => n3220, ZN => n3219);
   U2926 : AND2_X1 port map( A1 => DataP_alu_b_in_9_port, A2 => n3510, ZN => 
                           n2329);
   U2927 : NAND2_X1 port map( A1 => n3218, A2 => n2545, ZN => n2549);
   U2928 : NOR2_X1 port map( A1 => n2561, A2 => n2211, ZN => n3195);
   U2929 : OAI21_X1 port map( B1 => n2999, B2 => n85, A => n3192, ZN => n3196);
   U2930 : AOI22_X1 port map( A1 => n2997, A2 => DRAM_ADDRESS_10_port, B1 => 
                           n2991, B2 => DataP_alu_out_W_10_port, ZN => n3192);
   U2931 : OR2_X1 port map( A1 => n1846, A2 => n2334, ZN => n2333);
   U2932 : INV_X1 port map( A => n2336, ZN => n2334);
   U2933 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_9_port, ZN => n2391
                           );
   U2934 : NOR2_X1 port map( A1 => n2561, A2 => n2205, ZN => n3078);
   U2935 : OAI21_X1 port map( B1 => n3000, B2 => n97, A => n3077, ZN => n3079);
   U2936 : XNOR2_X1 port map( A => n3208, B => DataP_alu_b_in_7_port, ZN => 
                           n3209);
   U2937 : INV_X1 port map( A => n3214, ZN => DataP_alu_b_in_7_port);
   U2938 : NAND2_X1 port map( A1 => n3207, A2 => n1611, ZN => n3208);
   U2939 : NAND2_X1 port map( A1 => n3666, A2 => n3384, ZN => n3211);
   U2940 : INV_X1 port map( A => DataP_alu_a_in_6_port, ZN => n3667);
   U2941 : NAND2_X1 port map( A1 => n3206, A2 => n1920, ZN => n3381);
   U2942 : INV_X1 port map( A => DataP_alu_a_in_4_port, ZN => n3204);
   U2943 : NAND2_X1 port map( A1 => n2420, A2 => DataP_alu_a_in_2_port, ZN => 
                           n3370);
   U2944 : OR2_X1 port map( A1 => n1996, A2 => n2337, ZN => n3359);
   U2945 : OAI21_X1 port map( B1 => n125, B2 => n3193, A => n3112, ZN => n3114)
                           ;
   U2946 : NOR2_X1 port map( A1 => n2560, A2 => n2214, ZN => n3113);
   U2947 : NOR2_X1 port map( A1 => n2561, A2 => n2215, ZN => n3116);
   U2948 : AND2_X1 port map( A1 => n3376, A2 => n3375, ZN => n3205);
   U2949 : NOR2_X1 port map( A1 => n2563, A2 => n2212, ZN => n3109);
   U2950 : OAI21_X1 port map( B1 => n1837, B2 => n113, A => n3108, ZN => n3110)
                           ;
   U2951 : NOR2_X1 port map( A1 => n2506, A2 => n2505, ZN => n3203);
   U2952 : NOR2_X1 port map( A1 => n1837, A2 => n109, ZN => n3118);
   U2953 : OAI21_X1 port map( B1 => n2562, B2 => n2221, A => n3117, ZN => n3119
                           );
   U2954 : NAND2_X1 port map( A1 => n1888, A2 => n3382, ZN => n3212);
   U2955 : NOR2_X1 port map( A1 => n2563, A2 => n2198, ZN => n3121);
   U2956 : OAI21_X1 port map( B1 => n3000, B2 => n105, A => n3120, ZN => n3122)
                           ;
   U2957 : NAND2_X1 port map( A1 => n3210, A2 => DataP_alu_a_in_6_port, ZN => 
                           n3384);
   U2958 : NOR2_X1 port map( A1 => n1539, A2 => n2216, ZN => n3124);
   U2959 : OAI21_X1 port map( B1 => n3000, B2 => n101, A => n3123, ZN => n3125)
                           ;
   U2960 : NOR2_X1 port map( A1 => n3031, A2 => n3682, ZN => n3068);
   U2961 : NAND4_X1 port map( A1 => n520, A2 => n149, A3 => n145, A4 => n147, 
                           ZN => n3682);
   U2962 : NAND2_X1 port map( A1 => n3710, A2 => n3061, ZN => n3067);
   U2963 : INV_X1 port map( A => n3073, ZN => n3061);
   U2964 : XNOR2_X1 port map( A => n1871, B => n2156, ZN => n3058);
   U2965 : XNOR2_X1 port map( A => n529, B => DataP_Rs1_1_port, ZN => n3054);
   U2966 : NOR2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => n2134, ZN => 
                           n3198);
   U2967 : XNOR2_X1 port map( A => n3207, B => n1611, ZN => n2522);
   U2968 : OR2_X1 port map( A1 => n3002, A2 => n2182, ZN => n2499);
   U2969 : AND2_X1 port map( A1 => n3045, A2 => n3044, ZN => n2314);
   U2970 : NOR2_X1 port map( A1 => n3043, A2 => n3042, ZN => n3044);
   U2971 : XNOR2_X1 port map( A => DataP_Rs2_3_port, B => n2570, ZN => n3043);
   U2972 : NOR2_X1 port map( A1 => n3041, A2 => n3040, ZN => n3045);
   U2973 : XNOR2_X1 port map( A => DataP_Rs2_1_port, B => n529, ZN => n3040);
   U2974 : OAI21_X1 port map( B1 => n3018, B2 => n2479, A => n2355, ZN => n3050
                           );
   U2975 : NAND4_X1 port map( A1 => n1546, A2 => n1532, A3 => 
                           DataP_opcode_W_4_port, A4 => n2159, ZN => n2355);
   U2976 : XNOR2_X1 port map( A => DataP_Rs2_2_port, B => DataP_add_D_2_port, 
                           ZN => n3020);
   U2977 : XNOR2_X1 port map( A => DataP_Rs2_4_port, B => DataP_add_D_4_port, 
                           ZN => n3027);
   U2978 : INV_X1 port map( A => DataP_alu_b_in_9_port, ZN => n3218);
   U2979 : INV_X1 port map( A => n1537, ZN => n2838);
   U2980 : AND3_X1 port map( A1 => n1867, A2 => n3691, A3 => n3505, ZN => n2138
                           );
   U2981 : AND2_X1 port map( A1 => n1948, A2 => n3689, ZN => n2139);
   U2982 : NAND2_X1 port map( A1 => n2181, A2 => n1995, ZN => n3215);
   U2983 : XOR2_X1 port map( A => DataP_dest_M_4_port, B => n540, Z => n2140);
   U2984 : NAND2_X1 port map( A1 => n3067, A2 => n3066, ZN => n3191);
   U2985 : INV_X1 port map( A => n2434, ZN => n2349);
   U2986 : AND2_X1 port map( A1 => n1897, A2 => n1898, ZN => n2142);
   U2987 : AND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_18_port, ZN => 
                           n2145);
   U2988 : INV_X1 port map( A => n1880, ZN => n3395);
   U2989 : OR2_X1 port map( A1 => n3523, A2 => n1811, ZN => n2147);
   U2990 : AND2_X1 port map( A1 => n3347, A2 => n2433, ZN => n2148);
   U2991 : AND2_X1 port map( A1 => DataP_alu_a_in_13_port, A2 => n2544, ZN => 
                           n2149);
   U2992 : INV_X1 port map( A => n2407, ZN => n2281);
   U2993 : INV_X1 port map( A => n2548, ZN => n2546);
   U2994 : INV_X1 port map( A => n3353, ZN => n3356);
   U2995 : OR2_X1 port map( A1 => n3555, A2 => n3554, ZN => n2158);
   U2996 : NAND2_X1 port map( A1 => n2146, A2 => ALU_OPCODE_i_0_port, ZN => 
                           n3345);
   U2997 : INV_X1 port map( A => n3345, ZN => n3223);
   U2998 : XOR2_X1 port map( A => DataP_add_D_1_port, B => n2160, Z => n2163);
   U2999 : INV_X1 port map( A => n3660, ZN => n3679);
   U3000 : AND2_X1 port map( A1 => n1603, A2 => n3214, ZN => n2181);
   U3001 : AND2_X1 port map( A1 => DataP_alu_b_in_19_port, A2 => n2545, ZN => 
                           n2183);
   U3002 : AND2_X1 port map( A1 => n3005, A2 => DataP_alu_out_W_19_port, ZN => 
                           n2184);
   U3003 : NAND2_X1 port map( A1 => n3474, A2 => DataP_alu_a_in_26_port, ZN => 
                           n3505);
   U3004 : AND2_X1 port map( A1 => n3580, A2 => n2011, ZN => n2188);
   U3005 : INV_X1 port map( A => n3191, ZN => n2994);
   U3006 : XNOR2_X1 port map( A => n3400, B => n3395, ZN => n3264);
   U3007 : NOR2_X1 port map( A1 => n3910, A2 => n4020, ZN => n2223);
   U3008 : XNOR2_X1 port map( A => DataP_alu_a_in_11_port, B => n3254, ZN => 
                           n3318);
   U3009 : AND2_X1 port map( A1 => n2550, A2 => n2428, ZN => n2224);
   U3010 : AND2_X1 port map( A1 => n2136, A2 => n1556, ZN => n2235);
   U3011 : AND2_X1 port map( A1 => n2130, A2 => n1948, ZN => n2236);
   U3012 : AND3_X1 port map( A1 => n2469, A2 => n2470, A3 => 
                           DRAM_ADDRESS_0_port, ZN => n2237);
   U3013 : AND3_X1 port map( A1 => n2469, A2 => n2470, A3 => 
                           DRAM_ADDRESS_1_port, ZN => n2238);
   U3014 : AND2_X1 port map( A1 => n1878, A2 => n3611, ZN => n2239);
   U3015 : AND2_X1 port map( A1 => DataP_alu_a_in_4_port, A2 => n2461, ZN => 
                           n2240);
   U3016 : INV_X1 port map( A => n2312, ZN => n3496);
   U3017 : AND2_X1 port map( A1 => DataP_alu_a_in_17_port, A2 => n2538, ZN => 
                           n2242);
   U3018 : NAND2_X1 port map( A1 => n3272, A2 => n3271, ZN => n2244);
   U3019 : INV_X1 port map( A => Rst, ZN => n3012);
   U3020 : AOI22_X1 port map( A1 => n2149, A2 => n2546, B1 => n2542, B2 => 
                           n2481, ZN => n2282);
   U3021 : NAND2_X1 port map( A1 => n3397, A2 => n2149, ZN => n2283);
   U3022 : NAND2_X1 port map( A1 => n3264, A2 => n2542, ZN => n2284);
   U3023 : XNOR2_X1 port map( A => n2447, B => n3396, ZN => n3397);
   U3024 : NAND2_X1 port map( A1 => n3272, A2 => n2285, ZN => n3639);
   U3025 : AOI21_X1 port map( B1 => n2287, B2 => n2294, A => n2286, ZN => n2285
                           );
   U3026 : NAND2_X1 port map( A1 => n2289, A2 => n3271, ZN => n2286);
   U3027 : INV_X1 port map( A => n3264, ZN => n2287);
   U3028 : NAND2_X1 port map( A1 => n2290, A2 => n2225, ZN => n2425);
   U3029 : NAND2_X1 port map( A1 => n2291, A2 => n2370, ZN => n3576);
   U3030 : NAND2_X1 port map( A1 => n1992, A2 => n3510, ZN => n2291);
   U3031 : XNOR2_X1 port map( A => n2293, B => n2292, ZN => n2577);
   U3032 : INV_X1 port map( A => n3442, ZN => n2292);
   U3033 : NAND2_X1 port map( A1 => n3437, A2 => n2235, ZN => n2293);
   U3034 : AND2_X1 port map( A1 => DataP_alu_a_in_12_port, A2 => n2547, ZN => 
                           n2294);
   U3035 : NAND2_X1 port map( A1 => n2295, A2 => n3631, ZN => n3412);
   U3036 : NAND2_X1 port map( A1 => n3647, A2 => n3409, ZN => n2295);
   U3037 : NAND2_X1 port map( A1 => n2296, A2 => DataP_alu_a_in_18_port, ZN => 
                           n2304);
   U3038 : NAND2_X1 port map( A1 => n2298, A2 => n2297, ZN => n2296);
   U3039 : NAND2_X1 port map( A1 => DataP_alu_b_in_18_port, A2 => n2321, ZN => 
                           n2297);
   U3040 : NAND2_X1 port map( A1 => n3427, A2 => n3510, ZN => n2298);
   U3041 : INV_X1 port map( A => n2000, ZN => n2308);
   U3042 : AND2_X1 port map( A1 => n2354, A2 => n2299, ZN => n3612);
   U3043 : NOR2_X1 port map( A1 => n3426, A2 => n1918, ZN => n2301);
   U3044 : NAND2_X1 port map( A1 => n3281, A2 => n1521, ZN => n2302);
   U3045 : OAI22_X1 port map( A1 => n2305, A2 => n2303, B1 => n1610, B2 => 
                           n2381, ZN => n3459);
   U3046 : NAND4_X1 port map( A1 => n2304, A2 => n3612, A3 => n1552, A4 => 
                           n3611, ZN => n2303);
   U3047 : NAND4_X1 port map( A1 => n3577, A2 => n2378, A3 => n3458, A4 => 
                           n1557, ZN => n2305);
   U3048 : NOR2_X1 port map( A1 => n2184, A2 => n2307, ZN => n2306);
   U3049 : NAND2_X1 port map( A1 => n2403, A2 => n2461, ZN => n3669);
   U3050 : NAND2_X1 port map( A1 => n2309, A2 => n3510, ZN => n2403);
   U3051 : XNOR2_X1 port map( A => n3216, B => sra_131_SH_4_port, ZN => n2309);
   U3052 : NAND2_X1 port map( A1 => n1904, A2 => n2310, ZN => n3070);
   U3053 : NOR2_X1 port map( A1 => n2311, A2 => n3056, ZN => n2310);
   U3054 : OR2_X1 port map( A1 => n3054, A2 => n3055, ZN => n2311);
   U3055 : NAND2_X1 port map( A1 => n1839, A2 => DataP_B_s_12_port, ZN => n2387
                           );
   U3056 : XNOR2_X1 port map( A => n2317, B => n2316, ZN => n3455);
   U3057 : INV_X1 port map( A => n3495, ZN => n2316);
   U3058 : OAI21_X1 port map( B1 => n3565, B2 => n1516, A => n3463, ZN => n2317
                           );
   U3059 : NAND2_X1 port map( A1 => n2318, A2 => n3460, ZN => n3565);
   U3060 : NAND2_X1 port map( A1 => n3592, A2 => n2188, ZN => n2318);
   U3061 : NAND2_X1 port map( A1 => n3269, A2 => n2319, ZN => n2449);
   U3062 : NAND2_X1 port map( A1 => n1866, A2 => DataP_alu_a_in_7_port, ZN => 
                           n3265);
   U3063 : NAND2_X1 port map( A1 => n2322, A2 => n2320, ZN => n3213);
   U3064 : NAND2_X1 port map( A1 => n1950, A2 => n2321, ZN => n2320);
   U3065 : INV_X1 port map( A => n3510, ZN => n2321);
   U3066 : NAND2_X1 port map( A1 => n3209, A2 => n3510, ZN => n2322);
   U3067 : NAND4_X1 port map( A1 => n2323, A2 => n2549, A3 => n2326, A4 => 
                           n2327, ZN => n3220);
   U3068 : NAND2_X1 port map( A1 => n2324, A2 => n2329, ZN => n2323);
   U3069 : NAND2_X1 port map( A1 => n3663, A2 => n2325, ZN => n2324);
   U3070 : INV_X1 port map( A => n3216, ZN => n2325);
   U3071 : NAND2_X1 port map( A1 => n3215, A2 => n2329, ZN => n2326);
   U3072 : NAND4_X1 port map( A1 => n2510, A2 => n3218, A3 => n2328, A4 => 
                           n3663, ZN => n2327);
   U3073 : NOR2_X1 port map( A1 => n2543, A2 => n2003, ZN => n2328);
   U3074 : INV_X1 port map( A => DataP_alu_b_in_3_port, ZN => n2330);
   U3075 : INV_X1 port map( A => n3002, ZN => n2331);
   U3076 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_8_port, ZN => n2332
                           );
   U3077 : NOR2_X1 port map( A1 => DataP_alu_b_in_10_port, A2 => n1572, ZN => 
                           n3262);
   U3078 : NAND2_X1 port map( A1 => n2331, A2 => DRAM_ADDRESS_10_port, ZN => 
                           n2335);
   U3079 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_8_port, ZN => 
                           n2336);
   U3080 : NAND2_X1 port map( A1 => n2337, A2 => n1996, ZN => n3358);
   U3081 : NAND2_X1 port map( A1 => n2339, A2 => n2338, ZN => n2337);
   U3082 : NAND2_X1 port map( A1 => n1907, A2 => n3689, ZN => n2338);
   U3083 : INV_X1 port map( A => n2148, ZN => n2345);
   U3084 : OAI211_X1 port map( C1 => n1984, C2 => n2348, A => n2341, B => n2340
                           , ZN => DataP_PC_reg_N2);
   U3085 : NAND2_X1 port map( A1 => n2148, A2 => n2347, ZN => n2340);
   U3086 : AOI21_X1 port map( B1 => n2431, B2 => n2347, A => n2346, ZN => n2341
                           );
   U3087 : NAND3_X1 port map( A1 => n2436, A2 => n2434, A3 => n443, ZN => n2342
                           );
   U3088 : NAND2_X1 port map( A1 => n1919, A2 => n443, ZN => n2348);
   U3089 : NAND2_X1 port map( A1 => n3498, A2 => n2353, ZN => n3499);
   U3090 : OAI21_X1 port map( B1 => n2351, B2 => n2352, A => n2350, ZN => n3498
                           );
   U3091 : INV_X1 port map( A => n3564, ZN => n2350);
   U3092 : OAI21_X1 port map( B1 => n3462, B2 => n3461, A => n3460, ZN => n2351
                           );
   U3093 : NAND2_X1 port map( A1 => n2462, A2 => n2242, ZN => n2354);
   U3094 : NAND2_X1 port map( A1 => n2358, A2 => n2321, ZN => n2357);
   U3095 : INV_X1 port map( A => n1879, ZN => n2358);
   U3096 : XNOR2_X1 port map( A => n3249, B => n1879, ZN => n3233);
   U3097 : INV_X1 port map( A => n2359, ZN => n2550);
   U3098 : OAI211_X1 port map( C1 => n3532, C2 => n2361, A => n2360, B => n3508
                           , ZN => n2359);
   U3099 : NAND2_X1 port map( A1 => n2553, A2 => n3506, ZN => n2360);
   U3100 : NAND2_X1 port map( A1 => n3504, A2 => n3505, ZN => n3532);
   U3101 : NAND2_X1 port map( A1 => n3506, A2 => n3544, ZN => n2361);
   U3102 : NAND2_X1 port map( A1 => DataP_alu_b_in_20_port, A2 => n2321, ZN => 
                           n2364);
   U3103 : XNOR2_X1 port map( A => n3445, B => DataP_alu_b_in_20_port, ZN => 
                           n2365);
   U3104 : INV_X1 port map( A => DataP_alu_b_in_2_port, ZN => n3011);
   U3105 : NAND2_X1 port map( A1 => n3011, A2 => n3689, ZN => n2366);
   U3106 : OR2_X1 port map( A1 => n2503, A2 => n2467, ZN => n2367);
   U3107 : OAI21_X1 port map( B1 => n2467, B2 => n1550, A => n3510, ZN => n2368
                           );
   U3108 : NAND2_X1 port map( A1 => n3669, A2 => n3204, ZN => n3377);
   U3109 : INV_X1 port map( A => n1638, ZN => n2381);
   U3110 : NAND2_X1 port map( A1 => n3442, A2 => n2383, ZN => n2382);
   U3111 : INV_X1 port map( A => n3510, ZN => n2383);
   U3112 : NAND2_X1 port map( A1 => n1889, A2 => n1592, ZN => n3249);
   U3113 : OR2_X1 port map( A1 => n1988, A2 => n2394, ZN => n2392);
   U3114 : INV_X1 port map( A => n2401, ZN => n2394);
   U3115 : NAND3_X1 port map( A1 => n2422, A2 => n1988, A3 => n2138, ZN => 
                           n2395);
   U3116 : OAI22_X1 port map( A1 => n300, A2 => n3911, B1 => n3910, B2 => n4018
                           , ZN => DataP_PC_reg_N30);
   U3117 : NAND2_X1 port map( A1 => n2424, A2 => n2523, ZN => n3592);
   U3118 : NAND2_X1 port map( A1 => n1528, A2 => n2240, ZN => n3376);
   U3119 : OAI211_X1 port map( C1 => n3488, C2 => n2406, A => n2404, B => n3510
                           , ZN => n2474);
   U3120 : NAND2_X1 port map( A1 => n3488, A2 => n2405, ZN => n2404);
   U3121 : XNOR2_X1 port map( A => n2497, B => n2406, ZN => n2405);
   U3122 : INV_X1 port map( A => DataP_alu_b_in_27_port, ZN => n2406);
   U3123 : NAND2_X1 port map( A1 => n2474, A2 => n2445, ZN => n2444);
   U3124 : NAND2_X1 port map( A1 => n1934, A2 => n2383, ZN => n2407);
   U3125 : NAND3_X1 port map( A1 => n2503, A2 => n2133, A3 => n2241, ZN => 
                           n2409);
   U3126 : NAND2_X1 port map( A1 => n2408, A2 => n3510, ZN => n2457);
   U3127 : XNOR2_X1 port map( A => n2409, B => n1936, ZN => n2408);
   U3128 : XNOR2_X1 port map( A => n1908, B => n3511, ZN => n2413);
   U3129 : NAND2_X1 port map( A1 => n2410, A2 => n2411, ZN => DataP_PC_reg_N32)
                           ;
   U3130 : NAND2_X1 port map( A1 => n2413, A2 => n2412, ZN => n2410);
   U3131 : NAND3_X1 port map( A1 => n3466, A2 => n2131, A3 => n3467, ZN => 
                           n2422);
   U3132 : AOI21_X1 port map( B1 => n2551, B2 => n2224, A => n2427, ZN => n3685
                           );
   U3133 : NAND2_X1 port map( A1 => n1906, A2 => n2552, ZN => n2551);
   U3134 : OAI21_X1 port map( B1 => n2144, B2 => n2432, A => n3351, ZN => n2431
                           );
   U3135 : AOI22_X1 port map( A1 => n3342, A2 => n1876, B1 => n3343, B2 => 
                           n3356, ZN => n2432);
   U3136 : NOR2_X1 port map( A1 => n3356, A2 => n2132, ZN => n2433);
   U3137 : NOR2_X1 port map( A1 => n3357, A2 => n2435, ZN => n2434);
   U3138 : AND2_X1 port map( A1 => DataP_ALU_C_shifter_N82, A2 => n3675, ZN => 
                           n2435);
   U3139 : AOI21_X1 port map( B1 => n3354, B2 => n2438, A => n2437, ZN => n2436
                           );
   U3140 : NOR2_X1 port map( A1 => n3356, A2 => n3355, ZN => n2437);
   U3141 : NOR2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => n2146, ZN => 
                           n2438);
   U3142 : NOR2_X1 port map( A1 => n2440, A2 => n2439, ZN => n2441);
   U3143 : XNOR2_X1 port map( A => n3426, B => n1928, ZN => n3427);
   U3144 : NAND2_X1 port map( A1 => n2441, A2 => n1598, ZN => n3426);
   U3145 : OAI211_X1 port map( C1 => n2474, C2 => DataP_alu_a_in_27_port, A => 
                           n2444, B => n2443, ZN => n3506);
   U3146 : NAND2_X1 port map( A1 => n1912, A2 => n2446, ZN => n2443);
   U3147 : NOR2_X1 port map( A1 => n1912, A2 => n2446, ZN => n2445);
   U3148 : INV_X1 port map( A => n2473, ZN => n2446);
   U3149 : NAND4_X1 port map( A1 => n2142, A2 => n2504, A3 => n1995, A4 => 
                           n3395, ZN => n2447);
   U3150 : NAND2_X1 port map( A1 => n2455, A2 => n2450, ZN => n2448);
   U3151 : NAND2_X1 port map( A1 => n2452, A2 => n2478, ZN => n2451);
   U3152 : INV_X1 port map( A => n3318, ZN => n2452);
   U3153 : NAND2_X1 port map( A1 => n3250, A2 => n2454, ZN => n2453);
   U3154 : AND2_X1 port map( A1 => n1863, A2 => n3510, ZN => n2454);
   U3155 : NAND2_X1 port map( A1 => n2456, A2 => n3268, ZN => n2455);
   U3156 : NAND2_X1 port map( A1 => n3267, A2 => n3266, ZN => n2456);
   U3157 : NAND2_X1 port map( A1 => n2457, A2 => n2502, ZN => n3474);
   U3158 : NAND2_X1 port map( A1 => n2459, A2 => n2458, ZN => n3206);
   U3159 : AOI21_X1 port map( B1 => n2460, B2 => n2236, A => n2139, ZN => n2458
                           );
   U3160 : NAND2_X1 port map( A1 => n1574, A2 => n2460, ZN => n2459);
   U3161 : AOI21_X1 port map( B1 => n2003, B2 => n1948, A => n2375, ZN => n2460
                           );
   U3162 : NAND2_X1 port map( A1 => n3072, A2 => n3073, ZN => n2470);
   U3163 : AOI21_X1 port map( B1 => n2993, B2 => DataP_alu_out_W_0_port, A => 
                           n2237, ZN => n3112);
   U3164 : NOR2_X1 port map( A1 => n2464, A2 => n1938, ZN => n2463);
   U3165 : INV_X1 port map( A => n2493, ZN => n2464);
   U3166 : AND2_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => n2466, ZN => 
                           n2465);
   U3167 : OR2_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n3510, ZN => 
                           n2466);
   U3168 : AND2_X1 port map( A1 => n3470, A2 => DataP_alu_a_in_25_port, ZN => 
                           n3544);
   U3169 : INV_X1 port map( A => DataP_alu_b_in_25_port, ZN => n2467);
   U3170 : INV_X1 port map( A => Rst, ZN => n2468);
   U3171 : AOI21_X1 port map( B1 => n2993, B2 => DataP_alu_out_W_1_port, A => 
                           n2238, ZN => n3115);
   U3172 : NAND2_X1 port map( A1 => DataP_alu_b_in_27_port, A2 => n2478, ZN => 
                           n2473);
   U3173 : XNOR2_X1 port map( A => n2568, B => n523, ZN => n2476);
   U3174 : AND2_X1 port map( A1 => n3059, A2 => n3057, ZN => n2477);
   U3175 : NOR2_X1 port map( A1 => n1581, A2 => DataP_alu_b_in_2_port, ZN => 
                           n2501);
   U3176 : INV_X1 port map( A => n3510, ZN => n2478);
   U3177 : NAND2_X1 port map( A1 => n2571, A2 => n2162, ZN => n2479);
   U3178 : NAND4_X1 port map( A1 => n2480, A2 => n2186, A3 => n3023, A4 => 
                           n2140, ZN => n3063);
   U3179 : INV_X1 port map( A => n2547, ZN => n2481);
   U3180 : OR2_X1 port map( A1 => n3206, A2 => n1920, ZN => n3382);
   U3181 : NAND4_X1 port map( A1 => n1889, A2 => n2142, A3 => n2390, A4 => 
                           n2482, ZN => n2483);
   U3182 : NAND3_X1 port map( A1 => n2485, A2 => n2484, A3 => n2483, ZN => 
                           n3392);
   U3183 : OR2_X1 port map( A1 => n1889, A2 => n3417, ZN => n2484);
   U3184 : NAND2_X1 port map( A1 => n2486, A2 => DataP_alu_b_in_15_port, ZN => 
                           n2485);
   U3185 : NAND2_X1 port map( A1 => n2142, A2 => n2487, ZN => n2486);
   U3186 : OR2_X1 port map( A1 => n1563, A2 => DataP_alu_b_in_17_port, ZN => 
                           n2488);
   U3187 : NAND2_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n3424, ZN => 
                           n2493);
   U3188 : NAND2_X1 port map( A1 => n3437, A2 => n2495, ZN => n2494);
   U3189 : NOR2_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n1580, ZN => 
                           n2495);
   U3190 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_6_port, ZN => n2500
                           );
   U3191 : NAND3_X1 port map( A1 => n1598, A2 => n2136, A3 => n3421, ZN => 
                           n3445);
   U3192 : OAI21_X1 port map( B1 => n2522, B2 => n3689, A => n2521, ZN => n3210
                           );
   U3193 : NAND2_X1 port map( A1 => n3384, A2 => n3385, ZN => n3666);
   U3194 : OR2_X1 port map( A1 => n3210, A2 => DataP_alu_a_in_6_port, ZN => 
                           n3385);
   U3195 : NAND3_X1 port map( A1 => n3087, A2 => n3090, A3 => n3089, ZN => 
                           n2505);
   U3196 : NAND3_X1 port map( A1 => n2511, A2 => n2510, A3 => n3510, ZN => 
                           n2507);
   U3197 : INV_X1 port map( A => n3215, ZN => n2510);
   U3198 : NOR2_X1 port map( A1 => n2003, A2 => DataP_alu_b_in_8_port, ZN => 
                           n2511);
   U3199 : NAND2_X1 port map( A1 => n3425, A2 => n2478, ZN => n2512);
   U3200 : NAND2_X1 port map( A1 => DataP_alu_b_in_6_port, A2 => n3689, ZN => 
                           n2521);
   U3201 : NOR2_X1 port map( A1 => n2529, A2 => n2528, ZN => n297);
   U3202 : NOR2_X1 port map( A1 => n1609, A2 => n1909, ZN => n2528);
   U3203 : NAND2_X1 port map( A1 => n2530, A2 => n1990, ZN => n2529);
   U3204 : NAND2_X1 port map( A1 => n3708, A2 => n2153, ZN => n2530);
   U3205 : OAI211_X1 port map( C1 => n1991, C2 => n2533, A => n2531, B => n2537
                           , ZN => DataP_PC_reg_N33);
   U3206 : NAND2_X1 port map( A1 => n1909, A2 => n2532, ZN => n2531);
   U3207 : NOR2_X1 port map( A1 => n2534, A2 => n3911, ZN => n2532);
   U3208 : NAND2_X1 port map( A1 => n2536, A2 => n1919, ZN => n2533);
   U3209 : NOR2_X1 port map( A1 => n2535, A2 => n2153, ZN => n2534);
   U3210 : INV_X1 port map( A => n3707, ZN => n2535);
   U3211 : NAND2_X1 port map( A1 => n1990, A2 => n1609, ZN => n2536);
   U3212 : OR2_X1 port map( A1 => n3910, A2 => n4023, ZN => n2537);
   U3213 : AND2_X1 port map( A1 => DataP_ALU_C_shifter_N48, A2 => n3007, ZN => 
                           n2539);
   U3214 : NAND2_X1 port map( A1 => n3395, A2 => n2545, ZN => n2547);
   U3215 : NAND2_X1 port map( A1 => n1860, A2 => n2543, ZN => n2548);
   U3216 : INV_X1 port map( A => n3505, ZN => n2553);
   U3217 : INV_X1 port map( A => n3543, ZN => n2556);
   U3218 : OAI211_X1 port map( C1 => n1841, C2 => n3697, A => 
                           DataP_alu_b_in_15_port, B => n3660, ZN => n3403);
   U3219 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_7_port, ZN => n3082
                           );
   U3220 : NAND2_X1 port map( A1 => n1905, A2 => DataP_IMM_s_19_port, ZN => 
                           n3290);
   U3221 : XNOR2_X1 port map( A => DataP_alu_a_in_3_port, B => n1963, ZN => 
                           n3681);
   U3222 : OAI21_X1 port map( B1 => DataP_alu_a_in_13_port, B2 => n1860, A => 
                           n3697, ZN => n3650);
   U3223 : XNOR2_X1 port map( A => DataP_alu_a_in_13_port, B => n1860, ZN => 
                           n3651);
   U3224 : INV_X1 port map( A => DataP_alu_b_in_13_port, ZN => n3396);
   U3225 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_30_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_30_port, ZN => n3132);
   U3226 : AOI22_X1 port map( A1 => n2996, A2 => DRAM_ADDRESS_7_port, B1 => 
                           n2991, B2 => DataP_alu_out_W_7_port, ZN => n3077);
   U3227 : AOI22_X1 port map( A1 => n2996, A2 => DataP_alu_out_M_31_port, B1 =>
                           n2992, B2 => DataP_alu_out_W_31_port, ZN => n3129);
   U3228 : AOI22_X1 port map( A1 => n2995, A2 => DRAM_ADDRESS_9_port, B1 => 
                           n2992, B2 => DataP_alu_out_W_9_port, ZN => n3074);
   U3229 : AOI22_X1 port map( A1 => n2996, A2 => DRAM_ADDRESS_5_port, B1 => 
                           n2991, B2 => DataP_alu_out_W_5_port, ZN => n3120);
   U3230 : AOI22_X1 port map( A1 => n2996, A2 => DRAM_ADDRESS_6_port, B1 => 
                           n2991, B2 => DataP_alu_out_W_6_port, ZN => n3123);
   U3231 : AOI22_X1 port map( A1 => n2995, A2 => DRAM_ADDRESS_4_port, B1 => 
                           n2991, B2 => DataP_alu_out_W_4_port, ZN => n3117);
   U3232 : AOI22_X1 port map( A1 => n2995, A2 => DRAM_ADDRESS_3_port, B1 => 
                           n2992, B2 => DataP_alu_out_W_3_port, ZN => n3108);
   U3233 : AOI22_X1 port map( A1 => n2996, A2 => DRAM_ADDRESS_8_port, B1 => 
                           n2991, B2 => DataP_alu_out_W_8_port, ZN => n3126);
   U3234 : AOI22_X1 port map( A1 => n2995, A2 => DRAM_ADDRESS_2_port, B1 => 
                           n2993, B2 => DataP_alu_out_W_2_port, ZN => n3111);
   U3235 : NAND3_X1 port map( A1 => n1568, A2 => n432, A3 => n2998, ZN => n2560
                           );
   U3236 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_2_port, ZN => 
                           n3096);
   U3237 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_9_port, ZN => 
                           n3047);
   U3238 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_4_port, ZN => 
                           n3100);
   U3239 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_7_port, ZN => 
                           n3080);
   U3240 : NAND2_X1 port map( A1 => n3330, A2 => DataP_alu_out_W_0_port, ZN => 
                           n3088);
   U3241 : NAND2_X1 port map( A1 => n2006, A2 => DataP_alu_out_W_3_port, ZN => 
                           n3092);
   U3242 : NAND2_X1 port map( A1 => n3330, A2 => DataP_alu_out_W_1_port, ZN => 
                           n3084);
   U3243 : NAND2_X1 port map( A1 => n3327, A2 => DataP_B_s_11_port, ZN => n3247
                           );
   U3244 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_2_port, ZN => n3099)
                           ;
   U3245 : NAND2_X1 port map( A1 => n1839, A2 => DataP_B_s_10_port, ZN => n3231
                           );
   U3246 : NAND2_X1 port map( A1 => n1635, A2 => DataP_B_s_4_port, ZN => n3103)
                           ;
   U3247 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_7_port, ZN => n3083)
                           ;
   U3248 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_0_port, ZN => n3091)
                           ;
   U3249 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_3_port, ZN => n3095)
                           ;
   U3250 : NAND2_X1 port map( A1 => n1635, A2 => DataP_B_s_5_port, ZN => n3107)
                           ;
   U3251 : XNOR2_X1 port map( A => n536, B => n2154, ZN => n3059);
   U3252 : INV_X1 port map( A => n2005, ZN => n2566);
   U3253 : NAND2_X1 port map( A1 => n2011, A2 => n3576, ZN => n3582);
   U3254 : NAND2_X1 port map( A1 => n3593, A2 => n2011, ZN => n3461);
   U3255 : NAND2_X1 port map( A1 => n3443, A2 => n2011, ZN => n3460);
   U3256 : XNOR2_X1 port map( A => n1999, B => DataP_Rs1_2_port, ZN => n3055);
   U3257 : XNOR2_X1 port map( A => DataP_Rs2_2_port, B => n1999, ZN => n3042);
   U3258 : XNOR2_X1 port map( A => n530, B => n538, ZN => n3022);
   U3259 : NOR2_X1 port map( A1 => DataP_dest_M_4_port, A2 => 
                           DataP_dest_M_3_port, ZN => n3037);
   U3260 : INV_X1 port map( A => n2574, ZN => n2575);
   U3261 : XNOR2_X1 port map( A => n528, B => n2154, ZN => n3053);
   U3262 : XNOR2_X1 port map( A => n528, B => DataP_Rs2_0_port, ZN => n3041);
   U3263 : XNOR2_X1 port map( A => n528, B => n536, ZN => n3021);
   U3264 : XNOR2_X1 port map( A => n540, B => n524, ZN => n3057);
   U3265 : NAND2_X1 port map( A1 => n3034, A2 => n2161, ZN => n3035);
   U3266 : XNOR2_X1 port map( A => n1987, B => n2572, ZN => n3609);
   U3267 : XNOR2_X1 port map( A => DataP_add_D_1_port, B => DataP_Rs2_1_port, 
                           ZN => n3019);
   U3268 : XNOR2_X1 port map( A => DataP_dest_M_1_port, B => DataP_add_D_1_port
                           , ZN => n3023);
   U3269 : XNOR2_X1 port map( A => DataP_opcode_W_2_port, B => n2151, ZN => 
                           n3018);
   U3270 : XNOR2_X1 port map( A => n3428, B => n1559, ZN => n3436);
   U3271 : NAND2_X1 port map( A1 => n521, A2 => n520, ZN => n3060);
   U3272 : OAI21_X1 port map( B1 => n1948, B2 => n3671, A => n3694, ZN => n3379
                           );
   U3273 : XNOR2_X1 port map( A => DataP_alu_a_in_5_port, B => 
                           lt_x_134_B_5_port, ZN => n3380);
   U3274 : NAND2_X1 port map( A1 => n1518, A2 => DataP_B_s_1_port, ZN => n3087)
                           ;
   U3275 : XNOR2_X1 port map( A => n2568, B => DataP_Rs2_3_port, ZN => n3024);
   U3276 : NAND4_X1 port map( A1 => n1862, A2 => n1871, A3 => n540, A4 => n2568
                           , ZN => n3026);
   U3277 : OAI21_X1 port map( B1 => n2575, B2 => n3682, A => Rst, ZN => 
                           DataP_FORWARDING_BR_N12);
   U3278 : NAND2_X1 port map( A1 => n1850, A2 => n3502, ZN => n3545);
   U3279 : INV_X1 port map( A => n3445, ZN => n3438);
   U3280 : OAI211_X1 port map( C1 => DataP_opcode_M_4_port, C2 => 
                           DataP_opcode_M_0_port, A => DataP_opcode_M_1_port, B
                           => n1895, ZN => n3034);
   U3281 : OAI22_X1 port map( A1 => n1996, A2 => n3362, B1 => n1916, B2 => 
                           n3694, ZN => n3363);
   U3282 : XNOR2_X1 port map( A => DataP_alu_a_in_1_port, B => n1916, ZN => 
                           n3364);
   U3283 : NAND2_X1 port map( A1 => n3069, A2 => n3068, ZN => n3072);
   U3284 : OR2_X1 port map( A1 => n3069, A2 => n3065, ZN => n3066);
   U3285 : AOI21_X1 port map( B1 => n3498, B2 => n3496, A => n3495, ZN => n3466
                           );
   U3286 : AOI21_X1 port map( B1 => sra_131_SH_1_port, B2 => n3693, A => n3697,
                           ZN => n3362);
   U3287 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_11_port, ZN => 
                           n3246);
   U3288 : NAND2_X1 port map( A1 => n2565, A2 => DataP_ir_E_10_port, ZN => 
                           n3230);
   U3289 : OR2_X1 port map( A1 => n2228, A2 => n3002, ZN => n3048);
   U3290 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_4_port, ZN => n3102
                           );
   U3291 : OR2_X1 port map( A1 => n3002, A2 => n2230, ZN => n3081);
   U3292 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_2_port, ZN => n3098
                           );
   U3293 : NAND2_X1 port map( A1 => n2564, A2 => DataP_ir_E_3_port, ZN => n3094
                           );
   U3294 : NAND2_X1 port map( A1 => n3328, A2 => DataP_ir_E_5_port, ZN => n3106
                           );
   U3295 : NAND2_X1 port map( A1 => n3328, A2 => DataP_ir_E_0_port, ZN => n3090
                           );
   U3296 : NAND2_X1 port map( A1 => n3328, A2 => DataP_ir_E_1_port, ZN => n3086
                           );
   U3297 : NAND4_X1 port map( A1 => n2711, A2 => n1913, A3 => n1916, A4 => 
                           n1605, ZN => n2642);
   U3298 : NOR2_X1 port map( A1 => n2846, A2 => n2642, ZN => n2602);
   U3299 : NAND2_X1 port map( A1 => n1605, A2 => n2711, ZN => n2578);
   U3300 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_1_port, B1 => 
                           DataP_alu_a_in_2_port, B2 => n2711, ZN => n2580);
   U3301 : AOI22_X1 port map( A1 => n2839, A2 => n2578, B1 => n2580, B2 => 
                           n2988, ZN => n2591);
   U3302 : NAND2_X1 port map( A1 => n1913, A2 => n2591, ZN => n2612);
   U3303 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_3_port, B1 => 
                           DataP_alu_a_in_4_port, B2 => n2711, ZN => n2579);
   U3304 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_5_port, B1 => 
                           DataP_alu_a_in_6_port, B2 => n2711, ZN => n2582);
   U3305 : AOI22_X1 port map( A1 => n2713, A2 => n2579, B1 => n2582, B2 => 
                           n1916, ZN => n2590);
   U3306 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_7_port, B1 => 
                           DataP_alu_a_in_8_port, B2 => n2711, ZN => n2581);
   U3307 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_9_port, B1 => 
                           DataP_alu_a_in_10_port, B2 => n2711, ZN => n2583);
   U3308 : AOI22_X1 port map( A1 => n2713, A2 => n2581, B1 => n2583, B2 => 
                           n2988, ZN => n2593);
   U3309 : AOI22_X1 port map( A1 => n2842, A2 => n2590, B1 => n2593, B2 => 
                           n1913, ZN => n2611);
   U3310 : AOI22_X1 port map( A1 => n1915, A2 => n2612, B1 => n2611, B2 => 
                           n2064, ZN => n2654);
   U3311 : NOR2_X1 port map( A1 => lt_x_135_B_4_port, A2 => n2697, ZN => 
                           DataP_ALU_C_shifter_N28);
   U3312 : AOI22_X1 port map( A1 => n2709, A2 => n1605, B1 => 
                           DataP_alu_a_in_1_port, B2 => n2711, ZN => n2584);
   U3313 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_2_port, B1 => 
                           DataP_alu_a_in_3_port, B2 => n2710, ZN => n2586);
   U3314 : AOI22_X1 port map( A1 => n2713, A2 => n2584, B1 => n2586, B2 => 
                           n1916, ZN => n2595);
   U3315 : NAND2_X1 port map( A1 => n1913, A2 => n2595, ZN => n2616);
   U3316 : INV_X1 port map( A => n1907, ZN => n2713);
   U3317 : NAND2_X1 port map( A1 => n1930, A2 => n2763, ZN => n2780);
   U3318 : NOR2_X1 port map( A1 => n1915, A2 => n2780, ZN => n2792);
   U3319 : MUX2_X1 port map( A => n2748, B => n2792, S => lt_x_134_B_4_port, Z 
                           => DataP_ALU_C_shifter_N63);
   U3320 : NAND3_X1 port map( A1 => n2781, A2 => n2845, A3 => n2844, ZN => 
                           n2801);
   U3321 : AOI22_X1 port map( A1 => n2842, A2 => n2750, B1 => n2749, B2 => 
                           n1930, ZN => n2782);
   U3322 : AOI22_X1 port map( A1 => n2842, A2 => n2752, B1 => n2751, B2 => 
                           n1930, ZN => n2823);
   U3323 : AOI22_X1 port map( A1 => n1915, A2 => n2782, B1 => n2823, B2 => 
                           n2845, ZN => n2753);
   U3324 : NAND2_X1 port map( A1 => n2847, A2 => n2753, ZN => n2754);
   U3325 : OAI21_X1 port map( B1 => n2065, B2 => n2801, A => n2754, ZN => 
                           DataP_ALU_C_shifter_N64);
   U3326 : NAND3_X1 port map( A1 => n2784, A2 => n2127, A3 => n2844, ZN => 
                           n2802);
   U3327 : AOI22_X1 port map( A1 => n2842, A2 => n2756, B1 => n2755, B2 => 
                           n1930, ZN => n2785);
   U3328 : AOI22_X1 port map( A1 => n2842, A2 => n2758, B1 => n2757, B2 => 
                           n1930, ZN => n2827);
   U3329 : AOI22_X1 port map( A1 => n2846, A2 => n2785, B1 => n2827, B2 => 
                           n2064, ZN => n2759);
   U3330 : NAND2_X1 port map( A1 => n2065, A2 => n2759, ZN => n2760);
   U3331 : OAI21_X1 port map( B1 => n2065, B2 => n2802, A => n2760, ZN => 
                           DataP_ALU_C_shifter_N65);
   U3332 : AND2_X1 port map( A1 => n2065, A2 => n2761, ZN => 
                           DataP_ALU_C_shifter_N66);
   U3333 : AOI22_X1 port map( A1 => n2842, A2 => n2763, B1 => n2762, B2 => 
                           n1930, ZN => n2788);
   U3334 : AOI22_X1 port map( A1 => n2842, A2 => n2765, B1 => n2764, B2 => 
                           n1930, ZN => n2835);
   U3335 : AOI22_X1 port map( A1 => n2846, A2 => n2788, B1 => n2835, B2 => 
                           n2127, ZN => n2774);
   U3336 : AND2_X1 port map( A1 => n2847, A2 => n2774, ZN => 
                           DataP_ALU_C_shifter_N67);
   U3337 : AOI22_X1 port map( A1 => n2846, A2 => n2767, B1 => n2766, B2 => 
                           n2064, ZN => n2800);
   U3338 : AND2_X1 port map( A1 => n2847, A2 => n2800, ZN => 
                           DataP_ALU_C_shifter_N68);
   U3339 : AOI22_X1 port map( A1 => n2846, A2 => n2769, B1 => n2768, B2 => 
                           n2845, ZN => n2808);
   U3340 : AND2_X1 port map( A1 => n2847, A2 => n2808, ZN => 
                           DataP_ALU_C_shifter_N69);
   U3341 : AOI22_X1 port map( A1 => n1914, A2 => DataP_alu_a_in_10_port, B1 => 
                           DataP_alu_a_in_9_port, B2 => n1931, ZN => n2804);
   U3342 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2770, B1 => n2804
                           , B2 => n1916, ZN => n2816);
   U3343 : AOI22_X1 port map( A1 => n2842, A2 => n2771, B1 => n2816, B2 => 
                           n1930, ZN => n2834);
   U3344 : AOI22_X1 port map( A1 => n1914, A2 => DataP_alu_a_in_8_port, B1 => 
                           DataP_alu_a_in_7_port, B2 => n1931, ZN => n2803);
   U3345 : AOI22_X1 port map( A1 => n1914, A2 => DataP_alu_a_in_6_port, B1 => 
                           DataP_alu_a_in_5_port, B2 => n1931, ZN => n2806);
   U3346 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2803, B1 => n2806
                           , B2 => n1916, ZN => n2815);
   U3347 : AOI22_X1 port map( A1 => n1914, A2 => DataP_alu_a_in_4_port, B1 => 
                           DataP_alu_a_in_3_port, B2 => n1931, ZN => n2805);
   U3348 : AOI22_X1 port map( A1 => n2842, A2 => n2815, B1 => n2772, B2 => 
                           n1930, ZN => n2773);
   U3349 : AOI22_X1 port map( A1 => n2846, A2 => n2834, B1 => n2773, B2 => 
                           n2845, ZN => n2775);
   U3350 : MUX2_X1 port map( A => n2775, B => n2774, S => lt_x_134_B_4_port, Z 
                           => DataP_ALU_C_shifter_N51);
   U3351 : NAND2_X1 port map( A1 => n1930, A2 => n2776, ZN => n2778);
   U3352 : AOI22_X1 port map( A1 => n2846, A2 => n2778, B1 => n2777, B2 => 
                           n2064, ZN => n2813);
   U3353 : AND2_X1 port map( A1 => n2065, A2 => n2813, ZN => 
                           DataP_ALU_C_shifter_N70);
   U3354 : AOI22_X1 port map( A1 => n2846, A2 => n2780, B1 => n2779, B2 => 
                           n2064, ZN => n2819);
   U3355 : AND2_X1 port map( A1 => n2065, A2 => n2819, ZN => 
                           DataP_ALU_C_shifter_N71);
   U3356 : NAND2_X1 port map( A1 => n2781, A2 => n2844, ZN => n2783);
   U3357 : AOI22_X1 port map( A1 => n2846, A2 => n2783, B1 => n2782, B2 => 
                           n2127, ZN => n2824);
   U3358 : AND2_X1 port map( A1 => n2065, A2 => n2824, ZN => 
                           DataP_ALU_C_shifter_N72);
   U3359 : NAND2_X1 port map( A1 => n2784, A2 => n2844, ZN => n2786);
   U3360 : AOI22_X1 port map( A1 => n2846, A2 => n2786, B1 => n2785, B2 => 
                           n2127, ZN => n2828);
   U3361 : AND2_X1 port map( A1 => n2847, A2 => n2828, ZN => 
                           DataP_ALU_C_shifter_N73);
   U3362 : NOR2_X1 port map( A1 => n1915, A2 => n2787, ZN => n2832);
   U3363 : AND2_X1 port map( A1 => n2832, A2 => n2847, ZN => 
                           DataP_ALU_C_shifter_N74);
   U3364 : NOR2_X1 port map( A1 => n1915, A2 => n2788, ZN => n2836);
   U3365 : INV_X1 port map( A => n2126, ZN => n2840);
   U3366 : AOI22_X1 port map( A1 => n2713, A2 => n2853, B1 => n2856, B2 => 
                           n2126, ZN => n2867);
   U3367 : AOI22_X1 port map( A1 => n2841, A2 => n2865, B1 => n2867, B2 => 
                           n1913, ZN => n2918);
   U3368 : AOI22_X1 port map( A1 => n2986, A2 => DataP_alu_a_in_23_port, B1 => 
                           DataP_alu_a_in_22_port, B2 => n2985, ZN => n2855);
   U3369 : AOI22_X1 port map( A1 => n2986, A2 => DataP_alu_a_in_19_port, B1 => 
                           DataP_alu_a_in_18_port, B2 => n2985, ZN => n2857);
   U3370 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_17_port, B1 => 
                           DataP_alu_a_in_16_port, B2 => n2985, ZN => n2860);
   U3371 : AOI22_X1 port map( A1 => n2841, A2 => n2866, B1 => n2869, B2 => 
                           n1930, ZN => n2976);
   U3372 : AOI22_X1 port map( A1 => n1915, A2 => n2918, B1 => n2976, B2 => 
                           n2127, ZN => n2893);
   U3373 : AOI22_X1 port map( A1 => n2709, A2 => n1841, B1 => 
                           DataP_alu_a_in_14_port, B2 => n2710, ZN => n2859);
   U3374 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_13_port, B1 => 
                           DataP_alu_a_in_12_port, B2 => n2985, ZN => n2862);
   U3375 : AOI22_X1 port map( A1 => n2713, A2 => n2859, B1 => n2862, B2 => 
                           n2988, ZN => n2868);
   U3376 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_11_port, B1 => 
                           DataP_alu_a_in_10_port, B2 => n2711, ZN => n2861);
   U3377 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_9_port, B1 => 
                           DataP_alu_a_in_8_port, B2 => n2985, ZN => n2932);
   U3378 : AOI22_X1 port map( A1 => n2713, A2 => n2861, B1 => n2932, B2 => 
                           n2988, ZN => n2951);
   U3379 : AOI22_X1 port map( A1 => n2841, A2 => n2868, B1 => n2951, B2 => 
                           n1913, ZN => n2975);
   U3380 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_7_port, B1 => 
                           DataP_alu_a_in_6_port, B2 => n2985, ZN => n2931);
   U3381 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_5_port, B1 => 
                           DataP_alu_a_in_4_port, B2 => n2710, ZN => n2934);
   U3382 : AOI22_X1 port map( A1 => n2840, A2 => n2931, B1 => n2934, B2 => 
                           n2988, ZN => n2950);
   U3383 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_3_port, B1 => 
                           DataP_alu_a_in_2_port, B2 => n2711, ZN => n2933);
   U3384 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_1_port, B1 => 
                           n1605, B2 => n2711, ZN => n2848);
   U3385 : AOI221_X1 port map( B1 => n2933, B2 => n2839, C1 => n2848, C2 => 
                           n2988, A => n2842, ZN => n2849);
   U3386 : AOI21_X1 port map( B1 => n2842, B2 => n2950, A => n2849, ZN => n2850
                           );
   U3387 : AOI22_X1 port map( A1 => n2846, A2 => n2975, B1 => n2850, B2 => 
                           n2064, ZN => n2851);
   U3388 : MUX2_X1 port map( A => n2893, B => n2851, S => n2847, Z => 
                           DataP_ALU_C_shifter_N82);
   U3389 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n1923, B1 => n2852
                           , B2 => n2988, ZN => n2882);
   U3390 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2854, B1 => n2853
                           , B2 => n2988, ZN => n2884);
   U3391 : AOI22_X1 port map( A1 => n2841, A2 => n2882, B1 => n2884, B2 => 
                           n2989, ZN => n2900);
   U3392 : NAND2_X1 port map( A1 => n2846, A2 => DataP_alu_a_in_31_port, ZN => 
                           n2920);
   U3393 : OAI21_X1 port map( B1 => n1915, B2 => n2900, A => n2920, ZN => n2924
                           );
   U3394 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2856, B1 => n2855
                           , B2 => n2988, ZN => n2883);
   U3395 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2858, B1 => n2857
                           , B2 => n2988, ZN => n2886);
   U3396 : AOI22_X1 port map( A1 => n2841, A2 => n2883, B1 => n2886, B2 => 
                           n2989, ZN => n2899);
   U3397 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2860, B1 => n2859
                           , B2 => n2988, ZN => n2885);
   U3398 : AOI22_X1 port map( A1 => n2839, A2 => n2862, B1 => n2861, B2 => 
                           n2988, ZN => n2965);
   U3399 : AOI22_X1 port map( A1 => n2841, A2 => n2885, B1 => n2965, B2 => 
                           n2989, ZN => n2936);
   U3400 : AOI22_X1 port map( A1 => n2846, A2 => n2899, B1 => n2936, B2 => 
                           n2127, ZN => n2863);
   U3401 : MUX2_X1 port map( A => n2924, B => n2863, S => n2847, Z => 
                           DataP_ALU_C_shifter_N92);
   U3402 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_30_port, B1 => 
                           DataP_alu_a_in_29_port, B2 => n2985, ZN => n2871);
   U3403 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_28_port, B1 => 
                           DataP_alu_a_in_27_port, B2 => n2985, ZN => n2873);
   U3404 : AOI22_X1 port map( A1 => n2839, A2 => n2871, B1 => n2873, B2 => 
                           n2988, ZN => n2889);
   U3405 : NOR2_X1 port map( A1 => n1913, A2 => n1923, ZN => n2881);
   U3406 : AOI21_X1 port map( B1 => n1913, B2 => n2889, A => n2881, ZN => n2902
                           );
   U3407 : OAI21_X1 port map( B1 => n2846, B2 => n2902, A => n2920, ZN => n2925
                           );
   U3408 : AOI22_X1 port map( A1 => n2709, A2 => DataP_alu_a_in_26_port, B1 => 
                           DataP_alu_a_in_25_port, B2 => n2711, ZN => n2872);
   U3409 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_24_port, B1 => 
                           DataP_alu_a_in_23_port, B2 => n2710, ZN => n2875);
   U3410 : AOI22_X1 port map( A1 => n2839, A2 => n2872, B1 => n2875, B2 => 
                           n2988, ZN => n2888);
   U3411 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_22_port, B1 => 
                           DataP_alu_a_in_21_port, B2 => n2985, ZN => n2874);
   U3412 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_20_port, B1 => 
                           n1553, B2 => n2985, ZN => n2877);
   U3413 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2874, B1 => n2877
                           , B2 => n2988, ZN => n2891);
   U3414 : AOI22_X1 port map( A1 => n2841, A2 => n2888, B1 => n2891, B2 => 
                           n2989, ZN => n2901);
   U3415 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_18_port, B1 => 
                           DataP_alu_a_in_17_port, B2 => n2985, ZN => n2876);
   U3416 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_16_port, B1 => 
                           n1841, B2 => n2985, ZN => n2879);
   U3417 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2876, B1 => n2879
                           , B2 => n2988, ZN => n2890);
   U3418 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_14_port, B1 => 
                           DataP_alu_a_in_13_port, B2 => n2985, ZN => n2878);
   U3419 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_12_port, B1 => 
                           DataP_alu_a_in_11_port, B2 => n2711, ZN => n2903);
   U3420 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2878, B1 => n2903
                           , B2 => n2988, ZN => n2970);
   U3421 : AOI22_X1 port map( A1 => n2841, A2 => n2890, B1 => n2970, B2 => 
                           n1913, ZN => n2946);
   U3422 : AOI22_X1 port map( A1 => n1915, A2 => n2901, B1 => n2946, B2 => 
                           n2127, ZN => n2864);
   U3423 : MUX2_X1 port map( A => n2925, B => n2864, S => n2065, Z => 
                           DataP_ALU_C_shifter_N93);
   U3424 : AOI21_X1 port map( B1 => n2989, B2 => n2865, A => n2881, ZN => n2911
                           );
   U3425 : OAI21_X1 port map( B1 => n1915, B2 => n2911, A => n2920, ZN => n2927
                           );
   U3426 : AOI22_X1 port map( A1 => n2841, A2 => n2867, B1 => n2866, B2 => 
                           n1913, ZN => n2910);
   U3427 : AOI22_X1 port map( A1 => n2841, A2 => n2869, B1 => n2868, B2 => 
                           n1913, ZN => n2953);
   U3428 : AOI22_X1 port map( A1 => n1915, A2 => n2910, B1 => n2953, B2 => 
                           n2064, ZN => n2870);
   U3429 : MUX2_X1 port map( A => n2927, B => n2870, S => n2847, Z => 
                           DataP_ALU_C_shifter_N94);
   U3430 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n1923, B1 => n2871
                           , B2 => n2988, ZN => n2896);
   U3431 : AOI21_X1 port map( B1 => n1913, B2 => n2896, A => n2881, ZN => n2913
                           );
   U3432 : OAI21_X1 port map( B1 => n2846, B2 => n2913, A => n2920, ZN => n2929
                           );
   U3433 : AOI22_X1 port map( A1 => n2840, A2 => n2873, B1 => n2872, B2 => 
                           n2988, ZN => n2895);
   U3434 : AOI22_X1 port map( A1 => n2839, A2 => n2875, B1 => n2874, B2 => 
                           n2988, ZN => n2898);
   U3435 : AOI22_X1 port map( A1 => n2841, A2 => n2895, B1 => n2898, B2 => 
                           n1913, ZN => n2912);
   U3436 : AOI22_X1 port map( A1 => n2839, A2 => n2877, B1 => n2876, B2 => 
                           n2988, ZN => n2897);
   U3437 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2879, B1 => n2878
                           , B2 => n2988, ZN => n2904);
   U3438 : AOI22_X1 port map( A1 => n2841, A2 => n2897, B1 => n2904, B2 => 
                           n1913, ZN => n2960);
   U3439 : AOI22_X1 port map( A1 => n1915, A2 => n2912, B1 => n2960, B2 => 
                           n2064, ZN => n2880);
   U3440 : MUX2_X1 port map( A => n2929, B => n2880, S => n2065, Z => 
                           DataP_ALU_C_shifter_N95);
   U3441 : AOI21_X1 port map( B1 => n1913, B2 => n2882, A => n2881, ZN => n2915
                           );
   U3442 : OAI21_X1 port map( B1 => n1915, B2 => n2915, A => n2920, ZN => n2938
                           );
   U3443 : AOI22_X1 port map( A1 => n2841, A2 => n2884, B1 => n2883, B2 => 
                           n1913, ZN => n2914);
   U3444 : AOI22_X1 port map( A1 => n2841, A2 => n2886, B1 => n2885, B2 => 
                           n1913, ZN => n2966);
   U3445 : AOI22_X1 port map( A1 => n2846, A2 => n2914, B1 => n2966, B2 => 
                           n2127, ZN => n2887);
   U3446 : MUX2_X1 port map( A => n2938, B => n2887, S => n2847, Z => 
                           DataP_ALU_C_shifter_N96);
   U3447 : NAND2_X1 port map( A1 => lt_x_134_B_4_port, A2 => 
                           DataP_alu_a_in_31_port, ZN => n2923);
   U3448 : AOI22_X1 port map( A1 => n2841, A2 => n2889, B1 => n2888, B2 => 
                           n1913, ZN => n2916);
   U3449 : AOI22_X1 port map( A1 => n2841, A2 => n2891, B1 => n2890, B2 => 
                           n1913, ZN => n2972);
   U3450 : AOI221_X1 port map( B1 => n2916, B2 => n2846, C1 => n2972, C2 => 
                           n2064, A => lt_x_134_B_4_port, ZN => n2892);
   U3451 : OR2_X1 port map( A1 => n2981, A2 => n2892, ZN => 
                           DataP_ALU_C_shifter_N97);
   U3452 : AOI21_X1 port map( B1 => n2847, B2 => n2893, A => n2981, ZN => n2894
                           );
   U3453 : AOI22_X1 port map( A1 => n2841, A2 => n2896, B1 => n2895, B2 => 
                           n1913, ZN => n2921);
   U3454 : AOI22_X1 port map( A1 => n2841, A2 => n2898, B1 => n2897, B2 => 
                           n1913, ZN => n2979);
   U3455 : MUX2_X1 port map( A => n2921, B => n2979, S => n2064, Z => n2909);
   U3456 : OAI21_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2909, A => n2923,
                           ZN => DataP_ALU_C_shifter_N99);
   U3457 : MUX2_X1 port map( A => n2900, B => n2899, S => n2127, Z => n2937);
   U3458 : OAI21_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2937, A => n2923,
                           ZN => DataP_ALU_C_shifter_N100);
   U3459 : MUX2_X1 port map( A => n2902, B => n2901, S => n2064, Z => n2949);
   U3460 : OAI21_X1 port map( B1 => lt_x_135_B_4_port, B2 => n2949, A => n2923,
                           ZN => DataP_ALU_C_shifter_N101);
   U3461 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_10_port, B1 => 
                           DataP_alu_a_in_9_port, B2 => n2710, ZN => n2941);
   U3462 : AOI22_X1 port map( A1 => n1612, A2 => n2903, B1 => n2941, B2 => 
                           n2988, ZN => n2958);
   U3463 : AOI22_X1 port map( A1 => n2841, A2 => n2904, B1 => n2958, B2 => 
                           n2989, ZN => n2978);
   U3464 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_8_port, B1 => 
                           DataP_alu_a_in_7_port, B2 => n2710, ZN => n2940);
   U3465 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_6_port, B1 => 
                           DataP_alu_a_in_5_port, B2 => n2985, ZN => n2943);
   U3466 : AOI22_X1 port map( A1 => n2839, A2 => n2940, B1 => n2943, B2 => 
                           n2988, ZN => n2957);
   U3467 : AOI22_X1 port map( A1 => n2987, A2 => DataP_alu_a_in_4_port, B1 => 
                           DataP_alu_a_in_3_port, B2 => n2711, ZN => n2942);
   U3468 : AOI22_X1 port map( A1 => n2841, A2 => n2957, B1 => n2905, B2 => 
                           n2989, ZN => n2906);
   U3469 : AOI22_X1 port map( A1 => n1915, A2 => n2978, B1 => n2906, B2 => 
                           n2845, ZN => n2907);
   U3470 : NAND2_X1 port map( A1 => n2847, A2 => n2907, ZN => n2908);
   U3471 : OAI21_X1 port map( B1 => n2847, B2 => n2909, A => n2908, ZN => 
                           DataP_ALU_C_shifter_N83);
   U3472 : MUX2_X1 port map( A => n2911, B => n2910, S => n2127, Z => n2956);
   U3473 : OAI21_X1 port map( B1 => lt_x_135_B_4_port, B2 => n2956, A => n2923,
                           ZN => DataP_ALU_C_shifter_N102);
   U3474 : MUX2_X1 port map( A => n2913, B => n2912, S => n2064, Z => n2963);
   U3475 : OAI21_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2963, A => n2923,
                           ZN => DataP_ALU_C_shifter_N103);
   U3476 : MUX2_X1 port map( A => n2915, B => n2914, S => n2127, Z => n2968);
   U3477 : OAI21_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2968, A => n2923,
                           ZN => DataP_ALU_C_shifter_N104);
   U3478 : OAI21_X1 port map( B1 => n1915, B2 => n2916, A => n2920, ZN => n2917
                           );
   U3479 : OAI21_X1 port map( B1 => lt_x_135_B_4_port, B2 => n2982, A => n2923,
                           ZN => DataP_ALU_C_shifter_N105);
   U3480 : OAI21_X1 port map( B1 => n1915, B2 => n2918, A => n2920, ZN => n2919
                           );
   U3481 : OAI21_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2983, A => n2923,
                           ZN => DataP_ALU_C_shifter_N106);
   U3482 : OAI21_X1 port map( B1 => n2846, B2 => n2921, A => n2920, ZN => n2922
                           );
   U3483 : OAI21_X1 port map( B1 => lt_x_134_B_4_port, B2 => n2984, A => n2923,
                           ZN => DataP_ALU_C_shifter_N107);
   U3484 : AOI21_X1 port map( B1 => n2065, B2 => n2927, A => n2981, ZN => n2928
                           );
   U3485 : AOI22_X1 port map( A1 => sra_131_SH_1_port, A2 => n2932, B1 => n2931
                           , B2 => n2988, ZN => n2964);
   U3486 : AOI22_X1 port map( A1 => n1612, A2 => n2934, B1 => n2933, B2 => 
                           n2988, ZN => n2935);
   U3487 : AOI21_X1 port map( B1 => n2847, B2 => n2938, A => n2981, ZN => n2939
                           );
   U3488 : AOI22_X1 port map( A1 => n2840, A2 => n2941, B1 => n2940, B2 => 
                           n2988, ZN => n2969);
   U3489 : AOI22_X1 port map( A1 => n2839, A2 => n2943, B1 => n2942, B2 => 
                           n2988, ZN => n2944);
   U3490 : AOI22_X1 port map( A1 => n2841, A2 => n2969, B1 => n2944, B2 => 
                           n2989, ZN => n2945);
   U3491 : AOI22_X1 port map( A1 => n2846, A2 => n2946, B1 => n2945, B2 => 
                           n2064, ZN => n2947);
   U3492 : NAND2_X1 port map( A1 => n2065, A2 => n2947, ZN => n2948);
   U3493 : AOI22_X1 port map( A1 => n2841, A2 => n2951, B1 => n2950, B2 => 
                           n2989, ZN => n2952);
   U3494 : AOI22_X1 port map( A1 => n2846, A2 => n2953, B1 => n2952, B2 => 
                           n2845, ZN => n2954);
   U3495 : NAND2_X1 port map( A1 => n2847, A2 => n2954, ZN => n2955);
   U3496 : AOI22_X1 port map( A1 => n2842, A2 => n2958, B1 => n2957, B2 => 
                           n2989, ZN => n2959);
   U3497 : AOI22_X1 port map( A1 => n1915, A2 => n2960, B1 => n2959, B2 => 
                           n2845, ZN => n2961);
   U3498 : NAND2_X1 port map( A1 => n2065, A2 => n2961, ZN => n2962);
   U3499 : AOI22_X1 port map( A1 => n2841, A2 => n2970, B1 => n2969, B2 => 
                           n2989, ZN => n2971);
   U3500 : AOI22_X1 port map( A1 => n1915, A2 => n2972, B1 => n2971, B2 => 
                           n2845, ZN => n2973);
   U3501 : NAND2_X1 port map( A1 => n2847, A2 => n2973, ZN => n2974);
   U3502 : OAI21_X1 port map( B1 => n2065, B2 => n2982, A => n2974, ZN => 
                           DataP_ALU_C_shifter_N89);
   U3503 : INV_X1 port map( A => n2985, ZN => n2986);
   U3504 : INV_X1 port map( A => n2841, ZN => n2989);
   U3505 : INV_X1 port map( A => n2994, ZN => n2993);
   U3506 : INV_X1 port map( A => n1845, ZN => n2997);
   U3507 : XOR2_X1 port map( A => DataP_dest_M_4_port, B => n524, Z => n3052);
   U3508 : XOR2_X1 port map( A => DataP_dest_M_3_port, B => n523, Z => n3051);
   U3509 : NAND3_X1 port map( A1 => n3053, A2 => n3052, A3 => n3051, ZN => 
                           n3056);
   U3510 : NAND3_X1 port map( A1 => n2994, A2 => n432, A3 => n1844, ZN => n3194
                           );
   U3511 : NAND3_X1 port map( A1 => n3199, A2 => n443, A3 => 
                           ALU_OPCODE_i_3_port, ZN => n3200);
   U3512 : NAND3_X1 port map( A1 => ALU_OPCODE_i_0_port, A2 => 
                           ALU_OPCODE_i_3_port, A3 => n3222, ZN => n3695);
   U3513 : NAND3_X1 port map( A1 => DataP_alu_a_in_11_port, A2 => n3689, A3 => 
                           n1572, ZN => n3271);
   U3514 : XOR2_X1 port map( A => n3273, B => n1601, Z => n3279);
   U3515 : NAND3_X1 port map( A1 => DataP_alu_a_in_12_port, A2 => n3693, A3 => 
                           n1880, ZN => n3274);
   U3516 : MUX2_X1 port map( A => n3341, B => n3343, S => ALU_OPCODE_i_1_port, 
                           Z => n3342);
   U3517 : NAND3_X1 port map( A1 => n1602, A2 => n3343, A3 => n2144, ZN => 
                           n3344);
   U3518 : NAND3_X1 port map( A1 => n3348, A2 => ALU_OPCODE_i_3_port, A3 => 
                           n2150, ZN => n3355);
   U3519 : XOR2_X1 port map( A => n3361, B => n3360, Z => n3367);
   U3520 : MUX2_X1 port map( A => n3391, B => n3402, S => n3689, Z => n3393);
   U3521 : NAND3_X1 port map( A1 => n1841, A2 => n3689, A3 => 
                           DataP_alu_b_in_15_port, ZN => n3415);
   U3522 : NAND3_X1 port map( A1 => n3434, A2 => n3433, A3 => n3432, ZN => 
                           n3435);
   U3523 : NAND3_X1 port map( A1 => n3438, A2 => n3468, A3 => n1933, ZN => 
                           n3439);
   U3524 : MUX2_X1 port map( A => DataP_alu_b_in_23_port, B => n3440, S => 
                           n3510, Z => n3464);
   U3525 : MUX2_X1 port map( A => n3446, B => n1933, S => n3689, Z => n3447);
   U3526 : MUX2_X1 port map( A => n3469, B => DataP_alu_b_in_24_port, S => 
                           n3689, Z => n3471);
   U3527 : MUX2_X1 port map( A => n3492, B => n3491, S => n3510, Z => n3493);
   U3528 : NAND3_X1 port map( A1 => n1849, A2 => n3499, A3 => n3500, ZN => 
                           n3503);
   U3529 : NAND3_X1 port map( A1 => n3540, A2 => n3539, A3 => n3538, ZN => 
                           n3541);
   U3530 : XOR2_X1 port map( A => n3545, B => n3546, Z => n3553);
   U3531 : NAND3_X1 port map( A1 => n3551, A2 => n3550, A3 => n3549, ZN => 
                           n3552);
   U3532 : NAND3_X1 port map( A1 => n3561, A2 => n3560, A3 => n3559, ZN => 
                           n3562);
   U3533 : XOR2_X1 port map( A => n3582, B => n3581, Z => n3591);
   U3534 : XOR2_X1 port map( A => n1533, B => n1989, Z => n3601);
   U3535 : NAND3_X1 port map( A1 => n3599, A2 => n3598, A3 => n3597, ZN => 
                           n3600);
   U3536 : NAND3_X1 port map( A1 => n3619, A2 => n3618, A3 => n3617, ZN => 
                           n3620);
   U3537 : XOR2_X1 port map( A => n2239, B => n1986, Z => n3630);
   U3538 : NAND3_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => n3693, A3 => 
                           DataP_alu_b_in_16_port, ZN => n3623);
   U3539 : NAND3_X1 port map( A1 => n3628, A2 => n3627, A3 => n3626, ZN => 
                           n3629);
   U3540 : NAND3_X1 port map( A1 => DataP_alu_a_in_13_port, A2 => n3693, A3 => 
                           n1860, ZN => n3649);
   U3541 : MUX2_X1 port map( A => n3661, B => n3679, S => DataP_alu_a_in_8_port
                           , Z => n3664);
   U3542 : NAND3_X1 port map( A1 => n3696, A2 => n3695, A3 => n3694, ZN => 
                           n3698);
   U3543 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_30_port, B1 => 
                           DataP_pc_out_30_port, B2 => n3010, ZN => n3769);
   U3544 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_28_port, B1 => 
                           DataP_pc_out_28_port, B2 => n3010, ZN => n3753);
   U3545 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_26_port, B1 => 
                           DataP_pc_out_26_port, B2 => n3010, ZN => n3754);
   U3546 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_24_port, B1 => 
                           DataP_pc_out_24_port, B2 => n3010, ZN => n3764);
   U3547 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_22_port, B1 => 
                           DataP_pc_out_22_port, B2 => n3010, ZN => n3763);
   U3548 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_20_port, B1 => 
                           DataP_pc_out_20_port, B2 => n3010, ZN => n3760);
   U3549 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_18_port, B1 => 
                           DataP_pc_out_18_port, B2 => n3010, ZN => n3765);
   U3550 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_16_port, B1 => 
                           DataP_pc_out_16_port, B2 => n3010, ZN => n3759);
   U3551 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_14_port, B1 => DataP_pc_out_14_port, 
                           B2 => n3010, ZN => n3758);
   U3552 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_12_port, B1 => DataP_pc_out_12_port, 
                           B2 => n3010, ZN => n3766);
   U3553 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_10_port, B1 => 
                           DataP_pc_out_10_port, B2 => n3010, ZN => n3774);
   U3554 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_8_port, B1 => IRAM_ADDRESS_6_port, B2 
                           => n3010, ZN => n3736);
   U3555 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_6_port, B1 => IRAM_ADDRESS_4_port, B2 
                           => n3010, ZN => n3742);
   U3556 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_4_port, B1 => IRAM_ADDRESS_2_port, B2 
                           => n3010, ZN => n3749);
   U3557 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_2_port, B1 => IRAM_ADDRESS_0_port, B2 
                           => n3010, ZN => DataP_NPC_add_N3);
   U3558 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_3_port, B1 => IRAM_ADDRESS_1_port, B2 
                           => n3010, ZN => n3751);
   U3559 : NOR2_X1 port map( A1 => DataP_NPC_add_N3, A2 => n3751, ZN => n3750);
   U3560 : INV_X1 port map( A => n3750, ZN => n3748);
   U3561 : NOR2_X1 port map( A1 => n3749, A2 => n3748, ZN => n3747);
   U3562 : OAI221_X1 port map( B1 => n1940, B2 => IRAM_ADDRESS_3_port, C1 => 
                           n3010, C2 => DataP_npc_pre_5_port, A => n3747, ZN =>
                           n3743);
   U3563 : NOR2_X1 port map( A1 => n3742, A2 => n3743, ZN => n3741);
   U3564 : OAI221_X1 port map( B1 => n1940, B2 => IRAM_ADDRESS_5_port, C1 => 
                           n3010, C2 => DataP_npc_pre_7_port, A => n3741, ZN =>
                           n3737);
   U3565 : NOR2_X1 port map( A1 => n3736, A2 => n3737, ZN => n3735);
   U3566 : OAI221_X1 port map( B1 => n1940, B2 => IRAM_ADDRESS_7_port, C1 => 
                           n3010, C2 => DataP_npc_pre_9_port, A => n3735, ZN =>
                           n3773);
   U3567 : NOR2_X1 port map( A1 => n3774, A2 => n3773, ZN => n3731);
   U3568 : MUX2_X1 port map( A => DataP_pc_out_11_port, B => 
                           DataP_npc_pre_11_port, S => n1940, Z => n3770);
   U3569 : NAND2_X1 port map( A1 => n3731, A2 => n3770, ZN => n3730);
   U3570 : NOR2_X1 port map( A1 => n3766, A2 => n3730, ZN => n3729);
   U3571 : MUX2_X1 port map( A => DataP_pc_out_13_port, B => 
                           DataP_npc_pre_13_port, S => n1940, Z => n3761);
   U3572 : NAND2_X1 port map( A1 => n3729, A2 => n3761, ZN => n3728);
   U3573 : NOR2_X1 port map( A1 => n3758, A2 => n3728, ZN => n3727);
   U3574 : MUX2_X1 port map( A => DataP_pc_out_15_port, B => 
                           DataP_npc_pre_15_port, S => n1940, Z => n3757);
   U3575 : NAND2_X1 port map( A1 => n3727, A2 => n3757, ZN => n3726);
   U3576 : NOR2_X1 port map( A1 => n3759, A2 => n3726, ZN => n3725);
   U3577 : MUX2_X1 port map( A => DataP_pc_out_17_port, B => 
                           DataP_npc_pre_17_port, S => n1940, Z => n3767);
   U3578 : NAND2_X1 port map( A1 => n3725, A2 => n3767, ZN => n3724);
   U3579 : NOR2_X1 port map( A1 => n3765, A2 => n3724, ZN => n3723);
   U3580 : MUX2_X1 port map( A => DataP_pc_out_19_port, B => 
                           DataP_npc_pre_19_port, S => n1940, Z => n3762);
   U3581 : NAND2_X1 port map( A1 => n3723, A2 => n3762, ZN => n3722);
   U3582 : NOR2_X1 port map( A1 => n3760, A2 => n3722, ZN => n3721);
   U3583 : MUX2_X1 port map( A => DataP_pc_out_21_port, B => 
                           DataP_npc_pre_21_port, S => n1940, Z => n3771);
   U3584 : NAND2_X1 port map( A1 => n3721, A2 => n3771, ZN => n3720);
   U3585 : NOR2_X1 port map( A1 => n3763, A2 => n3720, ZN => n3719);
   U3586 : MUX2_X1 port map( A => DataP_pc_out_23_port, B => 
                           DataP_npc_pre_23_port, S => n1940, Z => n3772);
   U3587 : NAND2_X1 port map( A1 => n3719, A2 => n3772, ZN => n3718);
   U3588 : NOR2_X1 port map( A1 => n3764, A2 => n3718, ZN => n3717);
   U3589 : MUX2_X1 port map( A => DataP_pc_out_25_port, B => 
                           DataP_npc_pre_25_port, S => n1940, Z => n3755);
   U3590 : NAND2_X1 port map( A1 => n3717, A2 => n3755, ZN => n3716);
   U3591 : NOR2_X1 port map( A1 => n3754, A2 => n3716, ZN => n3715);
   U3592 : MUX2_X1 port map( A => DataP_pc_out_27_port, B => 
                           DataP_npc_pre_27_port, S => n1940, Z => n3756);
   U3593 : NAND2_X1 port map( A1 => n3715, A2 => n3756, ZN => n3714);
   U3594 : NOR2_X1 port map( A1 => n3753, A2 => n3714, ZN => n3713);
   U3595 : MUX2_X1 port map( A => DataP_pc_out_29_port, B => 
                           DataP_npc_pre_29_port, S => n1940, Z => n3768);
   U3596 : NAND2_X1 port map( A1 => n3713, A2 => n3768, ZN => n3712);
   U3597 : NOR2_X1 port map( A1 => n3769, A2 => n3712, ZN => n3752);
   U3598 : AOI21_X1 port map( B1 => n3769, B2 => n3712, A => n3752, ZN => 
                           DataP_NPC_add_N31);
   U3599 : XOR2_X1 port map( A => n3713, B => n3768, Z => DataP_NPC_add_N30);
   U3600 : AOI21_X1 port map( B1 => n3753, B2 => n3714, A => n3713, ZN => 
                           DataP_NPC_add_N29);
   U3601 : XOR2_X1 port map( A => n3715, B => n3756, Z => DataP_NPC_add_N28);
   U3602 : AOI21_X1 port map( B1 => n3754, B2 => n3716, A => n3715, ZN => 
                           DataP_NPC_add_N27);
   U3603 : XOR2_X1 port map( A => n3717, B => n3755, Z => DataP_NPC_add_N26);
   U3604 : AOI21_X1 port map( B1 => n3764, B2 => n3718, A => n3717, ZN => 
                           DataP_NPC_add_N25);
   U3605 : XOR2_X1 port map( A => n3719, B => n3772, Z => DataP_NPC_add_N24);
   U3606 : AOI21_X1 port map( B1 => n3763, B2 => n3720, A => n3719, ZN => 
                           DataP_NPC_add_N23);
   U3607 : XOR2_X1 port map( A => n3721, B => n3771, Z => DataP_NPC_add_N22);
   U3608 : AOI21_X1 port map( B1 => n3760, B2 => n3722, A => n3721, ZN => 
                           DataP_NPC_add_N21);
   U3609 : XOR2_X1 port map( A => n3723, B => n3762, Z => DataP_NPC_add_N20);
   U3610 : AOI21_X1 port map( B1 => n3765, B2 => n3724, A => n3723, ZN => 
                           DataP_NPC_add_N19);
   U3611 : XOR2_X1 port map( A => n3725, B => n3767, Z => DataP_NPC_add_N18);
   U3612 : AOI21_X1 port map( B1 => n3759, B2 => n3726, A => n3725, ZN => 
                           DataP_NPC_add_N17);
   U3613 : XOR2_X1 port map( A => n3727, B => n3757, Z => DataP_NPC_add_N16);
   U3614 : AOI21_X1 port map( B1 => n3758, B2 => n3728, A => n3727, ZN => 
                           DataP_NPC_add_N15);
   U3615 : XOR2_X1 port map( A => n3729, B => n3761, Z => DataP_NPC_add_N14);
   U3616 : AOI21_X1 port map( B1 => n3766, B2 => n3730, A => n3729, ZN => 
                           DataP_NPC_add_N13);
   U3617 : XOR2_X1 port map( A => n3731, B => n3770, Z => DataP_NPC_add_N12);
   U3618 : AOI21_X1 port map( B1 => n3774, B2 => n3773, A => n3731, ZN => 
                           DataP_NPC_add_N11);
   U3619 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_9_port, B1 => 
                           IRAM_ADDRESS_7_port, B2 => n3010, ZN => n3734);
   U3620 : INV_X1 port map( A => n3735, ZN => n3733);
   U3621 : INV_X1 port map( A => n3773, ZN => n3732);
   U3622 : AOI21_X1 port map( B1 => n3734, B2 => n3733, A => n3732, ZN => 
                           DataP_NPC_add_N10);
   U3623 : AOI21_X1 port map( B1 => n3736, B2 => n3737, A => n3735, ZN => 
                           DataP_NPC_add_N9);
   U3624 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_7_port, B1 => 
                           IRAM_ADDRESS_5_port, B2 => n3010, ZN => n3740);
   U3625 : INV_X1 port map( A => n3741, ZN => n3739);
   U3626 : INV_X1 port map( A => n3737, ZN => n3738);
   U3627 : AOI21_X1 port map( B1 => n3740, B2 => n3739, A => n3738, ZN => 
                           DataP_NPC_add_N8);
   U3628 : AOI21_X1 port map( B1 => n3742, B2 => n3743, A => n3741, ZN => 
                           DataP_NPC_add_N7);
   U3629 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_5_port, B1 => 
                           IRAM_ADDRESS_3_port, B2 => n3010, ZN => n3746);
   U3630 : INV_X1 port map( A => n3747, ZN => n3745);
   U3631 : INV_X1 port map( A => n3743, ZN => n3744);
   U3632 : AOI21_X1 port map( B1 => n3746, B2 => n3745, A => n3744, ZN => 
                           DataP_NPC_add_N6);
   U3633 : AOI21_X1 port map( B1 => n3749, B2 => n3748, A => n3747, ZN => 
                           DataP_NPC_add_N5);
   U3634 : AOI21_X1 port map( B1 => n3751, B2 => DataP_NPC_add_N3, A => n3750, 
                           ZN => DataP_NPC_add_N4);
   U3635 : AOI22_X1 port map( A1 => n1940, A2 => DataP_npc_pre_31_port, B1 => 
                           DataP_pc_out_31_port, B2 => n3010, ZN => n3775);
   U3636 : XNOR2_X1 port map( A => n3775, B => n3752, ZN => DataP_NPC_add_N32);
   n4024 <= '0';
   n1513 <= '1';
   U3639 : NAND2_X1 port map( A1 => IR_CU_28, A2 => n516, ZN => n3781);
   U3640 : NOR2_X1 port map( A1 => n3955, A2 => n3781, ZN => n606);
   U3641 : NAND2_X1 port map( A1 => IR_CU_27, A2 => n497, ZN => n3951);
   U3642 : NOR2_X1 port map( A1 => n514, A2 => n515, ZN => n3976);
   U3643 : NAND3_X1 port map( A1 => IR_CU_31, A2 => n3976, A3 => n510, ZN => 
                           n3813);
   U3644 : NOR2_X1 port map( A1 => IR_CU_27, A2 => n497, ZN => n3797);
   U3645 : INV_X1 port map( A => n3976, ZN => n3977);
   U3646 : NOR2_X1 port map( A1 => n3781, A2 => n3977, ZN => n3814);
   U3647 : NOR3_X1 port map( A1 => IR_CU_27, A2 => n3955, A3 => n516, ZN => 
                           n3847);
   U3648 : AOI22_X1 port map( A1 => IR_CU_31, A2 => n3966, B1 => n2141, B2 => 
                           n504, ZN => n3776);
   U3649 : NAND2_X1 port map( A1 => n515, A2 => n510, ZN => n3845);
   U3650 : NOR3_X1 port map( A1 => n514, A2 => n2129, A3 => n3781, ZN => n3796)
                           ;
   U3651 : AOI22_X1 port map( A1 => n3856, A2 => n606, B1 => n3853, B2 => n3796
                           , ZN => n3798);
   U3652 : OAI211_X1 port map( C1 => n3776, C2 => n3845, A => n3798, B => n3956
                           , ZN => n3777);
   U3653 : AOI211_X1 port map( C1 => n3797, C2 => n3814, A => n3847, B => n3777
                           , ZN => n3788);
   U3654 : NOR4_X1 port map( A1 => IR_CU_8_port, A2 => IR_CU_6_port, A3 => 
                           IR_CU_7_port, A4 => IR_CU_9_port, ZN => n3778);
   U3655 : NAND3_X1 port map( A1 => n3953, A2 => n484, A3 => n3778, ZN => n3790
                           );
   U3656 : NOR2_X1 port map( A1 => n479, A2 => n3790, ZN => n3824);
   U3657 : NAND2_X1 port map( A1 => IR_CU_5_port, A2 => n3824, ZN => n3802);
   U3658 : NOR3_X1 port map( A1 => n477, A2 => n2128, A3 => n3802, ZN => n3786)
                           ;
   U3659 : NOR3_X1 port map( A1 => n478, A2 => n3790, A3 => n2135, ZN => n3804)
                           ;
   U3660 : NAND2_X1 port map( A1 => n3804, A2 => n476, ZN => n3806);
   U3661 : OAI21_X1 port map( B1 => n476, B2 => n479, A => n2128, ZN => n3779);
   U3662 : OAI211_X1 port map( C1 => n479, C2 => n2128, A => n3779, B => n477, 
                           ZN => n3780);
   U3663 : NAND2_X1 port map( A1 => IR_CU_5_port, A2 => n480, ZN => n3836);
   U3664 : AOI221_X1 port map( B1 => n3790, B2 => n3806, C1 => n3780, C2 => 
                           n3806, A => n3836, ZN => n3785);
   U3665 : INV_X1 port map( A => n3786, ZN => n3833);
   U3666 : NOR3_X1 port map( A1 => n3795, A2 => n3955, A3 => n3951, ZN => n3821
                           );
   U3667 : INV_X1 port map( A => n3781, ZN => n3782);
   U3668 : NAND3_X1 port map( A1 => n514, A2 => n3782, A3 => n2129, ZN => n3817
                           );
   U3669 : NAND4_X1 port map( A1 => n3804, A2 => IR_CU_1_port, A3 => n480, A4 
                           => n482, ZN => n3827);
   U3670 : OAI21_X1 port map( B1 => n504, B2 => n3817, A => n3827, ZN => n3801)
                           ;
   U3671 : AOI211_X1 port map( C1 => n3856, C2 => n3796, A => n3821, B => n3801
                           , ZN => n3784);
   U3672 : NAND3_X1 port map( A1 => n3966, A2 => n3976, A3 => n510, ZN => n3783
                           );
   U3673 : OAI211_X1 port map( C1 => n3833, C2 => n476, A => n3784, B => n3783,
                           ZN => n3792);
   U3674 : AOI211_X1 port map( C1 => n3786, C2 => IR_CU_4_port, A => n3785, B 
                           => n3792, ZN => n3787);
   U3675 : OAI211_X1 port map( C1 => n3951, C2 => n3813, A => n3788, B => n3787
                           , ZN => CU_I_aluOpcode_i_0_port);
   U3676 : INV_X1 port map( A => n3795, ZN => n3968);
   U3677 : NAND2_X1 port map( A1 => n3968, A2 => IR_CU_27, ZN => n3954);
   U3678 : NOR2_X1 port map( A1 => IR_CU_1_port, A2 => n478, ZN => n3789);
   U3679 : AOI22_X1 port map( A1 => IR_CU_1_port, A2 => n478, B1 => n3789, B2 
                           => n476, ZN => n3803);
   U3680 : NOR3_X1 port map( A1 => n3803, A2 => n3836, A3 => n3790, ZN => n3791
                           );
   U3681 : AOI21_X1 port map( B1 => n3814, B2 => n3856, A => n3791, ZN => n3794
                           );
   U3682 : NOR3_X1 port map( A1 => IR_CU_1_port, A2 => n478, A3 => n3802, ZN =>
                           n3832);
   U3683 : NOR2_X1 port map( A1 => n516, A2 => n510, ZN => n3974);
   U3684 : NAND2_X1 port map( A1 => n3976, A2 => n3974, ZN => n3828);
   U3685 : AOI211_X1 port map( C1 => n3832, C2 => n476, A => n3792, B => n3807,
                           ZN => n3793);
   U3686 : OAI211_X1 port map( C1 => n514, C2 => n3954, A => n3794, B => n3793,
                           ZN => CU_I_aluOpcode_i_1_port);
   U3687 : INV_X1 port map( A => n3966, ZN => n3849);
   U3688 : NOR3_X1 port map( A1 => n3795, A2 => n3955, A3 => n3849, ZN => n3820
                           );
   U3689 : NOR3_X1 port map( A1 => n3795, A2 => n3837, A3 => n3977, ZN => n3831
                           );
   U3690 : INV_X1 port map( A => n3796, ZN => n3799);
   U3691 : INV_X1 port map( A => n3797, ZN => n3970);
   U3692 : OAI21_X1 port map( B1 => n3799, B2 => n3970, A => n3798, ZN => n3800
                           );
   U3693 : NOR4_X1 port map( A1 => n3820, A2 => n3831, A3 => n3801, A4 => n3800
                           , ZN => n3812);
   U3694 : NOR3_X1 port map( A1 => n3803, A2 => n3802, A3 => n480, ZN => n3810)
                           ;
   U3695 : NAND3_X1 port map( A1 => n478, A2 => n3824, A3 => n476, ZN => n3835)
                           ;
   U3696 : NAND2_X1 port map( A1 => n3804, A2 => IR_CU_0_port, ZN => n3805);
   U3697 : AOI211_X1 port map( C1 => n3835, C2 => n3805, A => IR_CU_1_port, B 
                           => n3836, ZN => n3809);
   U3698 : NOR3_X1 port map( A1 => IR_CU_4_port, A2 => n477, A3 => n3806, ZN =>
                           n3808);
   U3699 : NOR4_X1 port map( A1 => n3810, A2 => n3809, A3 => n3808, A4 => n3807
                           , ZN => n3811);
   U3700 : OAI211_X1 port map( C1 => n504, C2 => n3813, A => n3812, B => n3811,
                           ZN => CU_I_aluOpcode_i_2_port);
   U3701 : AOI211_X1 port map( C1 => IR_CU_31, C2 => n510, A => n3977, B => 
                           n3970, ZN => n3819);
   U3702 : NAND2_X1 port map( A1 => n3856, A2 => n3814, ZN => n3816);
   U3703 : NAND2_X1 port map( A1 => n606, A2 => n504, ZN => n3815);
   U3704 : OAI211_X1 port map( C1 => n3849, C2 => n3817, A => n3816, B => n3815
                           , ZN => n3818);
   U3705 : NOR4_X1 port map( A1 => n3821, A2 => n3820, A3 => n3819, A4 => n3818
                           , ZN => n3826);
   U3706 : OAI211_X1 port map( C1 => n2128, C2 => n480, A => IR_CU_5_port, B =>
                           IR_CU_0_port, ZN => n3822);
   U3707 : OAI21_X1 port map( B1 => n478, B2 => n3836, A => n3822, ZN => n3823)
                           ;
   U3708 : NAND3_X1 port map( A1 => n3824, A2 => n477, A3 => n3823, ZN => n3825
                           );
   U3709 : OAI211_X1 port map( C1 => n476, C2 => n3827, A => n3826, B => n3825,
                           ZN => CU_I_aluOpcode_i_3_port);
   U3710 : OAI211_X1 port map( C1 => n516, C2 => n2141, A => n510, B => n2129, 
                           ZN => n3829);
   U3711 : AOI22_X1 port map( A1 => IR_CU_27, A2 => n3829, B1 => n3828, B2 => 
                           n504, ZN => n3830);
   U3712 : AOI211_X1 port map( C1 => n3832, C2 => IR_CU_4_port, A => n3831, B 
                           => n3830, ZN => n3834);
   U3713 : OAI211_X1 port map( C1 => n3836, C2 => n3835, A => n3834, B => n3833
                           , ZN => CU_I_aluOpcode_i_4_port);
   U3714 : OAI211_X1 port map( C1 => IR_CU_26, C2 => n2129, A => IR_CU_28, B =>
                           IR_CU_27, ZN => n3839);
   U3715 : NOR3_X1 port map( A1 => n515, A2 => n510, A3 => n3837, ZN => n3838);
   U3716 : AOI21_X1 port map( B1 => n2141, B2 => n3839, A => n3838, ZN => n3857
                           );
   U3717 : NOR3_X1 port map( A1 => n515, A2 => n2141, A3 => n504, ZN => n3859);
   U3718 : INV_X1 port map( A => n3845, ZN => n3840);
   U3719 : AOI22_X1 port map( A1 => IR_CU_28, A2 => n3859, B1 => n3856, B2 => 
                           n3840, ZN => n3841);
   U3720 : AOI22_X1 port map( A1 => IR_CU_28, A2 => IR_CU_27, B1 => n504, B2 =>
                           n510, ZN => n3844);
   U3721 : NAND2_X1 port map( A1 => n3976, A2 => n3844, ZN => n3860);
   U3722 : OAI221_X1 port map( B1 => IR_CU_31, B2 => n3857, C1 => IR_CU_31, C2 
                           => n3841, A => n3860, ZN => n3846);
   U3723 : AOI21_X1 port map( B1 => n3968, B2 => n3966, A => n3846, ZN => n1371
                           );
   U3724 : AOI21_X1 port map( B1 => IR_CU_26, B2 => n510, A => n504, ZN => 
                           n3843);
   U3725 : INV_X1 port map( A => n3955, ZN => n3973);
   U3726 : NAND2_X1 port map( A1 => IR_CU_31, A2 => n3973, ZN => n3842);
   U3727 : OAI21_X1 port map( B1 => n3843, B2 => n3842, A => n1371, ZN => 
                           CU_I_cw_0_port);
   U3728 : AND3_X1 port map( A1 => n3973, A2 => n3844, A3 => n516, ZN => 
                           CU_I_cw_10_port);
   U3729 : NOR2_X1 port map( A1 => n516, A2 => n3845, ZN => n3850);
   U3730 : AOI21_X1 port map( B1 => n3951, B2 => n3850, A => n3847, ZN => n3862
                           );
   U3731 : INV_X1 port map( A => n3862, ZN => CU_I_cw_6_port);
   U3732 : OR2_X1 port map( A1 => n3846, A2 => CU_I_cw_6_port, ZN => 
                           CU_I_cw_1_port);
   U3733 : NAND2_X1 port map( A1 => n3850, A2 => n2141, ZN => n3852);
   U3734 : AOI22_X1 port map( A1 => n3850, A2 => n3856, B1 => n3847, B2 => n510
                           , ZN => n3848);
   U3735 : OAI21_X1 port map( B1 => n3849, B2 => n3852, A => n3848, ZN => 
                           CU_I_cw_3_port);
   U3736 : NAND2_X1 port map( A1 => n3973, A2 => n3974, ZN => n3854);
   U3737 : OAI211_X1 port map( C1 => n2141, C2 => n497, A => n3850, B => n504, 
                           ZN => n3851);
   U3738 : OAI21_X1 port map( B1 => n3970, B2 => n3854, A => n3851, ZN => 
                           CU_I_cw_4_port);
   U3739 : INV_X1 port map( A => n3854, ZN => n3855);
   U3740 : AOI21_X1 port map( B1 => n3856, B2 => n3855, A => CU_I_cw_7_port, ZN
                           => n1357);
   U3741 : INV_X1 port map( A => n3857, ZN => n3858);
   U3742 : AOI221_X1 port map( B1 => n3859, B2 => n516, C1 => n3858, C2 => n516
                           , A => CU_I_cw_10_port, ZN => n3861);
   U3743 : NAND3_X1 port map( A1 => n3862, A2 => n3861, A3 => n3860, ZN => 
                           CU_I_cw_9_port);
   U3744 : NAND3_X1 port map( A1 => n443, A2 => ALU_OPCODE_i_2_port, A3 => 
                           ALU_OPCODE_i_1_port, ZN => n3903);
   U3745 : OR2_X1 port map( A1 => n3903, A2 => ALU_OPCODE_i_0_port, ZN => n3984
                           );
   U3746 : NOR4_X1 port map( A1 => DataP_alu_out_W_12_port, A2 => 
                           DataP_alu_out_W_11_port, A3 => 
                           DataP_alu_out_W_10_port, A4 => 
                           DataP_alu_out_W_0_port, ZN => n3866);
   U3747 : NOR4_X1 port map( A1 => DataP_alu_out_W_15_port, A2 => 
                           DataP_alu_out_W_14_port, A3 => 
                           DataP_alu_out_W_13_port, A4 => 
                           DataP_alu_out_W_16_port, ZN => n3865);
   U3748 : NOR4_X1 port map( A1 => DataP_alu_out_W_17_port, A2 => 
                           DataP_alu_out_W_19_port, A3 => 
                           DataP_alu_out_W_18_port, A4 => 
                           DataP_alu_out_W_1_port, ZN => n3864);
   U3749 : NOR4_X1 port map( A1 => DataP_alu_out_W_23_port, A2 => 
                           DataP_alu_out_W_21_port, A3 => 
                           DataP_alu_out_W_20_port, A4 => 
                           DataP_alu_out_W_22_port, ZN => n3863);
   U3750 : NAND4_X1 port map( A1 => n3866, A2 => n3865, A3 => n3864, A4 => 
                           n3863, ZN => n3899);
   U3751 : INV_X1 port map( A => DataP_FWD_MUX_BR_S_0_port, ZN => n3871);
   U3752 : NAND2_X1 port map( A1 => n3871, A2 => DataP_FWD_MUX_BR_S_1_port, ZN 
                           => n3880);
   U3753 : INV_X1 port map( A => n3880, ZN => n3898);
   U3754 : NOR4_X1 port map( A1 => DataP_alu_out_W_27_port, A2 => 
                           DataP_alu_out_W_26_port, A3 => 
                           DataP_alu_out_W_25_port, A4 => 
                           DataP_alu_out_W_24_port, ZN => n3870);
   U3755 : NOR4_X1 port map( A1 => DataP_alu_out_W_30_port, A2 => 
                           DataP_alu_out_W_29_port, A3 => 
                           DataP_alu_out_W_28_port, A4 => 
                           DataP_alu_out_W_2_port, ZN => n3869);
   U3756 : NOR4_X1 port map( A1 => DataP_alu_out_W_31_port, A2 => 
                           DataP_alu_out_W_5_port, A3 => DataP_alu_out_W_4_port
                           , A4 => DataP_alu_out_W_3_port, ZN => n3868);
   U3757 : NOR4_X1 port map( A1 => DataP_alu_out_W_9_port, A2 => 
                           DataP_alu_out_W_8_port, A3 => DataP_alu_out_W_7_port
                           , A4 => DataP_alu_out_W_6_port, ZN => n3867);
   U3758 : NAND4_X1 port map( A1 => n3870, A2 => n3869, A3 => n3868, A4 => 
                           n3867, ZN => n3897);
   U3759 : NOR2_X1 port map( A1 => DataP_FWD_MUX_BR_S_1_port, A2 => n3871, ZN 
                           => n3895);
   U3760 : NOR4_X1 port map( A1 => DataP_A_s_27_port, A2 => DataP_A_s_26_port, 
                           A3 => DataP_A_s_25_port, A4 => DataP_A_s_24_port, ZN
                           => n3875);
   U3761 : NOR4_X1 port map( A1 => DataP_A_s_30_port, A2 => DataP_A_s_29_port, 
                           A3 => DataP_A_s_28_port, A4 => DataP_A_s_2_port, ZN 
                           => n3874);
   U3762 : NOR4_X1 port map( A1 => DataP_A_s_31_port, A2 => DataP_A_s_5_port, 
                           A3 => DataP_A_s_4_port, A4 => DataP_A_s_3_port, ZN 
                           => n3873);
   U3763 : NOR4_X1 port map( A1 => DataP_A_s_9_port, A2 => DataP_A_s_8_port, A3
                           => DataP_A_s_7_port, A4 => DataP_A_s_6_port, ZN => 
                           n3872);
   U3764 : NAND4_X1 port map( A1 => n3875, A2 => n3874, A3 => n3873, A4 => 
                           n3872, ZN => n3882);
   U3765 : NOR4_X1 port map( A1 => DataP_A_s_12_port, A2 => DataP_A_s_11_port, 
                           A3 => DataP_A_s_10_port, A4 => DataP_A_s_0_port, ZN 
                           => n3879);
   U3766 : NOR4_X1 port map( A1 => DataP_A_s_15_port, A2 => DataP_A_s_14_port, 
                           A3 => DataP_A_s_13_port, A4 => DataP_A_s_16_port, ZN
                           => n3878);
   U3767 : NOR4_X1 port map( A1 => DataP_A_s_17_port, A2 => DataP_A_s_19_port, 
                           A3 => DataP_A_s_18_port, A4 => DataP_A_s_1_port, ZN 
                           => n3877);
   U3768 : NOR4_X1 port map( A1 => DataP_A_s_23_port, A2 => DataP_A_s_21_port, 
                           A3 => DataP_A_s_20_port, A4 => DataP_A_s_22_port, ZN
                           => n3876);
   U3769 : NAND4_X1 port map( A1 => n3879, A2 => n3878, A3 => n3877, A4 => 
                           n3876, ZN => n3881);
   U3770 : OAI21_X1 port map( B1 => n3882, B2 => n3881, A => n3880, ZN => n3894
                           );
   U3771 : NOR4_X1 port map( A1 => DRAM_ADDRESS_11_port, A2 => 
                           DRAM_ADDRESS_10_port, A3 => DRAM_ADDRESS_1_port, A4 
                           => DRAM_ADDRESS_0_port, ZN => n3886);
   U3772 : NOR4_X1 port map( A1 => DRAM_ADDRESS_5_port, A2 => 
                           DRAM_ADDRESS_4_port, A3 => DRAM_ADDRESS_3_port, A4 
                           => DRAM_ADDRESS_2_port, ZN => n3885);
   U3773 : NOR4_X1 port map( A1 => DRAM_ADDRESS_9_port, A2 => 
                           DRAM_ADDRESS_8_port, A3 => DRAM_ADDRESS_7_port, A4 
                           => DRAM_ADDRESS_6_port, ZN => n3884);
   U3774 : NOR4_X1 port map( A1 => DataP_alu_out_M_15_port, A2 => 
                           DataP_alu_out_M_14_port, A3 => 
                           DataP_alu_out_M_13_port, A4 => 
                           DataP_alu_out_M_12_port, ZN => n3883);
   U3775 : NAND4_X1 port map( A1 => n3886, A2 => n3885, A3 => n3884, A4 => 
                           n3883, ZN => n3892);
   U3776 : NOR4_X1 port map( A1 => DataP_alu_out_M_16_port, A2 => 
                           DataP_alu_out_M_17_port, A3 => 
                           DataP_alu_out_M_19_port, A4 => 
                           DataP_alu_out_M_18_port, ZN => n3890);
   U3777 : NOR4_X1 port map( A1 => DataP_alu_out_M_23_port, A2 => 
                           DataP_alu_out_M_21_port, A3 => 
                           DataP_alu_out_M_20_port, A4 => 
                           DataP_alu_out_M_22_port, ZN => n3889);
   U3778 : NOR4_X1 port map( A1 => DataP_alu_out_M_27_port, A2 => 
                           DataP_alu_out_M_26_port, A3 => 
                           DataP_alu_out_M_25_port, A4 => 
                           DataP_alu_out_M_24_port, ZN => n3888);
   U3779 : NOR4_X1 port map( A1 => DataP_alu_out_M_31_port, A2 => 
                           DataP_alu_out_M_30_port, A3 => 
                           DataP_alu_out_M_29_port, A4 => 
                           DataP_alu_out_M_28_port, ZN => n3887);
   U3780 : NAND4_X1 port map( A1 => n3890, A2 => n3889, A3 => n3888, A4 => 
                           n3887, ZN => n3891);
   U3781 : OAI21_X1 port map( B1 => n3892, B2 => n3891, A => n3895, ZN => n3893
                           );
   U3782 : OAI21_X1 port map( B1 => n3895, B2 => n3894, A => n3893, ZN => n3896
                           );
   U3783 : AOI221_X1 port map( B1 => n3899, B2 => n3898, C1 => n3897, C2 => 
                           n3898, A => n3896, ZN => n3900);
   U3784 : XNOR2_X1 port map( A => DataP_pr_E, B => n3900, ZN => n3983);
   U3785 : NAND2_X1 port map( A1 => BR_EN_i, A2 => ALU_OPCODE_i_3_port, ZN => 
                           n3982);
   U3786 : NAND2_X1 port map( A1 => ALU_OPCODE_i_1_port, A2 => 
                           ALU_OPCODE_i_0_port, ZN => n3902);
   U3787 : INV_X1 port map( A => DataP_npc_8_port, ZN => n3998);
   U3788 : INV_X1 port map( A => DataP_npc_9_port, ZN => n3999);
   U3789 : OAI22_X1 port map( A1 => n341, A2 => n3911, B1 => n3910, B2 => n3999
                           , ZN => DataP_PC_reg_N11);
   U3790 : INV_X1 port map( A => DataP_npc_10_port, ZN => n4000);
   U3791 : OAI22_X1 port map( A1 => n340, A2 => n3911, B1 => n3910, B2 => n4000
                           , ZN => DataP_PC_reg_N12);
   U3792 : INV_X1 port map( A => DataP_npc_11_port, ZN => n4001);
   U3793 : OAI22_X1 port map( A1 => n2137, A2 => n3911, B1 => n3910, B2 => 
                           n4001, ZN => DataP_PC_reg_N13);
   U3794 : INV_X1 port map( A => DataP_npc_12_port, ZN => n4002);
   U3795 : OAI22_X1 port map( A1 => n337, A2 => n3911, B1 => n3910, B2 => n4002
                           , ZN => DataP_PC_reg_N14);
   U3796 : NAND3_X1 port map( A1 => n2222, A2 => n3907, A3 => n3906, ZN => 
                           n3905);
   U3797 : INV_X1 port map( A => DataP_npc_0_port, ZN => n3990);
   U3798 : INV_X1 port map( A => DataP_npc_1_port, ZN => n3991);
   U3799 : OAI22_X1 port map( A1 => n358, A2 => n3911, B1 => n3910, B2 => n3991
                           , ZN => DataP_PC_reg_N3);
   U3800 : INV_X1 port map( A => DataP_npc_2_port, ZN => n3992);
   U3801 : OAI22_X1 port map( A1 => n357, A2 => n3911, B1 => n3910, B2 => n3992
                           , ZN => DataP_PC_reg_N4);
   U3802 : INV_X1 port map( A => DataP_npc_3_port, ZN => n3993);
   U3803 : INV_X1 port map( A => DataP_npc_4_port, ZN => n3994);
   U3804 : INV_X1 port map( A => DataP_npc_5_port, ZN => n3995);
   U3805 : OAI22_X1 port map( A1 => n354, A2 => n3911, B1 => n3910, B2 => n3995
                           , ZN => DataP_PC_reg_N7);
   U3806 : INV_X1 port map( A => DataP_npc_6_port, ZN => n3996);
   U3807 : INV_X1 port map( A => DataP_npc_7_port, ZN => n3997);
   U3808 : OAI22_X1 port map( A1 => n350, A2 => n3911, B1 => n3910, B2 => n3997
                           , ZN => DataP_PC_reg_N9);
   U3809 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_0_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_0_port, ZN => n3912);
   U3810 : OAI21_X1 port map( B1 => n2272, B2 => n3946, A => n3912, ZN => 
                           DataP_WB_0_port);
   U3811 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_10_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_10_port, ZN => n3913)
                           ;
   U3812 : OAI21_X1 port map( B1 => n2257, B2 => n3946, A => n3913, ZN => 
                           DataP_WB_10_port);
   U3813 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_11_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_11_port, ZN => n3914)
                           ;
   U3814 : OAI21_X1 port map( B1 => n2251, B2 => n3946, A => n3914, ZN => 
                           DataP_WB_11_port);
   U3815 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_12_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_12_port, ZN => n3915)
                           ;
   U3816 : OAI21_X1 port map( B1 => n2246, B2 => n3946, A => n3915, ZN => 
                           DataP_WB_12_port);
   U3817 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_13_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_13_port, ZN => n3916)
                           ;
   U3818 : OAI21_X1 port map( B1 => n2258, B2 => n3946, A => n3916, ZN => 
                           DataP_WB_13_port);
   U3819 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_14_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_14_port, ZN => n3917)
                           ;
   U3820 : OAI21_X1 port map( B1 => n2252, B2 => n3946, A => n3917, ZN => 
                           DataP_WB_14_port);
   U3821 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_15_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_15_port, ZN => n3918)
                           ;
   U3822 : OAI21_X1 port map( B1 => n2247, B2 => n3946, A => n3918, ZN => 
                           DataP_WB_15_port);
   U3823 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_16_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_16_port, ZN => n3919)
                           ;
   U3824 : OAI21_X1 port map( B1 => n2263, B2 => n3946, A => n3919, ZN => 
                           DataP_WB_16_port);
   U3825 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_17_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_17_port, ZN => n3920)
                           ;
   U3826 : OAI21_X1 port map( B1 => n2248, B2 => n3946, A => n3920, ZN => 
                           DataP_WB_17_port);
   U3827 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_18_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_18_port, ZN => n3921)
                           ;
   U3828 : OAI21_X1 port map( B1 => n2259, B2 => n3946, A => n3921, ZN => 
                           DataP_WB_18_port);
   U3829 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_19_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_19_port, ZN => n3922)
                           ;
   U3830 : OAI21_X1 port map( B1 => n2253, B2 => n3946, A => n3922, ZN => 
                           DataP_WB_19_port);
   U3831 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_1_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_1_port, ZN => n3923);
   U3832 : OAI21_X1 port map( B1 => n2273, B2 => n3946, A => n3923, ZN => 
                           DataP_WB_1_port);
   U3833 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_20_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_20_port, ZN => n3924)
                           ;
   U3834 : OAI21_X1 port map( B1 => n2260, B2 => n3946, A => n3924, ZN => 
                           DataP_WB_20_port);
   U3835 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_21_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_21_port, ZN => n3925)
                           ;
   U3836 : OAI21_X1 port map( B1 => n2254, B2 => n3946, A => n3925, ZN => 
                           DataP_WB_21_port);
   U3837 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_22_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_22_port, ZN => n3926)
                           ;
   U3838 : OAI21_X1 port map( B1 => n2264, B2 => n3946, A => n3926, ZN => 
                           DataP_WB_22_port);
   U3839 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_23_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_23_port, ZN => n3927)
                           ;
   U3840 : OAI21_X1 port map( B1 => n2249, B2 => n3946, A => n3927, ZN => 
                           DataP_WB_23_port);
   U3841 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_24_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_24_port, ZN => n3928)
                           ;
   U3842 : OAI21_X1 port map( B1 => n2265, B2 => n3946, A => n3928, ZN => 
                           DataP_WB_24_port);
   U3843 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_25_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_25_port, ZN => n3929)
                           ;
   U3844 : OAI21_X1 port map( B1 => n2261, B2 => n3946, A => n3929, ZN => 
                           DataP_WB_25_port);
   U3845 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_26_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_26_port, ZN => n3930)
                           ;
   U3846 : OAI21_X1 port map( B1 => n2255, B2 => n3946, A => n3930, ZN => 
                           DataP_WB_26_port);
   U3847 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_27_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_27_port, ZN => n3931)
                           ;
   U3848 : OAI21_X1 port map( B1 => n2250, B2 => n3946, A => n3931, ZN => 
                           DataP_WB_27_port);
   U3849 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_28_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_28_port, ZN => n3932)
                           ;
   U3850 : OAI21_X1 port map( B1 => n2262, B2 => n3946, A => n3932, ZN => 
                           DataP_WB_28_port);
   U3851 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_29_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_29_port, ZN => n3933)
                           ;
   U3852 : OAI21_X1 port map( B1 => n2256, B2 => n3946, A => n3933, ZN => 
                           DataP_WB_29_port);
   U3853 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_2_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_2_port, ZN => n3934);
   U3854 : OAI21_X1 port map( B1 => n2276, B2 => n3946, A => n3934, ZN => 
                           DataP_WB_2_port);
   U3855 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_30_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_30_port, ZN => n3935)
                           ;
   U3856 : OAI21_X1 port map( B1 => n2266, B2 => n3946, A => n3935, ZN => 
                           DataP_WB_30_port);
   U3857 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_31_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_31_port, ZN => n3936)
                           ;
   U3858 : OAI21_X1 port map( B1 => n2267, B2 => n3946, A => n3936, ZN => 
                           DataP_WB_31_port);
   U3859 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_3_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_3_port, ZN => n3937);
   U3860 : OAI21_X1 port map( B1 => n2277, B2 => n3946, A => n3937, ZN => 
                           DataP_WB_3_port);
   U3861 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_4_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_4_port, ZN => n3938);
   U3862 : OAI21_X1 port map( B1 => n2274, B2 => n3946, A => n3938, ZN => 
                           DataP_WB_4_port);
   U3863 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_5_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_5_port, ZN => n3939);
   U3864 : OAI21_X1 port map( B1 => n2270, B2 => n3946, A => n3939, ZN => 
                           DataP_WB_5_port);
   U3865 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_6_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_6_port, ZN => n3940);
   U3866 : OAI21_X1 port map( B1 => n2268, B2 => n3946, A => n3940, ZN => 
                           DataP_WB_6_port);
   U3867 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_7_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_7_port, ZN => n3941);
   U3868 : OAI21_X1 port map( B1 => n2275, B2 => n3946, A => n3941, ZN => 
                           DataP_WB_7_port);
   U3869 : AOI22_X1 port map( A1 => n3944, A2 => DataP_LMD_out_8_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_8_port, ZN => n3942);
   U3870 : OAI21_X1 port map( B1 => n2271, B2 => n3946, A => n3942, ZN => 
                           DataP_WB_8_port);
   U3871 : AOI22_X1 port map( A1 => n3008, A2 => DataP_LMD_out_9_port, B1 => 
                           n3943, B2 => DataP_link_addr_W_9_port, ZN => n3945);
   U3872 : OAI21_X1 port map( B1 => n2269, B2 => n3946, A => n3945, ZN => 
                           DataP_WB_9_port);
   U3873 : INV_X1 port map( A => n144, ZN => n3952);
   U3874 : AOI211_X1 port map( C1 => n606, C2 => n504, A => CU_I_cw_7_port, B 
                           => n3953, ZN => n3950);
   U3875 : OAI211_X1 port map( C1 => n3952, C2 => n3951, A => Rst, B => n3950, 
                           ZN => n3964);
   U3876 : AND2_X1 port map( A1 => Rst, A2 => n3953, ZN => n3962);
   U3877 : NOR2_X1 port map( A1 => n3955, A2 => n3954, ZN => n3965);
   U3878 : NAND2_X1 port map( A1 => Rst, A2 => n3965, ZN => n3979);
   U3879 : OAI22_X1 port map( A1 => n497, A2 => n3979, B1 => n3956, B2 => n3964
                           , ZN => n3961);
   U3880 : AOI21_X1 port map( B1 => n3962, B2 => DataP_IR1_11_port, A => n3961,
                           ZN => n3957);
   U3881 : OAI21_X1 port map( B1 => n485, B2 => n3964, A => n3957, ZN => 
                           DataP_dest_D_0_port);
   U3882 : AOI21_X1 port map( B1 => n3962, B2 => DataP_IR1_12_port, A => n3961,
                           ZN => n3958);
   U3883 : OAI21_X1 port map( B1 => n486, B2 => n3964, A => n3958, ZN => 
                           DataP_dest_D_1_port);
   U3884 : AOI21_X1 port map( B1 => n3962, B2 => DataP_IR1_13_port, A => n3961,
                           ZN => n3959);
   U3885 : OAI21_X1 port map( B1 => n487, B2 => n3964, A => n3959, ZN => 
                           DataP_dest_D_2_port);
   U3886 : AOI21_X1 port map( B1 => n3962, B2 => DataP_IR1_14_port, A => n3961,
                           ZN => n3960);
   U3887 : OAI21_X1 port map( B1 => n488, B2 => n3964, A => n3960, ZN => 
                           DataP_dest_D_3_port);
   U3888 : AOI21_X1 port map( B1 => n3962, B2 => DataP_IR1_15_port, A => n3961,
                           ZN => n3963);
   U3889 : OAI21_X1 port map( B1 => n489, B2 => n3964, A => n3963, ZN => 
                           DataP_dest_D_4_port);
   U3890 : NAND2_X1 port map( A1 => IR_CU_28, A2 => n3966, ZN => n3971);
   U3891 : OAI21_X1 port map( B1 => n515, B2 => IR_CU_27, A => n2141, ZN => 
                           n3967);
   U3892 : AOI22_X1 port map( A1 => n3968, A2 => n497, B1 => n510, B2 => n3967,
                           ZN => n3969);
   U3893 : OAI221_X1 port map( B1 => n514, B2 => n3971, C1 => n2141, C2 => 
                           n3970, A => n3969, ZN => n3972);
   U3894 : AOI211_X1 port map( C1 => IR_CU_27, C2 => n3974, A => n3973, B => 
                           n3972, ZN => n3975);
   U3895 : OAI221_X1 port map( B1 => IR_CU_31, B2 => n3977, C1 => n516, C2 => 
                           n3976, A => n3975, ZN => n3978);
   U3896 : NAND4_X1 port map( A1 => Rst, A2 => DataP_IR1_15_port, A3 => n3981, 
                           A4 => n3978, ZN => n3980);
   U3897 : OAI21_X1 port map( B1 => n485, B2 => n3979, A => n3980, ZN => 
                           DataP_imm_out_16_port);
   U3898 : OAI21_X1 port map( B1 => n486, B2 => n3979, A => n3980, ZN => 
                           DataP_imm_out_17_port);
   U3899 : OAI21_X1 port map( B1 => n487, B2 => n3979, A => n3980, ZN => 
                           DataP_imm_out_18_port);
   U3900 : OAI21_X1 port map( B1 => n488, B2 => n3979, A => n3980, ZN => 
                           DataP_imm_out_19_port);
   U3901 : OAI21_X1 port map( B1 => n489, B2 => n3979, A => n3980, ZN => 
                           DataP_imm_out_20_port);
   U3902 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_21_port, ZN => n3989);
   U3903 : OAI21_X1 port map( B1 => n3981, B2 => n3989, A => n3980, ZN => 
                           DataP_imm_out_21_port);
   U3904 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_22_port, ZN => n3988);
   U3905 : OAI21_X1 port map( B1 => n3981, B2 => n3988, A => n3980, ZN => 
                           DataP_imm_out_22_port);
   U3906 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_23_port, ZN => n3987);
   U3907 : OAI21_X1 port map( B1 => n3981, B2 => n3987, A => n3980, ZN => 
                           DataP_imm_out_23_port);
   U3908 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_24_port, ZN => n3986);
   U3909 : OAI21_X1 port map( B1 => n3981, B2 => n3986, A => n3980, ZN => 
                           DataP_imm_out_24_port);
   U3910 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_25_port, ZN => n3985);
   U3911 : OAI21_X1 port map( B1 => n3981, B2 => n3985, A => n3980, ZN => 
                           DataP_imm_out_31_port);
   U3912 : MUX2_X1 port map( A => DataP_pc_out_0, B => DataP_npc_pre_0_port, S 
                           => n1940, Z => DataP_NPC_add_N1);
   U3913 : MUX2_X1 port map( A => DataP_pc_out_1, B => DataP_npc_pre_1_port, S 
                           => n1940, Z => DataP_NPC_add_N2);
   U3914 : NAND2_X1 port map( A1 => DataP_npc_0_port, A2 => n3009, ZN => n127);
   U3915 : AOI21_X1 port map( B1 => n3990, B2 => n4022, A => n3013, ZN => n126)
                           ;
   U3916 : NAND2_X1 port map( A1 => DataP_npc_1_port, A2 => n4021, ZN => n123);
   U3917 : AOI21_X1 port map( B1 => n3991, B2 => n4022, A => n3013, ZN => n122)
                           ;
   U3918 : NAND2_X1 port map( A1 => DataP_npc_2_port, A2 => n3009, ZN => n119);
   U3919 : AOI21_X1 port map( B1 => n3992, B2 => n4022, A => n3013, ZN => n118)
                           ;
   U3920 : NAND2_X1 port map( A1 => DataP_npc_3_port, A2 => n4021, ZN => n115);
   U3921 : AOI21_X1 port map( B1 => n3993, B2 => n4022, A => n3013, ZN => n114)
                           ;
   U3922 : NAND2_X1 port map( A1 => DataP_npc_4_port, A2 => n3009, ZN => n111);
   U3923 : AOI21_X1 port map( B1 => n3994, B2 => n4022, A => n3013, ZN => n110)
                           ;
   U3924 : NAND2_X1 port map( A1 => DataP_npc_5_port, A2 => n4021, ZN => n107);
   U3925 : AOI21_X1 port map( B1 => n3995, B2 => n4022, A => n3013, ZN => n106)
                           ;
   U3926 : NAND2_X1 port map( A1 => DataP_npc_6_port, A2 => n4021, ZN => n103);
   U3927 : AOI21_X1 port map( B1 => n3996, B2 => n4022, A => n3013, ZN => n102)
                           ;
   U3928 : NAND2_X1 port map( A1 => DataP_npc_7_port, A2 => n4021, ZN => n99);
   U3929 : AOI21_X1 port map( B1 => n3997, B2 => n4022, A => n3013, ZN => n98);
   U3930 : NAND2_X1 port map( A1 => DataP_npc_8_port, A2 => n4021, ZN => n95);
   U3931 : AOI21_X1 port map( B1 => n3998, B2 => n4022, A => n3013, ZN => n94);
   U3932 : NAND2_X1 port map( A1 => DataP_npc_9_port, A2 => n4021, ZN => n91);
   U3933 : AOI21_X1 port map( B1 => n3999, B2 => n4022, A => n3013, ZN => n90);
   U3934 : NAND2_X1 port map( A1 => DataP_npc_10_port, A2 => n4021, ZN => n87);
   U3935 : AOI21_X1 port map( B1 => n4000, B2 => n4022, A => n3014, ZN => n86);
   U3936 : NAND2_X1 port map( A1 => DataP_npc_11_port, A2 => n4021, ZN => n83);
   U3937 : AOI21_X1 port map( B1 => n4001, B2 => n4022, A => n3013, ZN => n82);
   U3938 : NAND2_X1 port map( A1 => DataP_npc_12_port, A2 => n3009, ZN => n79);
   U3939 : AOI21_X1 port map( B1 => n4002, B2 => n4022, A => n3013, ZN => n78);
   U3940 : NAND2_X1 port map( A1 => DataP_npc_13_port, A2 => n3009, ZN => n75);
   U3941 : AOI21_X1 port map( B1 => n4003, B2 => n4022, A => n3013, ZN => n74);
   U3942 : NAND2_X1 port map( A1 => DataP_npc_14_port, A2 => n3009, ZN => n71);
   U3943 : AOI21_X1 port map( B1 => n4004, B2 => n4022, A => n3013, ZN => n70);
   U3944 : NAND2_X1 port map( A1 => DataP_npc_15_port, A2 => n3009, ZN => n67);
   U3945 : AOI21_X1 port map( B1 => n4005, B2 => n4022, A => n3014, ZN => n66);
   U3946 : NAND2_X1 port map( A1 => DataP_npc_16_port, A2 => n3009, ZN => n63);
   U3947 : AOI21_X1 port map( B1 => n4006, B2 => n4022, A => n3014, ZN => n62);
   U3948 : NAND2_X1 port map( A1 => DataP_npc_17_port, A2 => n3009, ZN => n59);
   U3949 : AOI21_X1 port map( B1 => n4007, B2 => n4022, A => n3014, ZN => n58);
   U3950 : NAND2_X1 port map( A1 => DataP_npc_18_port, A2 => n3009, ZN => n55);
   U3951 : AOI21_X1 port map( B1 => n4008, B2 => n4022, A => n3014, ZN => n54);
   U3952 : NAND2_X1 port map( A1 => DataP_npc_19_port, A2 => n3009, ZN => n51);
   U3953 : AOI21_X1 port map( B1 => n4009, B2 => n4022, A => n3014, ZN => n50);
   U3954 : NAND2_X1 port map( A1 => DataP_npc_20_port, A2 => n3009, ZN => n47);
   U3955 : AOI21_X1 port map( B1 => n4010, B2 => n4022, A => n3014, ZN => n46);
   U3956 : NAND2_X1 port map( A1 => DataP_npc_21_port, A2 => n3009, ZN => n43);
   U3957 : AOI21_X1 port map( B1 => n4011, B2 => n4022, A => n3014, ZN => n42);
   U3958 : NAND2_X1 port map( A1 => DataP_npc_22_port, A2 => n4021, ZN => n39);
   U3959 : AOI21_X1 port map( B1 => n4012, B2 => n4022, A => n3014, ZN => n38);
   U3960 : NAND2_X1 port map( A1 => DataP_npc_23_port, A2 => n4021, ZN => n35);
   U3961 : AOI21_X1 port map( B1 => n4013, B2 => n4022, A => n3014, ZN => n34);
   U3962 : NAND2_X1 port map( A1 => DataP_npc_24_port, A2 => n3009, ZN => n31);
   U3963 : AOI21_X1 port map( B1 => n4014, B2 => n4022, A => n3014, ZN => n30);
   U3964 : NAND2_X1 port map( A1 => DataP_npc_25_port, A2 => n3009, ZN => n27);
   U3965 : AOI21_X1 port map( B1 => n4015, B2 => n4022, A => n3014, ZN => n26);
   U3966 : NAND2_X1 port map( A1 => DataP_npc_26_port, A2 => n3009, ZN => n23);
   U3967 : AOI21_X1 port map( B1 => n4016, B2 => n4022, A => n3014, ZN => n22);
   U3968 : NAND2_X1 port map( A1 => DataP_npc_27_port, A2 => n3009, ZN => n19);
   U3969 : AOI21_X1 port map( B1 => n4017, B2 => n4022, A => n3014, ZN => n18);
   U3970 : NAND2_X1 port map( A1 => DataP_npc_28_port, A2 => n3009, ZN => n15);
   U3971 : AOI21_X1 port map( B1 => n4018, B2 => n4022, A => n3014, ZN => n14);
   U3972 : NAND2_X1 port map( A1 => DataP_npc_29_port, A2 => n3009, ZN => n11);
   U3973 : AOI21_X1 port map( B1 => n4019, B2 => n4022, A => n3014, ZN => n10);
   U3974 : NAND2_X1 port map( A1 => DataP_npc_30_port, A2 => n3009, ZN => n7);
   U3975 : AOI21_X1 port map( B1 => n4020, B2 => n4022, A => n3014, ZN => n6);
   U3976 : NAND2_X1 port map( A1 => DataP_npc_31_port, A2 => n3009, ZN => n3);
   U3977 : AOI21_X1 port map( B1 => n4023, B2 => n4022, A => n3013, ZN => n2);

end SYN_structural;
