
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_syn is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, ADDS, SUBS, ANDS, ORS, XORS, LLS, LRS, SNE, SGE, SLE, J, 
   JAL, BEQZ, BNEZ, RAS, JR, JALR, SLT, SGT, SEQ, SLTU, SLEU, SGTU, SGEU);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111 11000";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX_syn;

package body CONV_PACK_DLX_syn is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return ADDS;
         when "00010" => return SUBS;
         when "00011" => return ANDS;
         when "00100" => return ORS;
         when "00101" => return XORS;
         when "00110" => return LLS;
         when "00111" => return LRS;
         when "01000" => return SNE;
         when "01001" => return SGE;
         when "01010" => return SLE;
         when "01011" => return J;
         when "01100" => return JAL;
         when "01101" => return BEQZ;
         when "01110" => return BNEZ;
         when "01111" => return RAS;
         when "10000" => return JR;
         when "10001" => return JALR;
         when "10010" => return SLT;
         when "10011" => return SGT;
         when "10100" => return SEQ;
         when "10101" => return SLTU;
         when "10110" => return SLEU;
         when "10111" => return SGTU;
         when "11000" => return SGEU;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when ADDS => return "00001";
         when SUBS => return "00010";
         when ANDS => return "00011";
         when ORS => return "00100";
         when XORS => return "00101";
         when LLS => return "00110";
         when LRS => return "00111";
         when SNE => return "01000";
         when SGE => return "01001";
         when SLE => return "01010";
         when J => return "01011";
         when JAL => return "01100";
         when BEQZ => return "01101";
         when BNEZ => return "01110";
         when RAS => return "01111";
         when JR => return "10000";
         when JALR => return "10001";
         when SLT => return "10010";
         when SGT => return "10011";
         when SEQ => return "10100";
         when SLTU => return "10101";
         when SLEU => return "10110";
         when SGTU => return "10111";
         when SGEU => return "11000";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_DLX_syn;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity add_sub_N32_DW01_sub_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end add_sub_N32_DW01_sub_2;

architecture SYN_cla of add_sub_N32_DW01_sub_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, DIFF_2_port, 
      DIFF_1_port, net26789, net26755, net26754, net26748, net37260, net37319, 
      net37512, net37522, net37543, net37600, net37602, net37633, net37685, 
      net37702, net37708, net37710, net37712, net37722, net37727, net37752, 
      net37871, net37882, net37954, net37922, net37353, net37243, net36877, 
      net26708, net26701, net36876, net26750, net39045, net37930, net37768, 
      net37416, net26732, net26707, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, DIFF_0_port, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_0_port );
   
   U3 : OR2_X1 port map( A1 => n10, A2 => n1, ZN => n89);
   U4 : NAND2_X1 port map( A1 => n2, A2 => net37319, ZN => n1);
   U5 : NOR2_X1 port map( A1 => net37602, A2 => net37712, ZN => n2);
   U6 : INV_X1 port map( A => n28, ZN => n3);
   U7 : INV_X1 port map( A => n3, ZN => n4);
   U8 : INV_X1 port map( A => n25, ZN => n5);
   U9 : CLKBUF_X1 port map( A => net37602, Z => n6);
   U10 : NOR2_X1 port map( A1 => n84, A2 => n85, ZN => n7);
   U11 : AND2_X1 port map( A1 => n37, A2 => n81, ZN => n8);
   U12 : XNOR2_X1 port map( A => net37543, B => n9, ZN => DIFF_6_port);
   U13 : NAND2_X1 port map( A1 => n64, A2 => net37512, ZN => n9);
   U14 : OR2_X1 port map( A1 => n88, A2 => net26748, ZN => n10);
   U15 : BUF_X1 port map( A => n33, Z => net37722);
   U16 : XNOR2_X1 port map( A => n11, B => net37954, ZN => DIFF_11_port);
   U17 : NOR2_X1 port map( A1 => n60, A2 => n43, ZN => n11);
   U18 : CLKBUF_X1 port map( A => net37243, Z => net37416);
   U19 : AND4_X2 port map( A1 => n71, A2 => n67, A3 => n70, A4 => n50, ZN => 
                           n53);
   U20 : XNOR2_X1 port map( A => n12, B => n81, ZN => DIFF_26_port);
   U21 : NAND2_X1 port map( A1 => n46, A2 => n37, ZN => n12);
   U22 : AND2_X1 port map( A1 => net37243, A2 => n13, ZN => n17);
   U23 : AND2_X1 port map( A1 => net39045, A2 => n18, ZN => n13);
   U24 : NOR2_X1 port map( A1 => net26707, A2 => net26708, ZN => n14);
   U25 : XNOR2_X1 port map( A => n14, B => B(20), ZN => DIFF_20_port);
   U26 : INV_X1 port map( A => net37768, ZN => net26707);
   U27 : NOR2_X1 port map( A1 => net37930, A2 => net26708, ZN => net37260);
   U28 : INV_X1 port map( A => B(17), ZN => n16);
   U29 : AND2_X1 port map( A1 => n16, A2 => n19, ZN => n18);
   U30 : NAND3_X1 port map( A1 => n19, A2 => n15, A3 => n16, ZN => net26708);
   U31 : INV_X1 port map( A => B(19), ZN => n15);
   U32 : INV_X1 port map( A => B(18), ZN => n19);
   U33 : AND2_X1 port map( A1 => net37600, A2 => net39045, ZN => net37768);
   U34 : CLKBUF_X1 port map( A => net26732, Z => net39045);
   U35 : XOR2_X1 port map( A => net37416, B => net39045, Z => DIFF_16_port);
   U36 : AND2_X1 port map( A1 => net37600, A2 => net39045, ZN => net37353);
   U37 : INV_X1 port map( A => B(16), ZN => net26732);
   U38 : NAND2_X1 port map( A1 => net26732, A2 => net26701, ZN => net37930);
   U39 : AND2_X1 port map( A1 => net26732, A2 => net37882, ZN => net37752);
   U40 : XNOR2_X1 port map( A => n17, B => B(19), ZN => DIFF_19_port);
   U41 : CLKBUF_X1 port map( A => B(18), Z => net37922);
   U42 : AND2_X1 port map( A1 => net37243, A2 => net37260, ZN => net37727);
   U43 : NOR2_X1 port map( A1 => n21, A2 => net26750, ZN => net36876);
   U44 : AND2_X1 port map( A1 => net36876, A2 => net36877, ZN => net37600);
   U45 : AND2_X1 port map( A1 => net36876, A2 => net36877, ZN => net37243);
   U46 : NAND4_X1 port map( A1 => n24, A2 => n28, A3 => n25, A4 => n20, ZN => 
                           net26750);
   U47 : INV_X1 port map( A => B(8), ZN => n20);
   U48 : NAND4_X1 port map( A1 => n24, A2 => n28, A3 => n25, A4 => n20, ZN => 
                           net37602);
   U49 : INV_X1 port map( A => B(9), ZN => n25);
   U50 : INV_X1 port map( A => B(10), ZN => n28);
   U51 : INV_X1 port map( A => B(11), ZN => n24);
   U52 : NAND4_X1 port map( A1 => n26, A2 => n27, A3 => n22, A4 => n23, ZN => 
                           n21);
   U53 : INV_X1 port map( A => B(13), ZN => n23);
   U54 : CLKBUF_X1 port map( A => n23, Z => net37633);
   U55 : AND2_X1 port map( A1 => n23, A2 => net26754, ZN => net37319);
   U56 : INV_X1 port map( A => B(12), ZN => n22);
   U57 : INV_X1 port map( A => B(15), ZN => n27);
   U58 : INV_X1 port map( A => B(14), ZN => n26);
   U59 : INV_X1 port map( A => B(8), ZN => net37702);
   U60 : CLKBUF_X1 port map( A => B(11), Z => net37954);
   U61 : CLKBUF_X1 port map( A => B(12), Z => net37712);
   U62 : CLKBUF_X1 port map( A => B(15), Z => net37710);
   U63 : CLKBUF_X1 port map( A => B(14), Z => net37708);
   U64 : INV_X1 port map( A => B(20), ZN => net26701);
   U65 : NOR2_X1 port map( A1 => net26708, A2 => B(20), ZN => net37522);
   U66 : OR2_X2 port map( A1 => n30, A2 => n88, ZN => n60);
   U67 : XNOR2_X1 port map( A => n29, B => n87, ZN => DIFF_23_port);
   U68 : NAND2_X1 port map( A1 => net37243, A2 => n49, ZN => n29);
   U69 : XOR2_X1 port map( A => n65, B => n86, Z => DIFF_22_port);
   U70 : NAND4_X1 port map( A1 => net37871, A2 => n32, A3 => n33, A4 => n31, ZN
                           => n30);
   U71 : NOR2_X1 port map( A1 => net37685, A2 => n34, ZN => net36877);
   U72 : NAND4_X1 port map( A1 => net37871, A2 => n32, A3 => n33, A4 => n31, ZN
                           => n34);
   U73 : INV_X1 port map( A => B(6), ZN => n31);
   U74 : NAND4_X1 port map( A1 => net37871, A2 => n32, A3 => n33, A4 => n31, ZN
                           => net26748);
   U75 : CLKBUF_X1 port map( A => n31, Z => net37543);
   U76 : INV_X1 port map( A => B(4), ZN => n33);
   U77 : INV_X1 port map( A => B(5), ZN => n32);
   U78 : CLKBUF_X1 port map( A => n32, Z => net37512);
   U79 : XNOR2_X1 port map( A => n35, B => net37922, ZN => DIFF_18_port);
   U80 : AND2_X1 port map( A1 => net37353, A2 => n16, ZN => n35);
   U81 : INV_X1 port map( A => B(0), ZN => n36);
   U82 : INV_X1 port map( A => B(25), ZN => n37);
   U83 : INV_X1 port map( A => B(3), ZN => n38);
   U84 : XNOR2_X1 port map( A => net37708, B => n90, ZN => DIFF_14_port);
   U85 : OR2_X1 port map( A1 => net37602, A2 => net37712, ZN => n55);
   U86 : AND2_X2 port map( A1 => n53, A2 => net37722, ZN => n64);
   U87 : OR2_X1 port map( A1 => n88, A2 => net26748, ZN => n59);
   U88 : INV_X1 port map( A => DIFF_0_port, ZN => n39);
   U89 : INV_X1 port map( A => n85, ZN => n40);
   U90 : NOR2_X1 port map( A1 => n41, A2 => n84, ZN => n46);
   U91 : NAND2_X1 port map( A1 => n83, A2 => n40, ZN => n41);
   U92 : OR2_X1 port map( A1 => n79, A2 => n42, ZN => n76);
   U93 : OR2_X1 port map( A1 => n80, A2 => B(28), ZN => n42);
   U94 : OR2_X1 port map( A1 => n58, A2 => B(10), ZN => n43);
   U95 : CLKBUF_X1 port map( A => n70, Z => n44);
   U96 : NOR2_X1 port map( A1 => B(21), A2 => B(22), ZN => net37882);
   U97 : INV_X1 port map( A => B(7), ZN => net37871);
   U98 : INV_X1 port map( A => B(21), ZN => n45);
   U99 : OR2_X1 port map( A1 => n47, A2 => n84, ZN => n79);
   U100 : OR2_X1 port map( A1 => n85, A2 => B(24), ZN => n47);
   U101 : NOR2_X1 port map( A1 => n60, A2 => n58, ZN => n92);
   U102 : NOR2_X1 port map( A1 => n6, A2 => n60, ZN => n91);
   U103 : AND2_X1 port map( A1 => net37522, A2 => net37752, ZN => n49);
   U104 : XNOR2_X1 port map( A => n48, B => n5, ZN => DIFF_9_port);
   U105 : NOR2_X1 port map( A1 => n59, A2 => net26789, ZN => n48);
   U106 : NAND4_X1 port map( A1 => n77, A2 => n38, A3 => n36, A4 => n70, ZN => 
                           net37685);
   U107 : INV_X1 port map( A => B(1), ZN => n50);
   U108 : NAND2_X1 port map( A1 => n64, A2 => n51, ZN => n68);
   U109 : AND2_X1 port map( A1 => net37512, A2 => net37543, ZN => n51);
   U110 : XNOR2_X1 port map( A => net37727, B => B(21), ZN => DIFF_21_port);
   U111 : CLKBUF_X1 port map( A => B(0), Z => DIFF_0_port);
   U112 : AND2_X1 port map( A1 => net37727, A2 => n45, ZN => n65);
   U113 : NOR2_X1 port map( A1 => n60, A2 => n55, ZN => n54);
   U114 : NOR2_X1 port map( A1 => n55, A2 => n10, ZN => n63);
   U115 : NOR2_X1 port map( A1 => n84, A2 => n85, ZN => n56);
   U116 : AND2_X1 port map( A1 => n7, A2 => n57, ZN => n66);
   U117 : AND2_X1 port map( A1 => n8, A2 => n83, ZN => n57);
   U118 : AND2_X1 port map( A1 => n63, A2 => net37633, ZN => n90);
   U119 : OR2_X1 port map( A1 => net26789, A2 => B(9), ZN => n58);
   U120 : NAND2_X1 port map( A1 => net37600, A2 => net37260, ZN => n84);
   U121 : XNOR2_X1 port map( A => n89, B => net26755, ZN => DIFF_15_port);
   U122 : INV_X1 port map( A => n60, ZN => n61);
   U123 : XOR2_X1 port map( A => n74, B => n75, Z => DIFF_30_port);
   U124 : NOR2_X1 port map( A1 => B(29), A2 => n76, ZN => n74);
   U125 : NAND4_X1 port map( A1 => n36, A2 => n71, A3 => n50, A4 => n70, ZN => 
                           n88);
   U126 : NOR2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U127 : AND2_X1 port map( A1 => n77, A2 => n67, ZN => n62);
   U128 : NAND2_X1 port map( A1 => n44, A2 => n62, ZN => n69);
   U129 : XOR2_X1 port map( A => net37702, B => n61, Z => DIFF_8_port);
   U130 : XOR2_X1 port map( A => n76, B => B(29), Z => DIFF_29_port);
   U131 : XNOR2_X1 port map( A => n72, B => n73, ZN => DIFF_31_port);
   U132 : INV_X1 port map( A => B(31), ZN => n73);
   U133 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => n72);
   U134 : XNOR2_X1 port map( A => n78, B => B(28), ZN => DIFF_28_port);
   U135 : XNOR2_X1 port map( A => n66, B => B(27), ZN => DIFF_27_port);
   U136 : XOR2_X1 port map( A => n44, B => n62, Z => DIFF_2_port);
   U137 : XOR2_X1 port map( A => net37512, B => n64, Z => DIFF_5_port);
   U138 : XOR2_X1 port map( A => n77, B => n39, Z => DIFF_1_port);
   U139 : INV_X1 port map( A => B(2), ZN => n70);
   U140 : INV_X1 port map( A => net37708, ZN => net26754);
   U141 : XOR2_X1 port map( A => n4, B => n92, Z => DIFF_10_port);
   U142 : INV_X1 port map( A => B(26), ZN => n81);
   U143 : INV_X1 port map( A => B(22), ZN => n86);
   U144 : INV_X1 port map( A => B(3), ZN => n71);
   U145 : INV_X1 port map( A => B(1), ZN => n77);
   U146 : INV_X1 port map( A => net37710, ZN => net26755);
   U147 : INV_X1 port map( A => B(24), ZN => n83);
   U148 : INV_X1 port map( A => B(30), ZN => n75);
   U149 : XNOR2_X1 port map( A => n56, B => B(24), ZN => DIFF_24_port);
   U150 : XOR2_X1 port map( A => n22, B => n91, Z => DIFF_12_port);
   U151 : XOR2_X1 port map( A => n53, B => net37722, Z => DIFF_4_port);
   U152 : XOR2_X1 port map( A => net37633, B => n54, Z => DIFF_13_port);
   U153 : XOR2_X1 port map( A => n37, B => n46, Z => DIFF_25_port);
   U154 : XOR2_X1 port map( A => net37353, B => n16, Z => DIFF_17_port);
   U155 : INV_X1 port map( A => B(23), ZN => n87);
   U156 : INV_X1 port map( A => B(27), ZN => n82);
   U157 : XNOR2_X1 port map( A => n38, B => n69, ZN => DIFF_3_port);
   U158 : XNOR2_X1 port map( A => net37871, B => n68, ZN => DIFF_7_port);
   U159 : INV_X1 port map( A => B(0), ZN => n67);
   U160 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n37, ZN => n80);
   U161 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n45, ZN => n85);
   U162 : INV_X1 port map( A => net37702, ZN => net26789);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor_DW01_add_3 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end branch_predictor_DW01_add_3;

architecture SYN_rpl of branch_predictor_DW01_add_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1036 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1036, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor_DW01_add_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end branch_predictor_DW01_add_2;

architecture SYN_rpl of branch_predictor_DW01_add_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n_1039 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1039, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end branch_predictor_DW01_add_1;

architecture SYN_rpl of branch_predictor_DW01_add_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, SUM_6_port, 
      SUM_7_port, SUM_8_port, SUM_9_port, SUM_10_port, SUM_11_port, SUM_12_port
      , SUM_13_port, SUM_15_port, SUM_16_port, SUM_17_port, SUM_18_port, 
      SUM_19_port, SUM_20_port, SUM_21_port, SUM_22_port, SUM_23_port, 
      SUM_24_port, SUM_25_port, SUM_26_port, SUM_14_port, SUM_27_port, 
      SUM_28_port, SUM_29_port, SUM_30_port, SUM_31_port, SUM_3_port, 
      SUM_4_port, SUM_5_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : AND2_X1 port map( A1 => A(6), A2 => n2, ZN => n1);
   U2 : AND2_X1 port map( A1 => A(5), A2 => n3, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A(30), A2 => n27, ZN => n57);
   U4 : AND2_X1 port map( A1 => A(4), A2 => n4, ZN => n3);
   U5 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n4);
   U6 : AND2_X1 port map( A1 => A(7), A2 => n1, ZN => n5);
   U7 : AND2_X1 port map( A1 => A(8), A2 => n5, ZN => n6);
   U8 : AND2_X1 port map( A1 => A(9), A2 => n6, ZN => n7);
   U9 : AND2_X1 port map( A1 => A(10), A2 => n7, ZN => n8);
   U10 : AND2_X1 port map( A1 => A(11), A2 => n8, ZN => n9);
   U11 : AND2_X1 port map( A1 => A(12), A2 => n9, ZN => n10);
   U12 : AND2_X1 port map( A1 => A(13), A2 => n10, ZN => n11);
   U13 : AND2_X1 port map( A1 => A(14), A2 => n11, ZN => n12);
   U14 : AND2_X1 port map( A1 => A(15), A2 => n12, ZN => n13);
   U15 : AND2_X1 port map( A1 => A(16), A2 => n13, ZN => n14);
   U16 : AND2_X1 port map( A1 => A(17), A2 => n14, ZN => n15);
   U17 : AND2_X1 port map( A1 => A(18), A2 => n15, ZN => n16);
   U18 : AND2_X1 port map( A1 => A(19), A2 => n16, ZN => n17);
   U19 : AND2_X1 port map( A1 => A(20), A2 => n17, ZN => n18);
   U20 : AND2_X1 port map( A1 => A(21), A2 => n18, ZN => n19);
   U21 : AND2_X1 port map( A1 => A(22), A2 => n19, ZN => n20);
   U22 : AND2_X1 port map( A1 => A(23), A2 => n20, ZN => n21);
   U23 : AND2_X1 port map( A1 => A(24), A2 => n21, ZN => n22);
   U24 : AND2_X1 port map( A1 => A(25), A2 => n22, ZN => n23);
   U25 : AND2_X1 port map( A1 => A(26), A2 => n23, ZN => n24);
   U26 : AND2_X1 port map( A1 => A(27), A2 => n24, ZN => n25);
   U27 : AND2_X1 port map( A1 => A(28), A2 => n25, ZN => n26);
   U28 : AND2_X1 port map( A1 => A(29), A2 => n26, ZN => n27);
   U29 : XOR2_X1 port map( A => A(6), B => n2, Z => SUM_6_port);
   U30 : XOR2_X1 port map( A => A(7), B => n1, Z => SUM_7_port);
   U31 : XOR2_X1 port map( A => A(8), B => n5, Z => SUM_8_port);
   U32 : XOR2_X1 port map( A => A(9), B => n6, Z => SUM_9_port);
   U33 : XOR2_X1 port map( A => A(10), B => n7, Z => SUM_10_port);
   U34 : XOR2_X1 port map( A => A(11), B => n8, Z => SUM_11_port);
   U35 : XOR2_X1 port map( A => A(12), B => n9, Z => SUM_12_port);
   U36 : XOR2_X1 port map( A => A(13), B => n10, Z => SUM_13_port);
   U37 : XOR2_X1 port map( A => A(15), B => n12, Z => SUM_15_port);
   U38 : XOR2_X1 port map( A => A(16), B => n13, Z => SUM_16_port);
   U39 : XOR2_X1 port map( A => A(17), B => n14, Z => SUM_17_port);
   U40 : XOR2_X1 port map( A => A(18), B => n15, Z => SUM_18_port);
   U41 : XOR2_X1 port map( A => A(19), B => n16, Z => SUM_19_port);
   U42 : XOR2_X1 port map( A => A(20), B => n17, Z => SUM_20_port);
   U43 : XOR2_X1 port map( A => A(21), B => n18, Z => SUM_21_port);
   U44 : XOR2_X1 port map( A => A(22), B => n19, Z => SUM_22_port);
   U45 : XOR2_X1 port map( A => A(23), B => n20, Z => SUM_23_port);
   U46 : XOR2_X1 port map( A => A(24), B => n21, Z => SUM_24_port);
   U47 : XOR2_X1 port map( A => A(25), B => n22, Z => SUM_25_port);
   U48 : XOR2_X1 port map( A => A(26), B => n23, Z => SUM_26_port);
   U49 : XOR2_X1 port map( A => A(14), B => n11, Z => SUM_14_port);
   U50 : XOR2_X1 port map( A => A(27), B => n24, Z => SUM_27_port);
   U51 : XOR2_X1 port map( A => A(28), B => n25, Z => SUM_28_port);
   U52 : XOR2_X1 port map( A => A(29), B => n26, Z => SUM_29_port);
   U53 : XOR2_X1 port map( A => A(30), B => n27, Z => SUM_30_port);
   U54 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U55 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U56 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U57 : XOR2_X1 port map( A => A(4), B => n4, Z => SUM_4_port);
   U58 : XOR2_X1 port map( A => A(5), B => n3, Z => SUM_5_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end branch_predictor_DW01_add_0;

architecture SYN_rpl of branch_predictor_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n2, n_1076 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1076, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity NPC_adder_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end NPC_adder_DW01_add_0;

architecture SYN_rpl of NPC_adder_DW01_add_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, SUM_3_port, 
      SUM_7_port, SUM_6_port, SUM_5_port, SUM_4_port, SUM_10_port, SUM_11_port,
      SUM_12_port, SUM_13_port, SUM_14_port, SUM_15_port, SUM_16_port, 
      SUM_17_port, SUM_18_port, SUM_19_port, SUM_20_port, SUM_21_port, 
      SUM_22_port, SUM_23_port, SUM_24_port, SUM_25_port, SUM_26_port, 
      SUM_27_port, SUM_28_port, SUM_29_port, SUM_30_port, SUM_8_port, 
      SUM_9_port, SUM_31_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : AND2_X1 port map( A1 => A(6), A2 => n2, ZN => n1);
   U2 : AND2_X1 port map( A1 => A(5), A2 => n3, ZN => n2);
   U3 : AND2_X1 port map( A1 => A(4), A2 => n25, ZN => n3);
   U4 : AND2_X1 port map( A1 => A(9), A2 => n27, ZN => n4);
   U5 : AND2_X1 port map( A1 => A(11), A2 => n15, ZN => n5);
   U6 : AND2_X1 port map( A1 => A(14), A2 => n12, ZN => n6);
   U7 : AND2_X1 port map( A1 => A(17), A2 => n13, ZN => n7);
   U8 : AND2_X1 port map( A1 => A(22), A2 => n11, ZN => n8);
   U9 : AND2_X1 port map( A1 => A(25), A2 => n17, ZN => n9);
   U10 : AND2_X1 port map( A1 => A(28), A2 => n18, ZN => n10);
   U11 : AND2_X1 port map( A1 => A(21), A2 => n16, ZN => n11);
   U12 : AND2_X1 port map( A1 => A(13), A2 => n19, ZN => n12);
   U13 : AND2_X1 port map( A1 => A(16), A2 => n20, ZN => n13);
   U14 : AND2_X1 port map( A1 => A(19), A2 => n21, ZN => n14);
   U15 : AND2_X1 port map( A1 => A(10), A2 => n4, ZN => n15);
   U16 : AND2_X1 port map( A1 => A(20), A2 => n14, ZN => n16);
   U17 : AND2_X1 port map( A1 => A(24), A2 => n22, ZN => n17);
   U18 : AND2_X1 port map( A1 => A(27), A2 => n23, ZN => n18);
   U19 : AND2_X1 port map( A1 => A(12), A2 => n5, ZN => n19);
   U20 : AND2_X1 port map( A1 => A(15), A2 => n6, ZN => n20);
   U21 : AND2_X1 port map( A1 => A(18), A2 => n7, ZN => n21);
   U22 : AND2_X1 port map( A1 => A(23), A2 => n8, ZN => n22);
   U23 : AND2_X1 port map( A1 => A(26), A2 => n9, ZN => n23);
   U24 : AND2_X1 port map( A1 => A(29), A2 => n10, ZN => n24);
   U25 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n25);
   U26 : AND2_X1 port map( A1 => A(7), A2 => n1, ZN => n26);
   U27 : AND2_X1 port map( A1 => A(8), A2 => n26, ZN => n27);
   U28 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U29 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U30 : XOR2_X1 port map( A => A(7), B => n1, Z => SUM_7_port);
   U31 : XOR2_X1 port map( A => A(6), B => n2, Z => SUM_6_port);
   U32 : XOR2_X1 port map( A => A(5), B => n3, Z => SUM_5_port);
   U33 : XOR2_X1 port map( A => A(4), B => n25, Z => SUM_4_port);
   U34 : XOR2_X1 port map( A => A(10), B => n4, Z => SUM_10_port);
   U35 : XOR2_X1 port map( A => A(11), B => n15, Z => SUM_11_port);
   U36 : XOR2_X1 port map( A => A(12), B => n5, Z => SUM_12_port);
   U37 : XOR2_X1 port map( A => A(13), B => n19, Z => SUM_13_port);
   U38 : XOR2_X1 port map( A => A(14), B => n12, Z => SUM_14_port);
   U39 : XOR2_X1 port map( A => A(15), B => n6, Z => SUM_15_port);
   U40 : XOR2_X1 port map( A => A(16), B => n20, Z => SUM_16_port);
   U41 : XOR2_X1 port map( A => A(17), B => n13, Z => SUM_17_port);
   U42 : XOR2_X1 port map( A => A(18), B => n7, Z => SUM_18_port);
   U43 : XOR2_X1 port map( A => A(19), B => n21, Z => SUM_19_port);
   U44 : XOR2_X1 port map( A => A(20), B => n14, Z => SUM_20_port);
   U45 : XOR2_X1 port map( A => A(21), B => n16, Z => SUM_21_port);
   U46 : XOR2_X1 port map( A => A(22), B => n11, Z => SUM_22_port);
   U47 : XOR2_X1 port map( A => A(23), B => n8, Z => SUM_23_port);
   U48 : XOR2_X1 port map( A => A(24), B => n22, Z => SUM_24_port);
   U49 : XOR2_X1 port map( A => A(25), B => n17, Z => SUM_25_port);
   U50 : XOR2_X1 port map( A => A(26), B => n9, Z => SUM_26_port);
   U51 : XOR2_X1 port map( A => A(27), B => n23, Z => SUM_27_port);
   U52 : XOR2_X1 port map( A => A(28), B => n18, Z => SUM_28_port);
   U53 : XOR2_X1 port map( A => A(29), B => n10, Z => SUM_29_port);
   U54 : XOR2_X1 port map( A => A(30), B => n24, Z => SUM_30_port);
   U55 : XOR2_X1 port map( A => A(8), B => n26, Z => SUM_8_port);
   U56 : XOR2_X1 port map( A => A(9), B => n27, Z => SUM_9_port);
   U57 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U58 : NAND2_X1 port map( A1 => A(30), A2 => n24, ZN => n57);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SHIFTER_GENERIC_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW01_ash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW01_ash_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => SH(4), Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => SH(4), Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => SH(4), Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => SH(4), Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => SH(4), Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => SH(4), Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => SH(4), Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => SH(4), Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n23, S => SH(4), Z 
                           => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n19, S => SH(4), Z 
                           => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n21, S => SH(4), Z 
                           => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n17, S => SH(4), Z 
                           => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n22, S => SH(4), Z 
                           => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n18, S => SH(4), Z 
                           => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n20, S => SH(4), Z 
                           => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n16, S => SH(4), Z 
                           => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n13, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n13, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n13, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n13, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n13, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n13, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n13, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n13, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n13, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n13, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n13, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n13, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n12, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n12, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n12, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n12, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n12, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n12, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n12, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n12, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n12, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n12, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n12, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n12, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n10, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n10, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n10, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n10, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n10, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n10, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n10, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n10, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n10, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n10, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n10, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n10, Z => ML_int_3_20_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n10, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n10, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n10, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n9, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n9, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n9, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n9, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n9, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n9, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n9, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n9, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n9, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n9, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n9, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n9, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n7, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n7, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n7, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n7, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n7, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n7, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n6, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n6, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n6, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n6, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n6, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n6, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n6, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n6, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n6, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n6, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n6, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n6, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n5, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n5, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n5, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n5, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n5, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n5, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n5, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n5, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n5, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n5, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n5, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n5, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n3, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n3, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n2, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n2, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n2, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n3, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n1, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n2, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n3, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n3, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n1, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n2, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n1, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n2, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n1, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n3, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n1, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n2, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n1, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n3, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n1, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n2, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n1, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n2, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n1, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n3, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n1, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n2, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n2, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n2, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n2, Z => 
                           ML_int_1_1_port);
   U3 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_19_port, S => 
                           n11, Z => ML_int_3_19_port);
   U4 : INV_X2 port map( A => n11, ZN => n10);
   U5 : INV_X1 port map( A => n11, ZN => n9);
   U6 : INV_X1 port map( A => n30, ZN => n20);
   U7 : INV_X1 port map( A => n31, ZN => n16);
   U8 : INV_X1 port map( A => n29, ZN => n18);
   U9 : INV_X1 port map( A => n28, ZN => n22);
   U10 : INV_X1 port map( A => n26, ZN => n21);
   U11 : INV_X1 port map( A => n27, ZN => n17);
   U12 : INV_X1 port map( A => n25, ZN => n19);
   U13 : INV_X1 port map( A => n24, ZN => n23);
   U14 : INV_X1 port map( A => SH(3), ZN => n14);
   U15 : INV_X1 port map( A => SH(1), ZN => n8);
   U16 : INV_X1 port map( A => SH(0), ZN => n4);
   U17 : INV_X2 port map( A => n4, ZN => n1);
   U18 : INV_X2 port map( A => n4, ZN => n2);
   U19 : INV_X2 port map( A => n8, ZN => n5);
   U20 : INV_X2 port map( A => n8, ZN => n6);
   U21 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => n8, ZN => n7);
   U23 : INV_X1 port map( A => SH(2), ZN => n11);
   U24 : INV_X1 port map( A => n14, ZN => n12);
   U25 : INV_X1 port map( A => n14, ZN => n13);
   U26 : INV_X1 port map( A => SH(4), ZN => n15);
   U27 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n15, ZN => B(9));
   U28 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n15, ZN => B(8));
   U29 : NOR2_X1 port map( A1 => SH(4), A2 => n24, ZN => B(7));
   U30 : NOR2_X1 port map( A1 => SH(4), A2 => n25, ZN => B(6));
   U31 : NOR2_X1 port map( A1 => SH(4), A2 => n26, ZN => B(5));
   U32 : NOR2_X1 port map( A1 => SH(4), A2 => n27, ZN => B(4));
   U33 : NOR2_X1 port map( A1 => SH(4), A2 => n28, ZN => B(3));
   U34 : NOR2_X1 port map( A1 => SH(4), A2 => n29, ZN => B(2));
   U35 : NOR2_X1 port map( A1 => SH(4), A2 => n30, ZN => B(1));
   U36 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n15, ZN => B(15));
   U37 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n15, ZN => B(14));
   U38 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n15, ZN => B(13));
   U39 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n15, ZN => B(12));
   U40 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n15, ZN => B(11));
   U41 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n15, ZN => B(10));
   U42 : NOR2_X1 port map( A1 => SH(4), A2 => n31, ZN => B(0));
   U43 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n14, ZN => n24);
   U44 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n14, ZN => n25);
   U45 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n14, ZN => n26);
   U46 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n14, ZN => n27);
   U47 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n14, ZN => n28);
   U48 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n14, ZN => n29);
   U49 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n14, ZN => n30);
   U50 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n14, ZN => n31);
   U51 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n11, ZN => 
                           ML_int_3_3_port);
   U52 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n11, ZN => 
                           ML_int_3_2_port);
   U53 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n11, ZN => 
                           ML_int_3_1_port);
   U54 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n11, ZN => 
                           ML_int_3_0_port);
   U55 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n8, ZN => 
                           ML_int_2_1_port);
   U56 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n8, ZN => 
                           ML_int_2_0_port);
   U57 : AND2_X1 port map( A1 => A(0), A2 => n4, ZN => ML_int_1_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SHIFTER_GENERIC_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW_rash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rash_0 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165 : std_logic;

begin
   
   U3 : CLKBUF_X1 port map( A => SH(4), Z => n5);
   U4 : AOI221_X1 port map( B1 => n54, B2 => A(7), C1 => n52, C2 => A(6), A => 
                           n165, ZN => n86);
   U5 : AOI221_X1 port map( B1 => n54, B2 => A(11), C1 => n52, C2 => A(10), A 
                           => n156, ZN => n67);
   U6 : AOI221_X1 port map( B1 => n54, B2 => A(13), C1 => n52, C2 => A(12), A 
                           => n153, ZN => n105);
   U7 : INV_X1 port map( A => n140, ZN => n57);
   U8 : AOI221_X1 port map( B1 => n54, B2 => A(10), C1 => n52, C2 => A(9), A =>
                           n99, ZN => n73);
   U9 : NAND2_X2 port map( A1 => SH(1), A2 => SH(0), ZN => n94);
   U10 : INV_X1 port map( A => n97, ZN => n53);
   U11 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n98);
   U12 : AOI221_X1 port map( B1 => n54, B2 => A(12), C1 => n52, C2 => A(11), A 
                           => n122, ZN => n58);
   U13 : NOR2_X2 port map( A1 => n2, A2 => SH(1), ZN => n97);
   U14 : INV_X1 port map( A => n59, ZN => n56);
   U15 : INV_X1 port map( A => SH(4), ZN => n6);
   U16 : INV_X1 port map( A => n89, ZN => n55);
   U17 : INV_X1 port map( A => n160, ZN => n32);
   U18 : INV_X1 port map( A => n126, ZN => n35);
   U19 : INV_X1 port map( A => n139, ZN => n27);
   U20 : INV_X1 port map( A => n94, ZN => n54);
   U21 : INV_X1 port map( A => n128, ZN => n33);
   U22 : INV_X1 port map( A => n95, ZN => n52);
   U23 : INV_X1 port map( A => n81, ZN => n16);
   U24 : INV_X1 port map( A => n138, ZN => B(12));
   U25 : AND2_X2 port map( A1 => n157, A2 => n3, ZN => n63);
   U26 : INV_X1 port map( A => n58, ZN => n8);
   U27 : INV_X1 port map( A => n105, ZN => n7);
   U28 : INV_X1 port map( A => n67, ZN => n10);
   U29 : INV_X1 port map( A => n93, ZN => n11);
   U30 : INV_X1 port map( A => n76, ZN => n18);
   U31 : INV_X1 port map( A => n62, ZN => n15);
   U32 : INV_X1 port map( A => n64, ZN => n21);
   U33 : INV_X1 port map( A => n82, ZN => n23);
   U34 : INV_X1 port map( A => n77, ZN => n25);
   U35 : INV_X1 port map( A => A(3), ZN => n44);
   U36 : INV_X1 port map( A => n125, ZN => n37);
   U37 : INV_X1 port map( A => A(14), ZN => n17);
   U38 : INV_X1 port map( A => A(23), ZN => n30);
   U39 : INV_X1 port map( A => A(12), ZN => n13);
   U40 : INV_X1 port map( A => A(6), ZN => n47);
   U41 : INV_X1 port map( A => A(7), ZN => n48);
   U42 : INV_X1 port map( A => A(31), ZN => n43);
   U43 : INV_X1 port map( A => A(17), ZN => n22);
   U44 : INV_X1 port map( A => A(21), ZN => n29);
   U45 : INV_X1 port map( A => A(20), ZN => n28);
   U46 : INV_X1 port map( A => A(15), ZN => n19);
   U47 : INV_X1 port map( A => A(16), ZN => n20);
   U48 : INV_X1 port map( A => A(29), ZN => n40);
   U49 : INV_X1 port map( A => A(27), ZN => n38);
   U50 : INV_X1 port map( A => A(26), ZN => n36);
   U51 : INV_X1 port map( A => A(30), ZN => n42);
   U52 : INV_X1 port map( A => A(28), ZN => n39);
   U53 : INV_X1 port map( A => A(18), ZN => n24);
   U54 : INV_X1 port map( A => A(19), ZN => n26);
   U55 : INV_X1 port map( A => A(9), ZN => n50);
   U56 : INV_X1 port map( A => A(8), ZN => n49);
   U57 : INV_X1 port map( A => A(10), ZN => n9);
   U58 : INV_X1 port map( A => A(11), ZN => n12);
   U59 : INV_X1 port map( A => A(24), ZN => n31);
   U60 : INV_X1 port map( A => A(25), ZN => n34);
   U61 : AND2_X1 port map( A1 => SH(2), A2 => n157, ZN => n65);
   U62 : INV_X1 port map( A => A(2), ZN => n41);
   U63 : NAND2_X1 port map( A1 => SH(1), A2 => n2, ZN => n95);
   U64 : INV_X1 port map( A => A(5), ZN => n46);
   U65 : INV_X1 port map( A => A(4), ZN => n45);
   U66 : NAND2_X1 port map( A1 => SH(1), A2 => n2, ZN => n1);
   U67 : INV_X1 port map( A => SH(0), ZN => n2);
   U68 : INV_X1 port map( A => SH(2), ZN => n3);
   U69 : INV_X1 port map( A => SH(3), ZN => n4);
   U70 : INV_X2 port map( A => n98, ZN => n51);
   U71 : OAI221_X1 port map( B1 => n58, B2 => n59, C1 => n60, C2 => n6, A => 
                           n61, ZN => B(9));
   U72 : AOI222_X1 port map( A1 => n55, A2 => n62, B1 => n63, B2 => n64, C1 => 
                           n65, C2 => n66, ZN => n61);
   U73 : OAI221_X1 port map( B1 => n67, B2 => n59, C1 => n68, C2 => n6, A => 
                           n69, ZN => B(8));
   U74 : AOI222_X1 port map( A1 => n55, A2 => n70, B1 => n63, B2 => n71, C1 => 
                           n65, C2 => n72, ZN => n69);
   U75 : OAI221_X1 port map( B1 => n73, B2 => n59, C1 => n74, C2 => n6, A => 
                           n75, ZN => B(7));
   U76 : AOI222_X1 port map( A1 => n55, A2 => n11, B1 => n63, B2 => n76, C1 => 
                           n65, C2 => n77, ZN => n75);
   U77 : OAI221_X1 port map( B1 => n78, B2 => n59, C1 => n79, C2 => n6, A => 
                           n80, ZN => B(6));
   U78 : AOI222_X1 port map( A1 => n55, A2 => n7, B1 => n63, B2 => n81, C1 => 
                           n65, C2 => n82, ZN => n80);
   U79 : OAI221_X1 port map( B1 => n83, B2 => n59, C1 => n84, C2 => n6, A => 
                           n85, ZN => B(5));
   U80 : AOI222_X1 port map( A1 => n55, A2 => n8, B1 => n63, B2 => n62, C1 => 
                           n65, C2 => n64, ZN => n85);
   U81 : OAI221_X1 port map( B1 => n86, B2 => n59, C1 => n87, C2 => n6, A => 
                           n88, ZN => B(4));
   U82 : AOI222_X1 port map( A1 => n55, A2 => n10, B1 => n63, B2 => n70, C1 => 
                           n65, C2 => n71, ZN => n88);
   U83 : OAI221_X1 port map( B1 => n73, B2 => n89, C1 => n90, C2 => n6, A => 
                           n91, ZN => B(3));
   U84 : AOI222_X1 port map( A1 => n65, A2 => n76, B1 => n56, B2 => n92, C1 => 
                           n63, C2 => n11, ZN => n91);
   U85 : OAI221_X1 port map( B1 => n94, B2 => n47, C1 => n95, C2 => n46, A => 
                           n96, ZN => n92);
   U86 : AOI22_X1 port map( A1 => A(4), A2 => n97, B1 => A(3), B2 => n98, ZN =>
                           n96);
   U87 : OAI22_X1 port map( A1 => n49, A2 => n53, B1 => n48, B2 => n51, ZN => 
                           n99);
   U88 : AND2_X1 port map( A1 => n56, A2 => n100, ZN => B(31));
   U89 : AND2_X1 port map( A1 => n101, A2 => n56, ZN => B(30));
   U90 : OAI221_X1 port map( B1 => n78, B2 => n89, C1 => n102, C2 => n6, A => 
                           n103, ZN => B(2));
   U91 : AOI222_X1 port map( A1 => n65, A2 => n81, B1 => n56, B2 => n104, C1 =>
                           n63, C2 => n7, ZN => n103);
   U92 : OAI221_X1 port map( B1 => n94, B2 => n46, C1 => n1, C2 => n45, A => 
                           n106, ZN => n104);
   U93 : AOI22_X1 port map( A1 => A(3), A2 => n97, B1 => A(2), B2 => n98, ZN =>
                           n106);
   U94 : AOI221_X1 port map( B1 => n54, B2 => A(9), C1 => n52, C2 => A(8), A =>
                           n107, ZN => n78);
   U95 : OAI22_X1 port map( A1 => n48, A2 => n53, B1 => n47, B2 => n51, ZN => 
                           n107);
   U96 : AND2_X1 port map( A1 => n108, A2 => n56, ZN => B(29));
   U97 : AND2_X1 port map( A1 => n109, A2 => n56, ZN => B(28));
   U98 : NOR3_X1 port map( A1 => n37, A2 => n5, A3 => SH(3), ZN => B(27));
   U99 : NOR2_X1 port map( A1 => n5, A2 => n110, ZN => B(26));
   U100 : NOR2_X1 port map( A1 => n5, A2 => n60, ZN => B(25));
   U101 : AOI22_X1 port map( A1 => n111, A2 => n57, B1 => n108, B2 => n112, ZN 
                           => n60);
   U102 : NOR2_X1 port map( A1 => n5, A2 => n68, ZN => B(24));
   U103 : AOI22_X1 port map( A1 => n113, A2 => n57, B1 => n109, B2 => n112, ZN 
                           => n68);
   U104 : NOR2_X1 port map( A1 => n5, A2 => n74, ZN => B(23));
   U105 : AOI222_X1 port map( A1 => n114, A2 => n112, B1 => n100, B2 => n115, 
                           C1 => n116, C2 => n57, ZN => n74);
   U106 : NOR2_X1 port map( A1 => n5, A2 => n79, ZN => B(22));
   U107 : AOI222_X1 port map( A1 => n117, A2 => n112, B1 => n101, B2 => n115, 
                           C1 => n118, C2 => n57, ZN => n79);
   U108 : NOR2_X1 port map( A1 => n5, A2 => n84, ZN => B(21));
   U109 : AOI222_X1 port map( A1 => n111, A2 => n112, B1 => n108, B2 => n115, 
                           C1 => n66, C2 => n57, ZN => n84);
   U110 : NOR2_X1 port map( A1 => n5, A2 => n87, ZN => B(20));
   U111 : AOI222_X1 port map( A1 => n113, A2 => n112, B1 => n109, B2 => n115, 
                           C1 => n72, C2 => n57, ZN => n87);
   U112 : OAI221_X1 port map( B1 => n83, B2 => n89, C1 => n119, C2 => n6, A => 
                           n120, ZN => B(1));
   U113 : AOI222_X1 port map( A1 => n65, A2 => n62, B1 => n56, B2 => n121, C1 
                           => n63, C2 => n8, ZN => n120);
   U114 : OAI22_X1 port map( A1 => n9, A2 => n53, B1 => n50, B2 => n51, ZN => 
                           n122);
   U115 : OAI221_X1 port map( B1 => n94, B2 => n45, C1 => n1, C2 => n44, A => 
                           n123, ZN => n121);
   U116 : AOI22_X1 port map( A1 => A(2), A2 => n97, B1 => A(1), B2 => n98, ZN 
                           => n123);
   U117 : AOI221_X1 port map( B1 => n54, B2 => A(8), C1 => n52, C2 => A(7), A 
                           => n124, ZN => n83);
   U118 : OAI22_X1 port map( A1 => n47, A2 => n53, B1 => n46, B2 => n51, ZN => 
                           n124);
   U119 : NOR2_X1 port map( A1 => n5, A2 => n90, ZN => B(19));
   U120 : AOI222_X1 port map( A1 => n77, A2 => n57, B1 => n116, B2 => n112, C1 
                           => n125, C2 => SH(3), ZN => n90);
   U121 : NOR2_X1 port map( A1 => n5, A2 => n102, ZN => B(18));
   U122 : AOI221_X1 port map( B1 => n118, B2 => n112, C1 => n82, C2 => n57, A 
                           => n35, ZN => n102);
   U123 : AOI22_X1 port map( A1 => n127, A2 => n101, B1 => n115, B2 => n117, ZN
                           => n126);
   U124 : NOR2_X1 port map( A1 => n5, A2 => n119, ZN => B(17));
   U125 : AOI221_X1 port map( B1 => n66, B2 => n112, C1 => n64, C2 => n57, A =>
                           n33, ZN => n119);
   U126 : AOI22_X1 port map( A1 => n127, A2 => n108, B1 => n115, B2 => n111, ZN
                           => n128);
   U127 : NOR2_X1 port map( A1 => n5, A2 => n129, ZN => B(16));
   U128 : OAI221_X1 port map( B1 => n25, B2 => n89, C1 => n18, C2 => n59, A => 
                           n130, ZN => B(15));
   U129 : AOI222_X1 port map( A1 => n65, A2 => n114, B1 => n131, B2 => n100, C1
                           => n63, C2 => n116, ZN => n130);
   U130 : OAI221_X1 port map( B1 => n23, B2 => n89, C1 => n16, C2 => n59, A => 
                           n132, ZN => B(14));
   U131 : AOI222_X1 port map( A1 => n65, A2 => n117, B1 => n131, B2 => n101, C1
                           => n63, C2 => n118, ZN => n132);
   U132 : OAI221_X1 port map( B1 => n21, B2 => n89, C1 => n15, C2 => n59, A => 
                           n133, ZN => B(13));
   U133 : AOI222_X1 port map( A1 => n65, A2 => n111, B1 => n131, B2 => n108, C1
                           => n63, C2 => n66, ZN => n133);
   U134 : OAI221_X1 port map( B1 => n94, B2 => n31, C1 => n95, C2 => n30, A => 
                           n134, ZN => n66);
   U135 : AOI22_X1 port map( A1 => A(22), A2 => n97, B1 => A(21), B2 => n98, ZN
                           => n134);
   U136 : OAI222_X1 port map( A1 => n53, A2 => n42, B1 => n95, B2 => n43, C1 =>
                           n51, C2 => n40, ZN => n108);
   U137 : OAI221_X1 port map( B1 => n94, B2 => n39, C1 => n1, C2 => n38, A => 
                           n135, ZN => n111);
   U138 : AOI22_X1 port map( A1 => A(26), A2 => n97, B1 => A(25), B2 => n98, ZN
                           => n135);
   U139 : OAI221_X1 port map( B1 => n94, B2 => n20, C1 => n95, C2 => n19, A => 
                           n136, ZN => n62);
   U140 : AOI22_X1 port map( A1 => A(14), A2 => n97, B1 => A(13), B2 => n98, ZN
                           => n136);
   U141 : OAI221_X1 port map( B1 => n94, B2 => n28, C1 => n1, C2 => n26, A => 
                           n137, ZN => n64);
   U142 : AOI22_X1 port map( A1 => A(18), A2 => n97, B1 => A(17), B2 => n98, ZN
                           => n137);
   U143 : AOI221_X1 port map( B1 => n71, B2 => n55, C1 => n70, C2 => n56, A => 
                           n27, ZN => n138);
   U144 : AOI222_X1 port map( A1 => n65, A2 => n113, B1 => n131, B2 => n109, C1
                           => n63, C2 => n72, ZN => n139);
   U145 : NOR2_X1 port map( A1 => n6, A2 => n140, ZN => n131);
   U146 : OAI221_X1 port map( B1 => n18, B2 => n89, C1 => n93, C2 => n59, A => 
                           n141, ZN => B(11));
   U147 : AOI221_X1 port map( B1 => n65, B2 => n116, C1 => n63, C2 => n77, A =>
                           n142, ZN => n141);
   U148 : NOR3_X1 port map( A1 => n6, A2 => SH(3), A3 => n37, ZN => n142);
   U149 : MUX2_X1 port map( A => n114, B => n100, S => SH(2), Z => n125);
   U150 : NOR2_X1 port map( A1 => n43, A2 => n51, ZN => n100);
   U151 : OAI221_X1 port map( B1 => n94, B2 => n42, C1 => n95, C2 => n40, A => 
                           n143, ZN => n114);
   U152 : AOI22_X1 port map( A1 => A(28), A2 => n97, B1 => A(27), B2 => n98, ZN
                           => n143);
   U153 : OAI221_X1 port map( B1 => n28, B2 => n53, C1 => n26, C2 => n51, A => 
                           n144, ZN => n77);
   U154 : AOI22_X1 port map( A1 => A(22), A2 => n54, B1 => A(21), B2 => n52, ZN
                           => n144);
   U155 : OAI221_X1 port map( B1 => n94, B2 => n36, C1 => n1, C2 => n34, A => 
                           n145, ZN => n116);
   U156 : AOI22_X1 port map( A1 => A(24), A2 => n97, B1 => A(23), B2 => n98, ZN
                           => n145);
   U157 : AOI221_X1 port map( B1 => n54, B2 => A(14), C1 => n52, C2 => A(13), A
                           => n146, ZN => n93);
   U158 : OAI22_X1 port map( A1 => n13, A2 => n53, B1 => n12, B2 => n51, ZN => 
                           n146);
   U159 : OAI221_X1 port map( B1 => n94, B2 => n24, C1 => n95, C2 => n22, A => 
                           n147, ZN => n76);
   U160 : AOI22_X1 port map( A1 => A(16), A2 => n97, B1 => A(15), B2 => n98, ZN
                           => n147);
   U161 : OAI221_X1 port map( B1 => n105, B2 => n59, C1 => n110, C2 => n6, A =>
                           n148, ZN => B(10));
   U162 : AOI222_X1 port map( A1 => n55, A2 => n81, B1 => n63, B2 => n82, C1 =>
                           n65, C2 => n118, ZN => n148);
   U163 : OAI221_X1 port map( B1 => n94, B2 => n34, C1 => n1, C2 => n31, A => 
                           n149, ZN => n118);
   U164 : AOI22_X1 port map( A1 => A(23), A2 => n97, B1 => A(22), B2 => n98, ZN
                           => n149);
   U165 : OAI221_X1 port map( B1 => n94, B2 => n29, C1 => n28, C2 => n1, A => 
                           n150, ZN => n82);
   U166 : AOI22_X1 port map( A1 => n97, A2 => A(19), B1 => n98, B2 => A(18), ZN
                           => n150);
   U167 : OAI221_X1 port map( B1 => n94, B2 => n22, C1 => n95, C2 => n20, A => 
                           n151, ZN => n81);
   U168 : AOI22_X1 port map( A1 => A(15), A2 => n97, B1 => A(14), B2 => n98, ZN
                           => n151);
   U169 : AOI22_X1 port map( A1 => n117, A2 => n57, B1 => n101, B2 => n112, ZN 
                           => n110);
   U170 : OAI22_X1 port map( A1 => n51, A2 => n42, B1 => n53, B2 => n43, ZN => 
                           n101);
   U171 : OAI221_X1 port map( B1 => n94, B2 => n40, C1 => n1, C2 => n39, A => 
                           n152, ZN => n117);
   U172 : AOI22_X1 port map( A1 => A(27), A2 => n97, B1 => A(26), B2 => n98, ZN
                           => n152);
   U173 : OAI22_X1 port map( A1 => n12, A2 => n53, B1 => n9, B2 => n51, ZN => 
                           n153);
   U174 : OAI221_X1 port map( B1 => n86, B2 => n89, C1 => n129, C2 => n6, A => 
                           n154, ZN => B(0));
   U175 : AOI222_X1 port map( A1 => n65, A2 => n70, B1 => n56, B2 => n155, C1 
                           => n63, C2 => n10, ZN => n154);
   U176 : OAI22_X1 port map( A1 => n50, A2 => n53, B1 => n49, B2 => n51, ZN => 
                           n156);
   U177 : OAI221_X1 port map( B1 => n94, B2 => n44, C1 => n95, C2 => n41, A => 
                           n158, ZN => n155);
   U178 : AOI22_X1 port map( A1 => A(1), A2 => n97, B1 => A(0), B2 => n98, ZN 
                           => n158);
   U179 : NAND2_X1 port map( A1 => n57, A2 => n6, ZN => n59);
   U180 : OAI221_X1 port map( B1 => n94, B2 => n19, C1 => n1, C2 => n17, A => 
                           n159, ZN => n70);
   U181 : AOI22_X1 port map( A1 => A(13), A2 => n97, B1 => A(12), B2 => n98, ZN
                           => n159);
   U182 : NOR2_X1 port map( A1 => n4, A2 => SH(4), ZN => n157);
   U183 : AOI221_X1 port map( B1 => n72, B2 => n112, C1 => n71, C2 => n57, A =>
                           n32, ZN => n129);
   U184 : AOI22_X1 port map( A1 => n127, A2 => n109, B1 => n115, B2 => n113, ZN
                           => n160);
   U185 : OAI221_X1 port map( B1 => n94, B2 => n38, C1 => n95, C2 => n36, A => 
                           n161, ZN => n113);
   U186 : AOI22_X1 port map( A1 => A(25), A2 => n97, B1 => A(24), B2 => n98, ZN
                           => n161);
   U187 : NOR2_X1 port map( A1 => n4, A2 => SH(2), ZN => n115);
   U188 : OAI221_X1 port map( B1 => n94, B2 => n43, C1 => n1, C2 => n42, A => 
                           n162, ZN => n109);
   U189 : AOI22_X1 port map( A1 => A(29), A2 => n97, B1 => A(28), B2 => n98, ZN
                           => n162);
   U190 : NOR2_X1 port map( A1 => n3, A2 => n4, ZN => n127);
   U191 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n140);
   U192 : OAI221_X1 port map( B1 => n94, B2 => n26, C1 => n1, C2 => n24, A => 
                           n163, ZN => n71);
   U193 : AOI22_X1 port map( A1 => A(17), A2 => n97, B1 => A(16), B2 => n98, ZN
                           => n163);
   U194 : OAI221_X1 port map( B1 => n53, B2 => n29, C1 => n28, C2 => n51, A => 
                           n164, ZN => n72);
   U195 : AOI22_X1 port map( A1 => A(23), A2 => n54, B1 => A(22), B2 => n52, ZN
                           => n164);
   U196 : NAND2_X1 port map( A1 => n112, A2 => n6, ZN => n89);
   U197 : NOR2_X1 port map( A1 => n3, A2 => SH(3), ZN => n112);
   U198 : OAI22_X1 port map( A1 => n46, A2 => n53, B1 => n45, B2 => n51, ZN => 
                           n165);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SHIFTER_GENERIC_N32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sra_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sra_0 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : INV_X1 port map( A => SH(1), ZN => n6);
   U3 : AOI221_X1 port map( B1 => n95, B2 => A(14), C1 => n96, C2 => A(15), A 
                           => n17, ZN => n150);
   U4 : AOI221_X1 port map( B1 => n95, B2 => A(8), C1 => n96, C2 => A(9), A => 
                           n107, ZN => n79);
   U5 : AOI221_X1 port map( B1 => n95, B2 => A(9), C1 => n96, C2 => A(10), A =>
                           n97, ZN => n74);
   U6 : AOI221_X1 port map( B1 => n95, B2 => A(11), C1 => n96, C2 => A(12), A 
                           => n131, ZN => n61);
   U7 : AOI221_X1 port map( B1 => n112, B2 => n113, C1 => n114, C2 => n115, A 
                           => n46, ZN => n63);
   U8 : NOR2_X2 port map( A1 => n6, A2 => SH(0), ZN => n95);
   U9 : AOI221_X1 port map( B1 => n118, B2 => n113, C1 => n119, C2 => n115, A 
                           => n46, ZN => n75);
   U10 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n115);
   U11 : INV_X1 port map( A => n99, ZN => n1);
   U12 : NAND2_X1 port map( A1 => n60, A2 => n12, ZN => n2);
   U13 : NAND2_X1 port map( A1 => n65, A2 => n16, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n67, A2 => n72, ZN => n4);
   U15 : AND3_X1 port map( A1 => n2, A2 => n3, A3 => n4, ZN => n88);
   U16 : INV_X1 port map( A => n99, ZN => n57);
   U17 : INV_X2 port map( A => n89, ZN => n60);
   U18 : AND2_X2 port map( A1 => SH(2), A2 => n167, ZN => n67);
   U19 : AOI221_X1 port map( B1 => n95, B2 => A(10), C1 => n96, C2 => A(11), A 
                           => n166, ZN => n69);
   U20 : INV_X2 port map( A => n98, ZN => n55);
   U21 : NAND2_X2 port map( A1 => n5, A2 => n6, ZN => n99);
   U22 : INV_X2 port map( A => n95, ZN => n58);
   U23 : NAND2_X2 port map( A1 => n115, A2 => n8, ZN => n62);
   U24 : INV_X1 port map( A => n96, ZN => n56);
   U25 : INV_X1 port map( A => SH(4), ZN => n8);
   U26 : INV_X1 port map( A => n62, ZN => n59);
   U27 : INV_X1 port map( A => n138, ZN => n24);
   U28 : INV_X1 port map( A => n139, ZN => n33);
   U29 : INV_X1 port map( A => n127, ZN => n39);
   U30 : INV_X1 port map( A => n135, ZN => n36);
   U31 : INV_X1 port map( A => n170, ZN => n32);
   U32 : INV_X1 port map( A => n126, ZN => n40);
   U33 : INV_X1 port map( A => n122, ZN => n43);
   U34 : NOR2_X2 port map( A1 => n5, A2 => n6, ZN => n96);
   U35 : INV_X1 port map( A => n101, ZN => n47);
   U36 : INV_X1 port map( A => n78, ZN => n26);
   U37 : AND2_X2 port map( A1 => n167, A2 => n7, ZN => n65);
   U38 : INV_X1 port map( A => n133, ZN => n18);
   U39 : INV_X1 port map( A => n150, ZN => n16);
   U40 : INV_X1 port map( A => n142, ZN => n20);
   U41 : INV_X1 port map( A => n136, ZN => n46);
   U42 : INV_X1 port map( A => n69, ZN => n12);
   U43 : INV_X1 port map( A => n61, ZN => n10);
   U44 : INV_X1 port map( A => n105, ZN => n9);
   U45 : INV_X1 port map( A => n93, ZN => n13);
   U46 : INV_X1 port map( A => n77, ZN => n22);
   U47 : INV_X1 port map( A => A(3), ZN => n48);
   U48 : INV_X1 port map( A => A(17), ZN => n23);
   U49 : INV_X1 port map( A => A(12), ZN => n15);
   U50 : INV_X1 port map( A => n149, ZN => n19);
   U51 : INV_X1 port map( A => n161, ZN => n21);
   U52 : INV_X1 port map( A => A(23), ZN => n30);
   U53 : INV_X1 port map( A => A(21), ZN => n29);
   U54 : INV_X1 port map( A => A(6), ZN => n51);
   U55 : INV_X1 port map( A => A(7), ZN => n52);
   U56 : INV_X1 port map( A => A(31), ZN => n45);
   U57 : INV_X1 port map( A => A(18), ZN => n25);
   U58 : INV_X1 port map( A => A(19), ZN => n27);
   U59 : INV_X1 port map( A => A(29), ZN => n41);
   U60 : INV_X1 port map( A => A(27), ZN => n37);
   U61 : INV_X1 port map( A => A(26), ZN => n35);
   U62 : INV_X1 port map( A => A(28), ZN => n38);
   U63 : INV_X1 port map( A => A(20), ZN => n28);
   U64 : INV_X1 port map( A => A(30), ZN => n44);
   U65 : INV_X1 port map( A => A(9), ZN => n54);
   U66 : INV_X1 port map( A => A(8), ZN => n53);
   U67 : INV_X1 port map( A => A(10), ZN => n11);
   U68 : INV_X1 port map( A => A(11), ZN => n14);
   U69 : INV_X1 port map( A => A(24), ZN => n31);
   U70 : INV_X1 port map( A => A(25), ZN => n34);
   U71 : INV_X1 port map( A => n169, ZN => n17);
   U72 : INV_X1 port map( A => A(2), ZN => n42);
   U73 : NAND2_X1 port map( A1 => SH(0), A2 => n6, ZN => n98);
   U74 : INV_X1 port map( A => A(5), ZN => n50);
   U75 : INV_X1 port map( A => A(4), ZN => n49);
   U76 : INV_X1 port map( A => SH(0), ZN => n5);
   U77 : INV_X1 port map( A => SH(2), ZN => n7);
   U78 : OAI221_X1 port map( B1 => n61, B2 => n62, C1 => n63, C2 => n8, A => 
                           n64, ZN => B_9_port);
   U79 : AOI222_X1 port map( A1 => n60, A2 => n18, B1 => n65, B2 => n66, C1 => 
                           n67, C2 => n68, ZN => n64);
   U80 : OAI221_X1 port map( B1 => n69, B2 => n62, C1 => n70, C2 => n8, A => 
                           n71, ZN => B_8_port);
   U81 : AOI222_X1 port map( A1 => n60, A2 => n16, B1 => n65, B2 => n72, C1 => 
                           n67, C2 => n73, ZN => n71);
   U82 : OAI221_X1 port map( B1 => n74, B2 => n62, C1 => n75, C2 => n8, A => 
                           n76, ZN => B_7_port);
   U83 : AOI222_X1 port map( A1 => n60, A2 => n13, B1 => n65, B2 => n77, C1 => 
                           n67, C2 => n78, ZN => n76);
   U84 : OAI221_X1 port map( B1 => n79, B2 => n62, C1 => n80, C2 => n8, A => 
                           n81, ZN => B_6_port);
   U85 : AOI222_X1 port map( A1 => n60, A2 => n9, B1 => n65, B2 => n20, C1 => 
                           n67, C2 => n82, ZN => n81);
   U86 : OAI221_X1 port map( B1 => n83, B2 => n62, C1 => n84, C2 => n8, A => 
                           n85, ZN => B_5_port);
   U87 : AOI222_X1 port map( A1 => n60, A2 => n10, B1 => n65, B2 => n18, C1 => 
                           n67, C2 => n66, ZN => n85);
   U88 : OAI221_X1 port map( B1 => n86, B2 => n62, C1 => n87, C2 => n8, A => 
                           n88, ZN => B_4_port);
   U89 : OAI221_X1 port map( B1 => n74, B2 => n89, C1 => n90, C2 => n8, A => 
                           n91, ZN => B_3_port);
   U90 : AOI222_X1 port map( A1 => n67, A2 => n77, B1 => n59, B2 => n92, C1 => 
                           n65, C2 => n13, ZN => n91);
   U91 : OAI221_X1 port map( B1 => n58, B2 => n50, C1 => n56, C2 => n51, A => 
                           n94, ZN => n92);
   U92 : AOI22_X1 port map( A1 => A(4), A2 => n55, B1 => A(3), B2 => n1, ZN => 
                           n94);
   U93 : OAI22_X1 port map( A1 => n53, A2 => n98, B1 => n52, B2 => n99, ZN => 
                           n97);
   U94 : OAI21_X1 port map( B1 => SH(4), B2 => n100, A => n101, ZN => B_30_port
                           );
   U95 : OAI221_X1 port map( B1 => n79, B2 => n89, C1 => n102, C2 => n8, A => 
                           n103, ZN => B_2_port);
   U96 : AOI222_X1 port map( A1 => n67, A2 => n20, B1 => n59, B2 => n104, C1 =>
                           n65, C2 => n9, ZN => n103);
   U97 : OAI221_X1 port map( B1 => n58, B2 => n49, C1 => n56, C2 => n50, A => 
                           n106, ZN => n104);
   U98 : AOI22_X1 port map( A1 => A(3), A2 => n55, B1 => A(2), B2 => n1, ZN => 
                           n106);
   U99 : OAI22_X1 port map( A1 => n52, A2 => n98, B1 => n51, B2 => n99, ZN => 
                           n107);
   U100 : OAI21_X1 port map( B1 => SH(4), B2 => n108, A => n101, ZN => 
                           B_29_port);
   U101 : OAI21_X1 port map( B1 => SH(4), B2 => n109, A => n101, ZN => 
                           B_28_port);
   U102 : OAI21_X1 port map( B1 => SH(4), B2 => n110, A => n101, ZN => 
                           B_27_port);
   U103 : OAI21_X1 port map( B1 => SH(4), B2 => n111, A => n101, ZN => 
                           B_26_port);
   U104 : OAI21_X1 port map( B1 => SH(4), B2 => n63, A => n101, ZN => B_25_port
                           );
   U105 : OAI21_X1 port map( B1 => SH(4), B2 => n70, A => n101, ZN => B_24_port
                           );
   U106 : AOI221_X1 port map( B1 => n116, B2 => n113, C1 => n117, C2 => n115, A
                           => n46, ZN => n70);
   U107 : OAI21_X1 port map( B1 => SH(4), B2 => n75, A => n101, ZN => B_23_port
                           );
   U108 : OAI21_X1 port map( B1 => SH(4), B2 => n80, A => n101, ZN => B_22_port
                           );
   U109 : AOI221_X1 port map( B1 => n120, B2 => n113, C1 => n121, C2 => n115, A
                           => n43, ZN => n80);
   U110 : AOI21_X1 port map( B1 => n123, B2 => n124, A => n125, ZN => n122);
   U111 : OAI21_X1 port map( B1 => SH(4), B2 => n84, A => n101, ZN => B_21_port
                           );
   U112 : AOI221_X1 port map( B1 => n114, B2 => n113, C1 => n68, C2 => n115, A 
                           => n40, ZN => n84);
   U113 : AOI21_X1 port map( B1 => n123, B2 => n112, A => n125, ZN => n126);
   U114 : OAI21_X1 port map( B1 => SH(4), B2 => n87, A => n101, ZN => B_20_port
                           );
   U115 : AOI221_X1 port map( B1 => n117, B2 => n113, C1 => n73, C2 => n115, A 
                           => n39, ZN => n87);
   U116 : AOI21_X1 port map( B1 => n123, B2 => n116, A => n125, ZN => n127);
   U117 : OAI221_X1 port map( B1 => n83, B2 => n89, C1 => n128, C2 => n8, A => 
                           n129, ZN => B_1_port);
   U118 : AOI222_X1 port map( A1 => n67, A2 => n18, B1 => n59, B2 => n130, C1 
                           => n65, C2 => n10, ZN => n129);
   U119 : OAI22_X1 port map( A1 => n11, A2 => n98, B1 => n54, B2 => n99, ZN => 
                           n131);
   U120 : OAI221_X1 port map( B1 => n58, B2 => n48, C1 => n56, C2 => n49, A => 
                           n132, ZN => n130);
   U121 : AOI22_X1 port map( A1 => A(2), A2 => n55, B1 => A(1), B2 => n1, ZN =>
                           n132);
   U122 : AOI221_X1 port map( B1 => n95, B2 => A(7), C1 => n96, C2 => A(8), A 
                           => n134, ZN => n83);
   U123 : OAI22_X1 port map( A1 => n51, A2 => n98, B1 => n50, B2 => n99, ZN => 
                           n134);
   U124 : OAI21_X1 port map( B1 => SH(4), B2 => n90, A => n101, ZN => B_19_port
                           );
   U125 : AOI221_X1 port map( B1 => n119, B2 => n113, C1 => n78, C2 => n115, A 
                           => n36, ZN => n90);
   U126 : AOI21_X1 port map( B1 => n123, B2 => n118, A => n125, ZN => n135);
   U127 : NOR2_X1 port map( A1 => n136, A2 => n7, ZN => n125);
   U128 : OAI21_X1 port map( B1 => SH(4), B2 => n102, A => n101, ZN => 
                           B_18_port);
   U129 : AOI221_X1 port map( B1 => n124, B2 => n137, C1 => n120, C2 => n123, A
                           => n24, ZN => n102);
   U130 : AOI22_X1 port map( A1 => n113, A2 => n121, B1 => n115, B2 => n82, ZN 
                           => n138);
   U131 : OAI21_X1 port map( B1 => SH(4), B2 => n128, A => n101, ZN => 
                           B_17_port);
   U132 : AOI221_X1 port map( B1 => n68, B2 => n113, C1 => n66, C2 => n115, A 
                           => n33, ZN => n128);
   U133 : AOI22_X1 port map( A1 => n137, A2 => n112, B1 => n123, B2 => n114, ZN
                           => n139);
   U134 : OAI21_X1 port map( B1 => SH(4), B2 => n140, A => n101, ZN => 
                           B_16_port);
   U135 : OAI221_X1 port map( B1 => n26, B2 => n89, C1 => n22, C2 => n62, A => 
                           n141, ZN => B_15_port);
   U136 : AOI221_X1 port map( B1 => n67, B2 => n118, C1 => n65, C2 => n119, A 
                           => n47, ZN => n141);
   U137 : NAND2_X1 port map( A1 => SH(4), A2 => A(31), ZN => n101);
   U138 : OAI221_X1 port map( B1 => n142, B2 => n62, C1 => n100, C2 => n8, A =>
                           n143, ZN => B_14_port);
   U139 : AOI222_X1 port map( A1 => n60, A2 => n82, B1 => n65, B2 => n121, C1 
                           => n67, C2 => n120, ZN => n143);
   U140 : AOI21_X1 port map( B1 => n124, B2 => n115, A => n144, ZN => n100);
   U141 : OAI221_X1 port map( B1 => n133, B2 => n62, C1 => n108, C2 => n8, A =>
                           n145, ZN => B_13_port);
   U142 : AOI222_X1 port map( A1 => n60, A2 => n66, B1 => n65, B2 => n68, C1 =>
                           n67, C2 => n114, ZN => n145);
   U143 : OAI221_X1 port map( B1 => n58, B2 => n37, C1 => n56, C2 => n38, A => 
                           n146, ZN => n114);
   U144 : AOI22_X1 port map( A1 => A(26), A2 => n55, B1 => A(25), B2 => n57, ZN
                           => n146);
   U145 : OAI221_X1 port map( B1 => n58, B2 => n30, C1 => n56, C2 => n31, A => 
                           n147, ZN => n68);
   U146 : AOI22_X1 port map( A1 => A(22), A2 => n55, B1 => A(21), B2 => n57, ZN
                           => n147);
   U147 : OAI221_X1 port map( B1 => n58, B2 => n27, C1 => n56, C2 => n28, A => 
                           n148, ZN => n66);
   U148 : AOI22_X1 port map( A1 => A(18), A2 => n55, B1 => A(17), B2 => n57, ZN
                           => n148);
   U149 : AOI21_X1 port map( B1 => n112, B2 => n115, A => n144, ZN => n108);
   U150 : OAI222_X1 port map( A1 => n99, A2 => n41, B1 => n98, B2 => n44, C1 =>
                           n6, C2 => n45, ZN => n112);
   U151 : AOI221_X1 port map( B1 => n95, B2 => A(15), C1 => n96, C2 => A(16), A
                           => n19, ZN => n133);
   U152 : AOI22_X1 port map( A1 => A(14), A2 => n55, B1 => A(13), B2 => n57, ZN
                           => n149);
   U153 : OAI221_X1 port map( B1 => n150, B2 => n62, C1 => n109, C2 => n8, A =>
                           n151, ZN => B_12_port);
   U154 : AOI222_X1 port map( A1 => n60, A2 => n72, B1 => n65, B2 => n73, C1 =>
                           n67, C2 => n117, ZN => n151);
   U155 : AOI21_X1 port map( B1 => n116, B2 => n115, A => n144, ZN => n109);
   U156 : OAI221_X1 port map( B1 => n93, B2 => n62, C1 => n110, C2 => n8, A => 
                           n152, ZN => B_11_port);
   U157 : AOI222_X1 port map( A1 => n60, A2 => n77, B1 => n65, B2 => n78, C1 =>
                           n67, C2 => n119, ZN => n152);
   U158 : OAI221_X1 port map( B1 => n58, B2 => n34, C1 => n56, C2 => n35, A => 
                           n153, ZN => n119);
   U159 : AOI22_X1 port map( A1 => A(24), A2 => n55, B1 => A(23), B2 => n57, ZN
                           => n153);
   U160 : OAI221_X1 port map( B1 => n28, B2 => n98, C1 => n27, C2 => n99, A => 
                           n154, ZN => n78);
   U161 : AOI22_X1 port map( A1 => A(21), A2 => n95, B1 => A(22), B2 => n96, ZN
                           => n154);
   U162 : OAI221_X1 port map( B1 => n58, B2 => n23, C1 => n56, C2 => n25, A => 
                           n155, ZN => n77);
   U163 : AOI22_X1 port map( A1 => A(16), A2 => n55, B1 => A(15), B2 => n1, ZN 
                           => n155);
   U164 : AOI21_X1 port map( B1 => n118, B2 => n115, A => n144, ZN => n110);
   U165 : OAI21_X1 port map( B1 => n7, B2 => n45, A => n136, ZN => n144);
   U166 : OAI221_X1 port map( B1 => n58, B2 => n41, C1 => n56, C2 => n44, A => 
                           n156, ZN => n118);
   U167 : AOI22_X1 port map( A1 => A(28), A2 => n55, B1 => A(27), B2 => n57, ZN
                           => n156);
   U168 : AOI221_X1 port map( B1 => n95, B2 => A(13), C1 => n96, C2 => A(14), A
                           => n157, ZN => n93);
   U169 : OAI22_X1 port map( A1 => n15, A2 => n98, B1 => n14, B2 => n99, ZN => 
                           n157);
   U170 : OAI221_X1 port map( B1 => n105, B2 => n62, C1 => n111, C2 => n8, A =>
                           n158, ZN => B_10_port);
   U171 : AOI222_X1 port map( A1 => n60, A2 => n20, B1 => n65, B2 => n82, C1 =>
                           n67, C2 => n121, ZN => n158);
   U172 : OAI221_X1 port map( B1 => n58, B2 => n31, C1 => n56, C2 => n34, A => 
                           n159, ZN => n121);
   U173 : AOI22_X1 port map( A1 => A(23), A2 => n55, B1 => A(22), B2 => n57, ZN
                           => n159);
   U174 : OAI221_X1 port map( B1 => n27, B2 => n98, C1 => n25, C2 => n99, A => 
                           n160, ZN => n82);
   U175 : AOI22_X1 port map( A1 => A(20), A2 => n95, B1 => A(21), B2 => n96, ZN
                           => n160);
   U176 : AOI221_X1 port map( B1 => n95, B2 => A(16), C1 => n96, C2 => A(17), A
                           => n21, ZN => n142);
   U177 : AOI22_X1 port map( A1 => A(15), A2 => n55, B1 => A(14), B2 => n57, ZN
                           => n161);
   U178 : AOI221_X1 port map( B1 => n124, B2 => n113, C1 => n120, C2 => n115, A
                           => n46, ZN => n111);
   U179 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n136);
   U180 : OAI221_X1 port map( B1 => n58, B2 => n38, C1 => n56, C2 => n41, A => 
                           n162, ZN => n120);
   U181 : AOI22_X1 port map( A1 => A(27), A2 => n55, B1 => A(26), B2 => n57, ZN
                           => n162);
   U182 : MUX2_X1 port map( A => A(30), B => A(31), S => n99, Z => n124);
   U183 : AOI221_X1 port map( B1 => n95, B2 => A(12), C1 => n96, C2 => A(13), A
                           => n163, ZN => n105);
   U184 : OAI22_X1 port map( A1 => n14, A2 => n98, B1 => n11, B2 => n99, ZN => 
                           n163);
   U185 : OAI221_X1 port map( B1 => n86, B2 => n89, C1 => n140, C2 => n8, A => 
                           n164, ZN => B_0_port);
   U186 : AOI222_X1 port map( A1 => n67, A2 => n16, B1 => n59, B2 => n165, C1 
                           => n65, C2 => n12, ZN => n164);
   U187 : OAI22_X1 port map( A1 => n54, A2 => n98, B1 => n53, B2 => n99, ZN => 
                           n166);
   U188 : OAI221_X1 port map( B1 => n58, B2 => n42, C1 => n56, C2 => n48, A => 
                           n168, ZN => n165);
   U189 : AOI22_X1 port map( A1 => A(1), A2 => n55, B1 => A(0), B2 => n1, ZN =>
                           n168);
   U190 : AOI22_X1 port map( A1 => A(13), A2 => n55, B1 => A(12), B2 => n57, ZN
                           => n169);
   U191 : AND2_X1 port map( A1 => SH(3), A2 => n8, ZN => n167);
   U192 : AOI221_X1 port map( B1 => n73, B2 => n113, C1 => n72, C2 => n115, A 
                           => n32, ZN => n140);
   U193 : AOI22_X1 port map( A1 => n137, A2 => n116, B1 => n123, B2 => n117, ZN
                           => n170);
   U194 : OAI221_X1 port map( B1 => n58, B2 => n35, C1 => n56, C2 => n37, A => 
                           n171, ZN => n117);
   U195 : AOI22_X1 port map( A1 => A(25), A2 => n55, B1 => A(24), B2 => n57, ZN
                           => n171);
   U196 : AND2_X1 port map( A1 => SH(3), A2 => n7, ZN => n123);
   U197 : OAI221_X1 port map( B1 => n58, B2 => n44, C1 => n56, C2 => n45, A => 
                           n172, ZN => n116);
   U198 : AOI22_X1 port map( A1 => A(29), A2 => n55, B1 => A(28), B2 => n57, ZN
                           => n172);
   U199 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n137);
   U200 : OAI221_X1 port map( B1 => n58, B2 => n25, C1 => n27, C2 => n56, A => 
                           n173, ZN => n72);
   U201 : AOI22_X1 port map( A1 => A(17), A2 => n55, B1 => A(16), B2 => n57, ZN
                           => n173);
   U202 : OAI221_X1 port map( B1 => n98, B2 => n29, C1 => n28, C2 => n99, A => 
                           n174, ZN => n73);
   U203 : AOI22_X1 port map( A1 => A(22), A2 => n95, B1 => A(23), B2 => n96, ZN
                           => n174);
   U204 : NAND2_X1 port map( A1 => n113, A2 => n8, ZN => n89);
   U205 : NOR2_X1 port map( A1 => n7, A2 => SH(3), ZN => n113);
   U206 : AOI221_X1 port map( B1 => n95, B2 => A(6), C1 => n96, C2 => A(7), A 
                           => n175, ZN => n86);
   U207 : OAI22_X1 port map( A1 => n50, A2 => n98, B1 => n49, B2 => n99, ZN => 
                           n175);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity comparator_N32_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_N32_DW01_cmp6_0;

architecture SYN_rpl of comparator_N32_DW01_cmp6_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A(0), ZN => n2);
   U2 : INV_X1 port map( A => A(1), ZN => n3);
   U3 : INV_X1 port map( A => B(1), ZN => n1);
   U4 : NOR4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => EQ);
   U5 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n7);
   U6 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n11);
   U7 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n10);
   U8 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n9);
   U9 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n8);
   U10 : NAND4_X1 port map( A1 => n12, A2 => n13, A3 => n14, A4 => n15, ZN => 
                           n6);
   U11 : OAI22_X1 port map( A1 => n16, A2 => n3, B1 => B(1), B2 => n16, ZN => 
                           n15);
   U12 : AND2_X1 port map( A1 => B(0), A2 => n2, ZN => n16);
   U13 : OAI22_X1 port map( A1 => A(1), A2 => n17, B1 => n17, B2 => n1, ZN => 
                           n14);
   U14 : NOR2_X1 port map( A1 => n2, A2 => B(0), ZN => n17);
   U15 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n13);
   U16 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n12);
   U17 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n5);
   U18 : NOR4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           n19);
   U19 : XOR2_X1 port map( A => B(10), B => A(10), Z => n23);
   U20 : XOR2_X1 port map( A => B(9), B => A(9), Z => n22);
   U21 : XOR2_X1 port map( A => B(8), B => A(8), Z => n21);
   U22 : XOR2_X1 port map( A => B(7), B => A(7), Z => n20);
   U23 : NOR4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           n18);
   U24 : XOR2_X1 port map( A => B(14), B => A(14), Z => n27);
   U25 : XOR2_X1 port map( A => B(13), B => A(13), Z => n26);
   U26 : XOR2_X1 port map( A => B(12), B => A(12), Z => n25);
   U27 : XOR2_X1 port map( A => B(11), B => A(11), Z => n24);
   U28 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n4);
   U29 : NOR4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => n35, ZN => 
                           n31);
   U30 : XOR2_X1 port map( A => B(18), B => A(18), Z => n35);
   U31 : XOR2_X1 port map( A => B(17), B => A(17), Z => n34);
   U32 : XOR2_X1 port map( A => B(16), B => A(16), Z => n33);
   U33 : XOR2_X1 port map( A => B(15), B => A(15), Z => n32);
   U34 : NOR4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => 
                           n30);
   U35 : XOR2_X1 port map( A => B(22), B => A(22), Z => n39);
   U36 : XOR2_X1 port map( A => B(21), B => A(21), Z => n38);
   U37 : XOR2_X1 port map( A => B(20), B => A(20), Z => n37);
   U38 : XOR2_X1 port map( A => B(19), B => A(19), Z => n36);
   U39 : NOR4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n29);
   U40 : XOR2_X1 port map( A => B(26), B => A(26), Z => n43);
   U41 : XOR2_X1 port map( A => B(25), B => A(25), Z => n42);
   U42 : XOR2_X1 port map( A => B(24), B => A(24), Z => n41);
   U43 : XOR2_X1 port map( A => B(23), B => A(23), Z => n40);
   U44 : NOR4_X1 port map( A1 => n44, A2 => n45, A3 => n46, A4 => n47, ZN => 
                           n28);
   U45 : XOR2_X1 port map( A => B(30), B => A(30), Z => n47);
   U46 : XOR2_X1 port map( A => B(29), B => A(29), Z => n46);
   U47 : XOR2_X1 port map( A => B(28), B => A(28), Z => n45);
   U48 : XOR2_X1 port map( A => B(27), B => A(27), Z => n44);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => n6, Z => n1);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n4, n5, n6, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n1, A2 => n9, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => S);
   U5 : INV_X1 port map( A => Ci, ZN => n1);
   U6 : INV_X1 port map( A => n9, ZN => n4);
   U7 : INV_X1 port map( A => n8, ZN => Co);
   U8 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n9, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => n1);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => n2);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n2, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => B, ZN => n3);
   U8 : OAI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U7 : INV_X1 port map( A => n5, ZN => n6);
   U8 : XOR2_X1 port map( A => n1, B => n6, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => n1, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U3 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n1, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n3, B2 => n2, ZN => Co);
   U7 : INV_X1 port map( A => n5, ZN => n6);
   U8 : XOR2_X1 port map( A => n6, B => n1, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => n1, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U4 : INV_X1 port map( A => n13, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U2 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U4 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U4 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => B(3), ZN => n2);
   U2 : NAND2_X1 port map( A1 => SEL, A2 => A(3), ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(3));
   U4 : INV_X1 port map( A => SEL, ZN => n1);
   U5 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U6 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U7 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_7;

architecture SYN_STRUCTURAL of carry_select_block_N4_7 is

   component MUX21_GENERIC_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1122, n_1123 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1122);
   RCA1 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1123);
   MUXSUM : MUX21_GENERIC_N4_7 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_6;

architecture SYN_STRUCTURAL of carry_select_block_N4_6 is

   component MUX21_GENERIC_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1124, n_1125 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1124);
   RCA1 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1125);
   MUXSUM : MUX21_GENERIC_N4_6 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_5;

architecture SYN_STRUCTURAL of carry_select_block_N4_5 is

   component MUX21_GENERIC_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1126, n_1127 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1126);
   RCA1 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1127);
   MUXSUM : MUX21_GENERIC_N4_5 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_4;

architecture SYN_STRUCTURAL of carry_select_block_N4_4 is

   component MUX21_GENERIC_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1128, n_1129 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1128);
   RCA1 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1129);
   MUXSUM : MUX21_GENERIC_N4_4 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_3;

architecture SYN_STRUCTURAL of carry_select_block_N4_3 is

   component MUX21_GENERIC_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1130, n_1131 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1130);
   RCA1 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1131);
   MUXSUM : MUX21_GENERIC_N4_3 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_2;

architecture SYN_STRUCTURAL of carry_select_block_N4_2 is

   component MUX21_GENERIC_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1132, n_1133 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1132);
   RCA1 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1133);
   MUXSUM : MUX21_GENERIC_N4_2 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_1;

architecture SYN_STRUCTURAL of carry_select_block_N4_1 is

   component MUX21_GENERIC_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1134, n_1135 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1134);
   RCA1 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1135);
   MUXSUM : MUX21_GENERIC_N4_1 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity BUFF_4 is

   port( IG, IP : in std_logic;  OG, OP : out std_logic);

end BUFF_4;

architecture SYN_BEHAVIORAL of BUFF_4 is

begin
   OG <= IG;
   OP <= IP;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity BUFF_3 is

   port( IG, IP : in std_logic;  OG, OP : out std_logic);

end BUFF_3;

architecture SYN_BEHAVIORAL of BUFF_3 is

begin
   OG <= IG;
   OP <= IP;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity BUFF_2 is

   port( IG, IP : in std_logic;  OG, OP : out std_logic);

end BUFF_2;

architecture SYN_BEHAVIORAL of BUFF_2 is

begin
   OG <= IG;
   OP <= IP;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity BUFF_1 is

   port( IG, IP : in std_logic;  OG, OP : out std_logic);

end BUFF_1;

architecture SYN_BEHAVIORAL of BUFF_1 is

begin
   OG <= IG;
   OP <= IP;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_26 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_26;

architecture SYN_BEHAVIORAL of PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n3);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_25 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_25;

architecture SYN_BEHAVIORAL of PG_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n3);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_24 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_24;

architecture SYN_BEHAVIORAL of PG_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U2 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_23 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_23;

architecture SYN_BEHAVIORAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_22 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_22;

architecture SYN_BEHAVIORAL of PG_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_21 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_21;

architecture SYN_BEHAVIORAL of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_20 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_20;

architecture SYN_BEHAVIORAL of PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_19 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_19;

architecture SYN_BEHAVIORAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_18 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_18;

architecture SYN_BEHAVIORAL of PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => PA, A2 => GA, ZN => n2);
   U2 : NOR2_X1 port map( A1 => GB, A2 => GA, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => G);
   U4 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_17 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_17;

architecture SYN_BEHAVIORAL of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_16 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_16;

architecture SYN_BEHAVIORAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_15 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_15;

architecture SYN_BEHAVIORAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_14 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_14;

architecture SYN_BEHAVIORAL of PG_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U2 : INV_X1 port map( A => n3, ZN => G);
   U3 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_13 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_13;

architecture SYN_BEHAVIORAL of PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U2 : INV_X1 port map( A => n3, ZN => G);
   U3 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_12 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_12;

architecture SYN_BEHAVIORAL of PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n2, A2 => GA, ZN => G);
   U2 : AND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_11 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_11;

architecture SYN_BEHAVIORAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n2, A2 => GA, ZN => G);
   U2 : AND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_10 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_10;

architecture SYN_BEHAVIORAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_9 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_9;

architecture SYN_BEHAVIORAL of PG_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U2 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);
   U3 : INV_X1 port map( A => GA, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_8 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_8;

architecture SYN_BEHAVIORAL of PG_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GA, ZN => n1);
   U2 : NAND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => G);
   U4 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_7 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_7;

architecture SYN_BEHAVIORAL of PG_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GA, ZN => n1);
   U2 : NAND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_6 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_6;

architecture SYN_BEHAVIORAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n3);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_5 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_5;

architecture SYN_BEHAVIORAL of PG_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => GA, ZN => n1);
   U2 : NAND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_4 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_4;

architecture SYN_BEHAVIORAL of PG_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_3 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_3;

architecture SYN_BEHAVIORAL of PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U2 : INV_X1 port map( A => n3, ZN => G);
   U3 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_2 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_2;

architecture SYN_BEHAVIORAL of PG_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => GB, A2 => PA, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => G);
   U3 : AND2_X1 port map( A1 => PA, A2 => PB, ZN => P);
   U4 : INV_X1 port map( A => GA, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_1 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_1;

architecture SYN_BEHAVIORAL of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U3 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_31 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_31;

architecture SYN_behavioral of and_gate_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_30 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_30;

architecture SYN_behavioral of and_gate_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_29 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_29;

architecture SYN_behavioral of and_gate_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_28 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_28;

architecture SYN_behavioral of and_gate_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_27 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_27;

architecture SYN_behavioral of and_gate_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_26 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_26;

architecture SYN_behavioral of and_gate_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_25 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_25;

architecture SYN_behavioral of and_gate_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_24 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_24;

architecture SYN_behavioral of and_gate_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_23 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_23;

architecture SYN_behavioral of and_gate_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_22 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_22;

architecture SYN_behavioral of and_gate_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_21 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_21;

architecture SYN_behavioral of and_gate_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_20 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_20;

architecture SYN_behavioral of and_gate_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_19 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_19;

architecture SYN_behavioral of and_gate_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_18 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_18;

architecture SYN_behavioral of and_gate_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_17 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_17;

architecture SYN_behavioral of and_gate_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_16 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_16;

architecture SYN_behavioral of and_gate_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_15 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_15;

architecture SYN_behavioral of and_gate_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_14 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_14;

architecture SYN_behavioral of and_gate_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_13 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_13;

architecture SYN_behavioral of and_gate_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_12 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_12;

architecture SYN_behavioral of and_gate_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_11 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_11;

architecture SYN_behavioral of and_gate_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_10 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_10;

architecture SYN_behavioral of and_gate_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_9 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_9;

architecture SYN_behavioral of and_gate_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_8 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_8;

architecture SYN_behavioral of and_gate_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_7 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_7;

architecture SYN_behavioral of and_gate_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_6 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_6;

architecture SYN_behavioral of and_gate_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_5 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_5;

architecture SYN_behavioral of and_gate_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_4 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_4;

architecture SYN_behavioral of and_gate_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_3 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_3;

architecture SYN_behavioral of and_gate_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_2 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_2;

architecture SYN_behavioral of and_gate_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_1 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_1;

architecture SYN_behavioral of and_gate_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_31 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_31;

architecture SYN_behavioral of xor_gate_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_30 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_30;

architecture SYN_behavioral of xor_gate_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_29 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_29;

architecture SYN_behavioral of xor_gate_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_28 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_28;

architecture SYN_behavioral of xor_gate_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_27 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_27;

architecture SYN_behavioral of xor_gate_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_26 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_26;

architecture SYN_behavioral of xor_gate_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_25 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_25;

architecture SYN_behavioral of xor_gate_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_24 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_24;

architecture SYN_behavioral of xor_gate_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_23 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_23;

architecture SYN_behavioral of xor_gate_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => O);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_22 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_22;

architecture SYN_behavioral of xor_gate_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_21 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_21;

architecture SYN_behavioral of xor_gate_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_20 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_20;

architecture SYN_behavioral of xor_gate_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_19 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_19;

architecture SYN_behavioral of xor_gate_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_18 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_18;

architecture SYN_behavioral of xor_gate_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_17 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_17;

architecture SYN_behavioral of xor_gate_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => O);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_16 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_16;

architecture SYN_behavioral of xor_gate_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_15 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_15;

architecture SYN_behavioral of xor_gate_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_14 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_14;

architecture SYN_behavioral of xor_gate_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_13 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_13;

architecture SYN_behavioral of xor_gate_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_12 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_12;

architecture SYN_behavioral of xor_gate_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_11 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_11;

architecture SYN_behavioral of xor_gate_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_10 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_10;

architecture SYN_behavioral of xor_gate_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_9 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_9;

architecture SYN_behavioral of xor_gate_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => O);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_8 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_8;

architecture SYN_behavioral of xor_gate_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_7 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_7;

architecture SYN_behavioral of xor_gate_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_6 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_6;

architecture SYN_behavioral of xor_gate_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_5 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_5;

architecture SYN_behavioral of xor_gate_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_4 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_4;

architecture SYN_behavioral of xor_gate_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_3 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_3;

architecture SYN_behavioral of xor_gate_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_2 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_2;

architecture SYN_behavioral of xor_gate_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_1 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_1;

architecture SYN_behavioral of xor_gate_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_9 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_9;

architecture SYN_BEHAVIORAL of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_8 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_8;

architecture SYN_BEHAVIORAL of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_7 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_7;

architecture SYN_BEHAVIORAL of G_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PA, A2 => GB, ZN => n2);
   U2 : OR2_X1 port map( A1 => n2, A2 => GA, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_6 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_6;

architecture SYN_BEHAVIORAL of G_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_5 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_5;

architecture SYN_BEHAVIORAL of G_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X2 port map( A1 => GA, A2 => n2, ZN => G);
   U2 : AND2_X1 port map( A1 => GB, A2 => PA, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_4 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_4;

architecture SYN_BEHAVIORAL of G_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_3 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_3;

architecture SYN_BEHAVIORAL of G_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_2 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_2;

architecture SYN_BEHAVIORAL of G_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NAND2_X2 port map( A1 => n1, A2 => n2, ZN => G);
   U2 : NAND2_X1 port map( A1 => GB, A2 => PA, ZN => n2);
   U3 : INV_X1 port map( A => GA, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_1 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_1;

architecture SYN_BEHAVIORAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FWD_CAM_1 is

   port( RST : in std_logic;  DATA_IN_1, DATA_IN_2, DATA_IN_3 : in 
         std_logic_vector (5 downto 0);  MATCH_1, MATCH_2, MATCH_3 : out 
         std_logic);

end FWD_CAM_1;

architecture SYN_Behavioral of FWD_CAM_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45 : std_logic;

begin
   
   U27 : NAND3_X1 port map( A1 => DATA_IN_3(3), A2 => n42, A3 => DATA_IN_3(4), 
                           ZN => n43);
   U28 : NAND3_X1 port map( A1 => DATA_IN_2(3), A2 => n35, A3 => DATA_IN_2(4), 
                           ZN => n36);
   U29 : NAND3_X1 port map( A1 => DATA_IN_1(3), A2 => n28, A3 => DATA_IN_1(4), 
                           ZN => n29);
   U3 : AND2_X1 port map( A1 => RST, A2 => n31, ZN => MATCH_1);
   U4 : OAI21_X1 port map( B1 => DATA_IN_1(5), B2 => n30, A => n29, ZN => n31);
   U5 : AOI22_X1 port map( A1 => n27, A2 => DATA_IN_1(4), B1 => DATA_IN_1(3), 
                           B2 => n26, ZN => n30);
   U6 : AND2_X1 port map( A1 => RST, A2 => n45, ZN => MATCH_3);
   U7 : OAI21_X1 port map( B1 => DATA_IN_3(5), B2 => n44, A => n43, ZN => n45);
   U8 : AND2_X1 port map( A1 => RST, A2 => n38, ZN => MATCH_2);
   U9 : OAI21_X1 port map( B1 => DATA_IN_2(5), B2 => n37, A => n36, ZN => n38);
   U10 : AND2_X1 port map( A1 => n32, A2 => DATA_IN_2(2), ZN => n34);
   U11 : XNOR2_X1 port map( A => DATA_IN_2(2), B => n2, ZN => n35);
   U12 : AND2_X1 port map( A1 => n39, A2 => DATA_IN_3(2), ZN => n41);
   U13 : XNOR2_X1 port map( A => DATA_IN_3(2), B => n1, ZN => n42);
   U14 : OAI211_X1 port map( C1 => DATA_IN_2(4), C2 => DATA_IN_2(0), A => 
                           DATA_IN_2(2), B => DATA_IN_2(1), ZN => n33);
   U15 : INV_X1 port map( A => DATA_IN_2(1), ZN => n2);
   U16 : OAI211_X1 port map( C1 => DATA_IN_3(4), C2 => DATA_IN_3(0), A => 
                           DATA_IN_3(2), B => DATA_IN_3(1), ZN => n40);
   U17 : INV_X1 port map( A => DATA_IN_3(1), ZN => n1);
   U18 : AOI22_X1 port map( A1 => n41, A2 => DATA_IN_3(4), B1 => DATA_IN_3(3), 
                           B2 => n40, ZN => n44);
   U19 : OAI22_X1 port map( A1 => DATA_IN_3(0), A2 => DATA_IN_3(1), B1 => n1, 
                           B2 => DATA_IN_3(3), ZN => n39);
   U20 : INV_X1 port map( A => DATA_IN_1(1), ZN => n3);
   U21 : OAI22_X1 port map( A1 => DATA_IN_1(0), A2 => DATA_IN_1(1), B1 => n3, 
                           B2 => DATA_IN_1(3), ZN => n25);
   U22 : AOI22_X1 port map( A1 => n34, A2 => DATA_IN_2(4), B1 => DATA_IN_2(3), 
                           B2 => n33, ZN => n37);
   U23 : OAI22_X1 port map( A1 => DATA_IN_2(0), A2 => DATA_IN_2(1), B1 => n2, 
                           B2 => DATA_IN_2(3), ZN => n32);
   U24 : AND2_X1 port map( A1 => n25, A2 => DATA_IN_1(2), ZN => n27);
   U25 : OAI211_X1 port map( C1 => DATA_IN_1(4), C2 => DATA_IN_1(0), A => 
                           DATA_IN_1(2), B => DATA_IN_1(1), ZN => n26);
   U26 : XNOR2_X1 port map( A => DATA_IN_1(2), B => n3, ZN => n28);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity mux_3to1_N32_3 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux_3to1_N32_3;

architecture SYN_BEHAVIORAL of mux_3to1_N32_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27986, net28019, net29531, net29543, net29814, net37145, net37292,
      net37339, net37338, net37714, net37887, net37925, net37961, net38041, 
      net38078, net38213, net38721, net38782, net38796, net39109, net43925, 
      net28020, net45622, net37351, net37209, net28024, n3, n6, n7, n8, n9, n10
      , n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n28, n29, n30, n31, n32, n33, n35, n36, n37, n40, n41, n42, n45, n46
      , n47, n50, n51, n52, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, 
      n66, n67, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105 : std_logic;

begin
   
   U1 : OR3_X2 port map( A1 => n35, A2 => n37, A3 => n36, ZN => Y(18));
   U2 : NAND3_X2 port map( A1 => n14, A2 => n15, A3 => n16, ZN => Y(23));
   U3 : CLKBUF_X1 port map( A => net27986, Z => net29543);
   U4 : CLKBUF_X1 port map( A => net27986, Z => net37714);
   U5 : NAND3_X1 port map( A1 => n54, A2 => n55, A3 => n56, ZN => Y(22));
   U6 : OR3_X1 port map( A1 => n17, A2 => n18, A3 => n19, ZN => Y(25));
   U7 : BUF_X1 port map( A => net27986, Z => net43925);
   U8 : CLKBUF_X1 port map( A => SEL(0), Z => net37351);
   U9 : CLKBUF_X1 port map( A => net28019, Z => net38721);
   U10 : OR3_X2 port map( A1 => n50, A2 => n51, A3 => n52, ZN => Y(21));
   U11 : CLKBUF_X1 port map( A => net37145, Z => n3);
   U12 : CLKBUF_X1 port map( A => net37145, Z => net37887);
   U13 : NAND3_X1 port map( A1 => n74, A2 => n75, A3 => n76, ZN => Y(17));
   U14 : NAND2_X1 port map( A1 => SEL(1), A2 => n6, ZN => net28019);
   U15 : INV_X1 port map( A => SEL(0), ZN => n6);
   U16 : INV_X1 port map( A => SEL(1), ZN => net28024);
   U17 : NAND3_X1 port map( A1 => n8, A2 => n7, A3 => n9, ZN => Y(0));
   U18 : NAND2_X1 port map( A1 => net27986, A2 => C(0), ZN => n9);
   U19 : INV_X1 port map( A => net28019, ZN => net27986);
   U20 : NAND2_X1 port map( A1 => B(0), A2 => net29814, ZN => n7);
   U21 : OR2_X1 port map( A1 => n10, A2 => net29814, ZN => n8);
   U22 : NAND2_X1 port map( A1 => net37209, A2 => A(0), ZN => n10);
   U23 : BUF_X1 port map( A => net28019, Z => net37209);
   U24 : INV_X1 port map( A => net37209, ZN => net37292);
   U25 : AND2_X1 port map( A1 => net28024, A2 => net37351, ZN => net29814);
   U26 : AND2_X2 port map( A1 => net28024, A2 => net37351, ZN => net37925);
   U27 : NAND2_X1 port map( A1 => net28024, A2 => net37351, ZN => net28020);
   U28 : INV_X1 port map( A => net38721, ZN => net45622);
   U29 : INV_X1 port map( A => net38721, ZN => net38796);
   U30 : OR3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => Y(19));
   U31 : AND2_X2 port map( A1 => net28020, A2 => net28019, ZN => net37145);
   U32 : AND2_X2 port map( A1 => net28019, A2 => net28020, ZN => net38041);
   U33 : OR3_X2 port map( A1 => n12, A2 => n11, A3 => n13, ZN => Y(14));
   U34 : AND2_X1 port map( A1 => net27986, A2 => C(14), ZN => n13);
   U35 : AND2_X1 port map( A1 => B(14), A2 => net29814, ZN => n11);
   U36 : AND2_X1 port map( A1 => net37145, A2 => A(14), ZN => n12);
   U37 : CLKBUF_X1 port map( A => net37145, Z => net39109);
   U38 : NAND2_X1 port map( A1 => B(23), A2 => net37961, ZN => n14);
   U39 : NAND2_X1 port map( A1 => A(23), A2 => net37887, ZN => n15);
   U40 : NAND2_X1 port map( A1 => C(23), A2 => net37714, ZN => n16);
   U41 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => Y(13));
   U42 : AND2_X1 port map( A1 => B(25), A2 => net37961, ZN => n17);
   U43 : AND2_X1 port map( A1 => A(25), A2 => net37887, ZN => n18);
   U44 : AND2_X1 port map( A1 => C(25), A2 => net29543, ZN => n19);
   U45 : BUF_X1 port map( A => net29814, Z => net37961);
   U46 : NAND3_X1 port map( A1 => n78, A2 => n77, A3 => n79, ZN => Y(3));
   U47 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => Y(15));
   U48 : NAND2_X1 port map( A1 => net39109, A2 => A(15), ZN => n20);
   U49 : NAND2_X1 port map( A1 => net43925, A2 => C(15), ZN => n21);
   U50 : NAND2_X1 port map( A1 => B(15), A2 => net29814, ZN => n22);
   U51 : NAND3_X1 port map( A1 => n91, A2 => n90, A3 => n92, ZN => Y(8));
   U52 : NAND3_X1 port map( A1 => n23, A2 => n24, A3 => n25, ZN => Y(11));
   U53 : NAND2_X1 port map( A1 => net38041, A2 => A(11), ZN => n23);
   U54 : NAND2_X1 port map( A1 => net43925, A2 => C(11), ZN => n24);
   U55 : NAND2_X1 port map( A1 => net29814, A2 => B(11), ZN => n25);
   U56 : CLKBUF_X1 port map( A => net37145, Z => net38782);
   U57 : NAND3_X1 port map( A1 => n40, A2 => n41, A3 => n42, ZN => Y(12));
   U58 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => Y(7));
   U59 : NAND2_X1 port map( A1 => net38041, A2 => A(7), ZN => n28);
   U60 : NAND2_X1 port map( A1 => net38796, A2 => C(7), ZN => n29);
   U61 : NAND2_X1 port map( A1 => B(7), A2 => net37925, ZN => n30);
   U62 : CLKBUF_X1 port map( A => net29543, Z => net38213);
   U63 : CLKBUF_X1 port map( A => net37145, Z => net38078);
   U64 : NAND2_X1 port map( A1 => B(20), A2 => net37961, ZN => n31);
   U65 : NAND2_X1 port map( A1 => A(20), A2 => net38078, ZN => n32);
   U66 : NAND2_X1 port map( A1 => C(20), A2 => net37292, ZN => n33);
   U67 : AND3_X1 port map( A1 => n31, A2 => n32, A3 => n33, ZN => n98);
   U68 : CLKBUF_X1 port map( A => net37925, Z => net29531);
   U69 : AND2_X1 port map( A1 => B(18), A2 => net37925, ZN => n35);
   U70 : AND2_X1 port map( A1 => net37145, A2 => A(18), ZN => n36);
   U71 : AND2_X1 port map( A1 => net27986, A2 => C(18), ZN => n37);
   U72 : NAND3_X1 port map( A1 => n82, A2 => n81, A3 => n80, ZN => Y(2));
   U73 : INV_X1 port map( A => net37338, ZN => net37339);
   U74 : NAND2_X1 port map( A1 => B(12), A2 => net37925, ZN => n40);
   U75 : NAND2_X1 port map( A1 => net38041, A2 => A(12), ZN => n41);
   U76 : NAND2_X1 port map( A1 => net37292, A2 => C(12), ZN => n42);
   U77 : NAND3_X1 port map( A1 => n87, A2 => n88, A3 => n89, ZN => Y(10));
   U78 : AND2_X1 port map( A1 => B(19), A2 => net37925, ZN => n45);
   U79 : AND2_X1 port map( A1 => net37145, A2 => A(19), ZN => n46);
   U80 : AND2_X1 port map( A1 => net27986, A2 => C(19), ZN => n47);
   U81 : NAND3_X1 port map( A1 => n57, A2 => n58, A3 => n59, ZN => Y(4));
   U82 : AND2_X1 port map( A1 => B(21), A2 => net37925, ZN => n50);
   U83 : AND2_X1 port map( A1 => n3, A2 => A(21), ZN => n51);
   U84 : AND2_X1 port map( A1 => C(21), A2 => net37292, ZN => n52);
   U85 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => Y(5));
   U86 : NAND2_X1 port map( A1 => B(22), A2 => net37961, ZN => n54);
   U87 : NAND2_X1 port map( A1 => A(22), A2 => net37887, ZN => n55);
   U88 : NAND2_X1 port map( A1 => C(22), A2 => net37714, ZN => n56);
   U89 : NAND3_X1 port map( A1 => n94, A2 => n95, A3 => n96, ZN => Y(1));
   U90 : NAND2_X1 port map( A1 => B(4), A2 => net37925, ZN => n57);
   U91 : NAND2_X1 port map( A1 => net38041, A2 => A(4), ZN => n58);
   U92 : NAND2_X1 port map( A1 => C(4), A2 => net45622, ZN => n59);
   U93 : NAND3_X1 port map( A1 => n83, A2 => n84, A3 => n85, ZN => Y(9));
   U94 : NAND3_X1 port map( A1 => n65, A2 => n66, A3 => n67, ZN => Y(6));
   U95 : NAND2_X1 port map( A1 => net37925, A2 => B(5), ZN => n62);
   U96 : NAND2_X1 port map( A1 => net38041, A2 => A(5), ZN => n63);
   U97 : NAND2_X1 port map( A1 => net38796, A2 => C(5), ZN => n64);
   U98 : NAND2_X1 port map( A1 => B(6), A2 => net37925, ZN => n65);
   U99 : NAND2_X1 port map( A1 => net38041, A2 => A(6), ZN => n66);
   U100 : NAND2_X1 port map( A1 => net37292, A2 => C(6), ZN => n67);
   U101 : NAND2_X1 port map( A1 => B(13), A2 => net37925, ZN => n71);
   U102 : NAND2_X1 port map( A1 => net38041, A2 => A(13), ZN => n72);
   U103 : NAND2_X1 port map( A1 => C(13), A2 => net37292, ZN => n73);
   U104 : NAND2_X1 port map( A1 => B(17), A2 => net37925, ZN => n74);
   U105 : NAND2_X1 port map( A1 => n3, A2 => A(17), ZN => n75);
   U106 : NAND2_X1 port map( A1 => C(17), A2 => net38796, ZN => n76);
   U107 : NAND2_X1 port map( A1 => B(3), A2 => net29814, ZN => n77);
   U108 : NAND2_X1 port map( A1 => net38041, A2 => A(3), ZN => n78);
   U109 : NAND2_X1 port map( A1 => net38796, A2 => C(3), ZN => n79);
   U110 : INV_X1 port map( A => net38041, ZN => net37338);
   U111 : NAND2_X1 port map( A1 => net37925, A2 => B(2), ZN => n80);
   U112 : NAND2_X1 port map( A1 => net37145, A2 => A(2), ZN => n81);
   U113 : NAND2_X1 port map( A1 => net45622, A2 => C(2), ZN => n82);
   U114 : NAND2_X1 port map( A1 => B(9), A2 => net37925, ZN => n83);
   U115 : NAND2_X1 port map( A1 => net37145, A2 => A(9), ZN => n84);
   U116 : NAND2_X1 port map( A1 => net27986, A2 => C(9), ZN => n85);
   U117 : NAND2_X1 port map( A1 => B(10), A2 => net37925, ZN => n87);
   U118 : NAND2_X1 port map( A1 => net38041, A2 => A(10), ZN => n88);
   U119 : NAND2_X1 port map( A1 => C(10), A2 => net45622, ZN => n89);
   U120 : NAND2_X1 port map( A1 => B(8), A2 => net37925, ZN => n90);
   U121 : NAND2_X1 port map( A1 => net38041, A2 => A(8), ZN => n91);
   U122 : NAND2_X1 port map( A1 => net37292, A2 => C(8), ZN => n92);
   U123 : NAND2_X1 port map( A1 => B(1), A2 => net37925, ZN => n94);
   U124 : NAND2_X1 port map( A1 => net37145, A2 => A(1), ZN => n95);
   U125 : NAND2_X1 port map( A1 => C(1), A2 => net27986, ZN => n96);
   U126 : AOI222_X1 port map( A1 => B(16), A2 => net37925, B1 => net38782, B2 
                           => A(16), C1 => net37714, C2 => C(16), ZN => n97);
   U127 : INV_X1 port map( A => n97, ZN => Y(16));
   U128 : INV_X1 port map( A => n98, ZN => Y(20));
   U129 : AOI222_X1 port map( A1 => B(24), A2 => net29531, B1 => A(24), B2 => 
                           net37339, C1 => C(24), C2 => net29543, ZN => n99);
   U130 : INV_X1 port map( A => n99, ZN => Y(24));
   U131 : AOI222_X1 port map( A1 => B(26), A2 => net37961, B1 => A(26), B2 => 
                           net37339, C1 => C(26), C2 => net29543, ZN => n100);
   U132 : INV_X1 port map( A => n100, ZN => Y(26));
   U133 : AOI222_X1 port map( A1 => B(27), A2 => net29531, B1 => A(27), B2 => 
                           net37339, C1 => C(27), C2 => net29543, ZN => n101);
   U134 : INV_X1 port map( A => n101, ZN => Y(27));
   U135 : AOI222_X1 port map( A1 => B(28), A2 => net29531, B1 => A(28), B2 => 
                           net37339, C1 => C(28), C2 => net29543, ZN => n102);
   U136 : INV_X1 port map( A => n102, ZN => Y(28));
   U137 : AOI222_X1 port map( A1 => B(29), A2 => net29531, B1 => A(29), B2 => 
                           net37339, C1 => C(29), C2 => net38213, ZN => n103);
   U138 : INV_X1 port map( A => n103, ZN => Y(29));
   U139 : AOI222_X1 port map( A1 => B(30), A2 => net29531, B1 => A(30), B2 => 
                           net37339, C1 => C(30), C2 => net29543, ZN => n104);
   U140 : INV_X1 port map( A => n104, ZN => Y(30));
   U141 : AOI222_X1 port map( A1 => B(31), A2 => net29531, B1 => A(31), B2 => 
                           net37339, C1 => C(31), C2 => net38213, ZN => n105);
   U142 : INV_X1 port map( A => n105, ZN => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity mux_3to1_N32_2 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux_3to1_N32_2;

architecture SYN_BEHAVIORAL of mux_3to1_N32_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n109, Z => n1);
   U2 : BUF_X1 port map( A => n109, Z => n2);
   U3 : BUF_X1 port map( A => n109, Z => n3);
   U4 : NOR2_X1 port map( A1 => n6, A2 => n7, ZN => n109);
   U5 : INV_X1 port map( A => n93, ZN => Y(23));
   U6 : INV_X1 port map( A => n92, ZN => Y(22));
   U7 : INV_X1 port map( A => n91, ZN => Y(21));
   U8 : INV_X1 port map( A => n112, ZN => Y(9));
   U9 : INV_X1 port map( A => n108, ZN => Y(8));
   U10 : INV_X1 port map( A => n107, ZN => Y(7));
   U11 : INV_X1 port map( A => n89, ZN => Y(1));
   U12 : INV_X1 port map( A => n88, ZN => Y(19));
   U13 : INV_X1 port map( A => n87, ZN => Y(18));
   U14 : INV_X1 port map( A => n105, ZN => Y(5));
   U15 : INV_X1 port map( A => n104, ZN => Y(4));
   U16 : INV_X1 port map( A => n103, ZN => Y(3));
   U17 : INV_X1 port map( A => n85, ZN => Y(16));
   U18 : INV_X1 port map( A => n84, ZN => Y(15));
   U19 : INV_X1 port map( A => n83, ZN => Y(14));
   U20 : INV_X1 port map( A => n101, ZN => Y(30));
   U21 : INV_X1 port map( A => n100, ZN => Y(2));
   U22 : INV_X1 port map( A => n99, ZN => Y(29));
   U23 : INV_X1 port map( A => n81, ZN => Y(12));
   U24 : INV_X1 port map( A => n80, ZN => Y(11));
   U25 : INV_X1 port map( A => n79, ZN => Y(10));
   U26 : INV_X1 port map( A => n97, ZN => Y(27));
   U27 : INV_X1 port map( A => n96, ZN => Y(26));
   U28 : INV_X1 port map( A => n95, ZN => Y(25));
   U29 : BUF_X1 port map( A => n110, Z => n6);
   U30 : BUF_X1 port map( A => n110, Z => n4);
   U31 : BUF_X1 port map( A => n110, Z => n5);
   U32 : BUF_X1 port map( A => n111, Z => n9);
   U33 : BUF_X1 port map( A => n111, Z => n7);
   U34 : BUF_X1 port map( A => n111, Z => n8);
   U35 : AOI222_X1 port map( A1 => B(14), A2 => n7, B1 => C(14), B2 => n6, C1 
                           => A(14), C2 => n1, ZN => n83);
   U36 : AOI222_X1 port map( A1 => B(15), A2 => n7, B1 => C(15), B2 => n6, C1 
                           => A(15), C2 => n1, ZN => n84);
   U37 : AOI222_X1 port map( A1 => B(16), A2 => n7, B1 => C(16), B2 => n6, C1 
                           => A(16), C2 => n1, ZN => n85);
   U38 : AOI222_X1 port map( A1 => B(10), A2 => n7, B1 => C(10), B2 => n6, C1 
                           => A(10), C2 => n1, ZN => n79);
   U39 : AOI222_X1 port map( A1 => B(11), A2 => n7, B1 => C(11), B2 => n6, C1 
                           => A(11), C2 => n1, ZN => n80);
   U40 : AOI222_X1 port map( A1 => B(12), A2 => n7, B1 => C(12), B2 => n6, C1 
                           => A(12), C2 => n1, ZN => n81);
   U41 : AOI222_X1 port map( A1 => B(21), A2 => n8, B1 => C(21), B2 => n5, C1 
                           => A(21), C2 => n2, ZN => n91);
   U42 : AOI222_X1 port map( A1 => B(22), A2 => n8, B1 => C(22), B2 => n5, C1 
                           => A(22), C2 => n2, ZN => n92);
   U43 : AOI222_X1 port map( A1 => B(23), A2 => n8, B1 => C(23), B2 => n5, C1 
                           => A(23), C2 => n2, ZN => n93);
   U44 : AOI222_X1 port map( A1 => B(18), A2 => n7, B1 => C(18), B2 => n5, C1 
                           => A(18), C2 => n1, ZN => n87);
   U45 : AOI222_X1 port map( A1 => B(19), A2 => n7, B1 => C(19), B2 => n5, C1 
                           => A(19), C2 => n1, ZN => n88);
   U46 : AOI222_X1 port map( A1 => B(1), A2 => n8, B1 => C(1), B2 => n5, C1 => 
                           A(1), C2 => n1, ZN => n89);
   U47 : AOI222_X1 port map( A1 => B(7), A2 => n9, B1 => C(7), B2 => n4, C1 => 
                           A(7), C2 => n3, ZN => n107);
   U48 : AOI222_X1 port map( A1 => B(8), A2 => n9, B1 => C(8), B2 => n4, C1 => 
                           A(8), C2 => n3, ZN => n108);
   U49 : AOI222_X1 port map( A1 => B(9), A2 => n9, B1 => C(9), B2 => n4, C1 => 
                           A(9), C2 => n3, ZN => n112);
   U50 : AOI222_X1 port map( A1 => B(3), A2 => n9, B1 => C(3), B2 => n4, C1 => 
                           A(3), C2 => n3, ZN => n103);
   U51 : AOI222_X1 port map( A1 => B(4), A2 => n9, B1 => C(4), B2 => n4, C1 => 
                           A(4), C2 => n3, ZN => n104);
   U52 : AOI222_X1 port map( A1 => B(5), A2 => n9, B1 => C(5), B2 => n4, C1 => 
                           A(5), C2 => n3, ZN => n105);
   U53 : AOI222_X1 port map( A1 => B(29), A2 => n8, B1 => C(29), B2 => n4, C1 
                           => A(29), C2 => n2, ZN => n99);
   U54 : AOI222_X1 port map( A1 => B(2), A2 => n8, B1 => C(2), B2 => n4, C1 => 
                           A(2), C2 => n2, ZN => n100);
   U55 : AOI222_X1 port map( A1 => B(30), A2 => n9, B1 => C(30), B2 => n4, C1 
                           => A(30), C2 => n2, ZN => n101);
   U56 : AOI222_X1 port map( A1 => B(25), A2 => n8, B1 => C(25), B2 => n5, C1 
                           => A(25), C2 => n2, ZN => n95);
   U57 : AOI222_X1 port map( A1 => B(26), A2 => n8, B1 => C(26), B2 => n5, C1 
                           => A(26), C2 => n2, ZN => n96);
   U58 : AOI222_X1 port map( A1 => B(27), A2 => n8, B1 => C(27), B2 => n5, C1 
                           => A(27), C2 => n2, ZN => n97);
   U59 : INV_X1 port map( A => n86, ZN => Y(17));
   U60 : AOI222_X1 port map( A1 => B(17), A2 => n7, B1 => C(17), B2 => n5, C1 
                           => A(17), C2 => n1, ZN => n86);
   U61 : INV_X1 port map( A => n98, ZN => Y(28));
   U62 : AOI222_X1 port map( A1 => B(28), A2 => n8, B1 => C(28), B2 => n4, C1 
                           => A(28), C2 => n2, ZN => n98);
   U63 : INV_X1 port map( A => n94, ZN => Y(24));
   U64 : AOI222_X1 port map( A1 => B(24), A2 => n8, B1 => C(24), B2 => n5, C1 
                           => A(24), C2 => n2, ZN => n94);
   U65 : INV_X1 port map( A => n82, ZN => Y(13));
   U66 : AOI222_X1 port map( A1 => B(13), A2 => n7, B1 => C(13), B2 => n6, C1 
                           => A(13), C2 => n1, ZN => n82);
   U67 : INV_X1 port map( A => n78, ZN => Y(0));
   U68 : AOI222_X1 port map( A1 => B(0), A2 => n7, B1 => C(0), B2 => n6, C1 => 
                           A(0), C2 => n1, ZN => n78);
   U69 : INV_X1 port map( A => n90, ZN => Y(20));
   U70 : AOI222_X1 port map( A1 => B(20), A2 => n8, B1 => C(20), B2 => n5, C1 
                           => A(20), C2 => n2, ZN => n90);
   U71 : INV_X1 port map( A => n106, ZN => Y(6));
   U72 : AOI222_X1 port map( A1 => B(6), A2 => n9, B1 => C(6), B2 => n4, C1 => 
                           A(6), C2 => n3, ZN => n106);
   U73 : INV_X1 port map( A => n102, ZN => Y(31));
   U74 : AOI222_X1 port map( A1 => B(31), A2 => n9, B1 => C(31), B2 => n4, C1 
                           => A(31), C2 => n3, ZN => n102);
   U75 : NOR2_X1 port map( A1 => n77, A2 => SEL(1), ZN => n111);
   U76 : AND2_X1 port map( A1 => SEL(1), A2 => n77, ZN => n110);
   U77 : INV_X1 port map( A => SEL(0), ZN => n77);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity mux_3to1_N32_1 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux_3to1_N32_1;

architecture SYN_BEHAVIORAL of mux_3to1_N32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n109, Z => n1);
   U2 : BUF_X1 port map( A => n109, Z => n2);
   U3 : BUF_X1 port map( A => n109, Z => n3);
   U4 : NOR2_X1 port map( A1 => n6, A2 => n7, ZN => n109);
   U5 : BUF_X1 port map( A => n110, Z => n6);
   U6 : BUF_X1 port map( A => n110, Z => n5);
   U7 : BUF_X1 port map( A => n110, Z => n4);
   U8 : BUF_X1 port map( A => n111, Z => n9);
   U9 : BUF_X1 port map( A => n111, Z => n7);
   U10 : BUF_X1 port map( A => n111, Z => n8);
   U11 : NOR2_X1 port map( A1 => n77, A2 => SEL(1), ZN => n111);
   U12 : AND2_X1 port map( A1 => SEL(1), A2 => n77, ZN => n110);
   U13 : INV_X1 port map( A => n78, ZN => Y(0));
   U14 : AOI222_X1 port map( A1 => B(0), A2 => n7, B1 => C(0), B2 => n6, C1 => 
                           A(0), C2 => n1, ZN => n78);
   U15 : INV_X1 port map( A => n89, ZN => Y(1));
   U16 : AOI222_X1 port map( A1 => B(1), A2 => n8, B1 => C(1), B2 => n5, C1 => 
                           A(1), C2 => n1, ZN => n89);
   U17 : INV_X1 port map( A => n100, ZN => Y(2));
   U18 : AOI222_X1 port map( A1 => B(2), A2 => n8, B1 => C(2), B2 => n4, C1 => 
                           A(2), C2 => n2, ZN => n100);
   U19 : INV_X1 port map( A => n103, ZN => Y(3));
   U20 : AOI222_X1 port map( A1 => B(3), A2 => n9, B1 => C(3), B2 => n4, C1 => 
                           A(3), C2 => n3, ZN => n103);
   U21 : INV_X1 port map( A => n104, ZN => Y(4));
   U22 : AOI222_X1 port map( A1 => B(4), A2 => n9, B1 => C(4), B2 => n4, C1 => 
                           A(4), C2 => n3, ZN => n104);
   U23 : INV_X1 port map( A => n105, ZN => Y(5));
   U24 : AOI222_X1 port map( A1 => B(5), A2 => n9, B1 => C(5), B2 => n4, C1 => 
                           A(5), C2 => n3, ZN => n105);
   U25 : INV_X1 port map( A => n106, ZN => Y(6));
   U26 : AOI222_X1 port map( A1 => B(6), A2 => n9, B1 => C(6), B2 => n4, C1 => 
                           A(6), C2 => n3, ZN => n106);
   U27 : INV_X1 port map( A => n107, ZN => Y(7));
   U28 : AOI222_X1 port map( A1 => B(7), A2 => n9, B1 => C(7), B2 => n4, C1 => 
                           A(7), C2 => n3, ZN => n107);
   U29 : INV_X1 port map( A => n108, ZN => Y(8));
   U30 : AOI222_X1 port map( A1 => B(8), A2 => n9, B1 => C(8), B2 => n4, C1 => 
                           A(8), C2 => n3, ZN => n108);
   U31 : INV_X1 port map( A => n112, ZN => Y(9));
   U32 : AOI222_X1 port map( A1 => B(9), A2 => n9, B1 => C(9), B2 => n4, C1 => 
                           A(9), C2 => n3, ZN => n112);
   U33 : INV_X1 port map( A => n79, ZN => Y(10));
   U34 : AOI222_X1 port map( A1 => B(10), A2 => n7, B1 => C(10), B2 => n6, C1 
                           => A(10), C2 => n1, ZN => n79);
   U35 : INV_X1 port map( A => n80, ZN => Y(11));
   U36 : AOI222_X1 port map( A1 => B(11), A2 => n7, B1 => C(11), B2 => n6, C1 
                           => A(11), C2 => n1, ZN => n80);
   U37 : INV_X1 port map( A => n81, ZN => Y(12));
   U38 : AOI222_X1 port map( A1 => B(12), A2 => n7, B1 => C(12), B2 => n6, C1 
                           => A(12), C2 => n1, ZN => n81);
   U39 : INV_X1 port map( A => n82, ZN => Y(13));
   U40 : AOI222_X1 port map( A1 => B(13), A2 => n7, B1 => C(13), B2 => n6, C1 
                           => A(13), C2 => n1, ZN => n82);
   U41 : INV_X1 port map( A => n83, ZN => Y(14));
   U42 : AOI222_X1 port map( A1 => B(14), A2 => n7, B1 => C(14), B2 => n6, C1 
                           => A(14), C2 => n1, ZN => n83);
   U43 : INV_X1 port map( A => n84, ZN => Y(15));
   U44 : AOI222_X1 port map( A1 => B(15), A2 => n7, B1 => C(15), B2 => n6, C1 
                           => A(15), C2 => n1, ZN => n84);
   U45 : INV_X1 port map( A => n85, ZN => Y(16));
   U46 : AOI222_X1 port map( A1 => B(16), A2 => n7, B1 => C(16), B2 => n6, C1 
                           => A(16), C2 => n1, ZN => n85);
   U47 : INV_X1 port map( A => n86, ZN => Y(17));
   U48 : AOI222_X1 port map( A1 => B(17), A2 => n7, B1 => C(17), B2 => n5, C1 
                           => A(17), C2 => n1, ZN => n86);
   U49 : INV_X1 port map( A => n87, ZN => Y(18));
   U50 : AOI222_X1 port map( A1 => B(18), A2 => n7, B1 => C(18), B2 => n5, C1 
                           => A(18), C2 => n1, ZN => n87);
   U51 : INV_X1 port map( A => n88, ZN => Y(19));
   U52 : AOI222_X1 port map( A1 => B(19), A2 => n7, B1 => C(19), B2 => n5, C1 
                           => A(19), C2 => n1, ZN => n88);
   U53 : INV_X1 port map( A => n90, ZN => Y(20));
   U54 : AOI222_X1 port map( A1 => B(20), A2 => n8, B1 => C(20), B2 => n5, C1 
                           => A(20), C2 => n2, ZN => n90);
   U55 : INV_X1 port map( A => n91, ZN => Y(21));
   U56 : AOI222_X1 port map( A1 => B(21), A2 => n8, B1 => C(21), B2 => n5, C1 
                           => A(21), C2 => n2, ZN => n91);
   U57 : INV_X1 port map( A => n92, ZN => Y(22));
   U58 : AOI222_X1 port map( A1 => B(22), A2 => n8, B1 => C(22), B2 => n5, C1 
                           => A(22), C2 => n2, ZN => n92);
   U59 : INV_X1 port map( A => n93, ZN => Y(23));
   U60 : AOI222_X1 port map( A1 => B(23), A2 => n8, B1 => C(23), B2 => n5, C1 
                           => A(23), C2 => n2, ZN => n93);
   U61 : INV_X1 port map( A => n94, ZN => Y(24));
   U62 : AOI222_X1 port map( A1 => B(24), A2 => n8, B1 => C(24), B2 => n5, C1 
                           => A(24), C2 => n2, ZN => n94);
   U63 : INV_X1 port map( A => n95, ZN => Y(25));
   U64 : AOI222_X1 port map( A1 => B(25), A2 => n8, B1 => C(25), B2 => n5, C1 
                           => A(25), C2 => n2, ZN => n95);
   U65 : INV_X1 port map( A => n96, ZN => Y(26));
   U66 : AOI222_X1 port map( A1 => B(26), A2 => n8, B1 => C(26), B2 => n5, C1 
                           => A(26), C2 => n2, ZN => n96);
   U67 : INV_X1 port map( A => n97, ZN => Y(27));
   U68 : AOI222_X1 port map( A1 => B(27), A2 => n8, B1 => C(27), B2 => n5, C1 
                           => A(27), C2 => n2, ZN => n97);
   U69 : INV_X1 port map( A => n98, ZN => Y(28));
   U70 : AOI222_X1 port map( A1 => B(28), A2 => n8, B1 => C(28), B2 => n4, C1 
                           => A(28), C2 => n2, ZN => n98);
   U71 : INV_X1 port map( A => n99, ZN => Y(29));
   U72 : AOI222_X1 port map( A1 => B(29), A2 => n8, B1 => C(29), B2 => n4, C1 
                           => A(29), C2 => n2, ZN => n99);
   U73 : INV_X1 port map( A => n101, ZN => Y(30));
   U74 : AOI222_X1 port map( A1 => B(30), A2 => n9, B1 => C(30), B2 => n4, C1 
                           => A(30), C2 => n2, ZN => n101);
   U75 : INV_X1 port map( A => n102, ZN => Y(31));
   U76 : AOI222_X1 port map( A1 => B(31), A2 => n9, B1 => C(31), B2 => n4, C1 
                           => A(31), C2 => n3, ZN => n102);
   U77 : INV_X1 port map( A => SEL(0), ZN => n77);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N32_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n10, Z => n3);
   U2 : BUF_X1 port map( A => n10, Z => n2);
   U3 : BUF_X1 port map( A => n10, Z => n8);
   U4 : BUF_X1 port map( A => n8, Z => n7);
   U5 : BUF_X1 port map( A => n9, Z => n6);
   U6 : BUF_X1 port map( A => n3, Z => n5);
   U7 : BUF_X1 port map( A => n10, Z => n4);
   U8 : BUF_X1 port map( A => n10, Z => n9);
   U9 : INV_X1 port map( A => n1, ZN => n10);
   U10 : BUF_X1 port map( A => SEL, Z => n1);
   U11 : INV_X1 port map( A => n97, ZN => Y(2));
   U12 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n4, ZN => 
                           n97);
   U13 : INV_X1 port map( A => n103, ZN => Y(6));
   U14 : AOI22_X1 port map( A1 => A(6), A2 => SEL, B1 => B(6), B2 => n2, ZN => 
                           n103);
   U15 : INV_X1 port map( A => n102, ZN => Y(5));
   U16 : AOI22_X1 port map( A1 => A(5), A2 => n1, B1 => B(5), B2 => n3, ZN => 
                           n102);
   U17 : INV_X1 port map( A => n101, ZN => Y(4));
   U18 : AOI22_X1 port map( A1 => A(4), A2 => SEL, B1 => B(4), B2 => n3, ZN => 
                           n101);
   U19 : INV_X1 port map( A => n106, ZN => Y(9));
   U20 : AOI22_X1 port map( A1 => n1, A2 => A(9), B1 => B(9), B2 => n2, ZN => 
                           n106);
   U21 : INV_X1 port map( A => n77, ZN => Y(11));
   U22 : AOI22_X1 port map( A1 => A(11), A2 => SEL, B1 => B(11), B2 => n9, ZN 
                           => n77);
   U23 : INV_X1 port map( A => n80, ZN => Y(14));
   U24 : AOI22_X1 port map( A1 => A(14), A2 => n1, B1 => B(14), B2 => n8, ZN =>
                           n80);
   U25 : INV_X1 port map( A => n83, ZN => Y(17));
   U26 : AOI22_X1 port map( A1 => A(17), A2 => SEL, B1 => B(17), B2 => n7, ZN 
                           => n83);
   U27 : INV_X1 port map( A => n89, ZN => Y(22));
   U28 : AOI22_X1 port map( A1 => A(22), A2 => n1, B1 => B(22), B2 => n6, ZN =>
                           n89);
   U29 : INV_X1 port map( A => n92, ZN => Y(25));
   U30 : AOI22_X1 port map( A1 => A(25), A2 => n1, B1 => B(25), B2 => n5, ZN =>
                           n92);
   U31 : INV_X1 port map( A => n95, ZN => Y(28));
   U32 : AOI22_X1 port map( A1 => A(28), A2 => n1, B1 => B(28), B2 => n4, ZN =>
                           n95);
   U33 : INV_X1 port map( A => n88, ZN => Y(21));
   U34 : AOI22_X1 port map( A1 => A(21), A2 => n1, B1 => B(21), B2 => n6, ZN =>
                           n88);
   U35 : INV_X1 port map( A => n79, ZN => Y(13));
   U36 : AOI22_X1 port map( A1 => A(13), A2 => n1, B1 => B(13), B2 => n8, ZN =>
                           n79);
   U37 : INV_X1 port map( A => n82, ZN => Y(16));
   U38 : AOI22_X1 port map( A1 => A(16), A2 => SEL, B1 => B(16), B2 => n8, ZN 
                           => n82);
   U39 : INV_X1 port map( A => n85, ZN => Y(19));
   U40 : AOI22_X1 port map( A1 => A(19), A2 => n1, B1 => B(19), B2 => n7, ZN =>
                           n85);
   U41 : INV_X1 port map( A => n91, ZN => Y(24));
   U42 : AOI22_X1 port map( A1 => A(24), A2 => n1, B1 => B(24), B2 => n5, ZN =>
                           n91);
   U43 : INV_X1 port map( A => n94, ZN => Y(27));
   U44 : AOI22_X1 port map( A1 => A(27), A2 => n1, B1 => B(27), B2 => n5, ZN =>
                           n94);
   U45 : INV_X1 port map( A => n98, ZN => Y(30));
   U46 : AOI22_X1 port map( A1 => A(30), A2 => n1, B1 => B(30), B2 => n4, ZN =>
                           n98);
   U47 : INV_X1 port map( A => n87, ZN => Y(20));
   U48 : AOI22_X1 port map( A1 => A(20), A2 => n1, B1 => B(20), B2 => n6, ZN =>
                           n87);
   U49 : INV_X1 port map( A => n76, ZN => Y(10));
   U50 : AOI22_X1 port map( A1 => A(10), A2 => SEL, B1 => B(10), B2 => n9, ZN 
                           => n76);
   U51 : INV_X1 port map( A => n78, ZN => Y(12));
   U52 : AOI22_X1 port map( A1 => A(12), A2 => n1, B1 => B(12), B2 => n9, ZN =>
                           n78);
   U53 : INV_X1 port map( A => n81, ZN => Y(15));
   U54 : AOI22_X1 port map( A1 => A(15), A2 => SEL, B1 => B(15), B2 => n8, ZN 
                           => n81);
   U55 : INV_X1 port map( A => n84, ZN => Y(18));
   U56 : AOI22_X1 port map( A1 => A(18), A2 => n1, B1 => B(18), B2 => n7, ZN =>
                           n84);
   U57 : INV_X1 port map( A => n90, ZN => Y(23));
   U58 : AOI22_X1 port map( A1 => A(23), A2 => n1, B1 => B(23), B2 => n6, ZN =>
                           n90);
   U59 : INV_X1 port map( A => n93, ZN => Y(26));
   U60 : AOI22_X1 port map( A1 => A(26), A2 => n1, B1 => B(26), B2 => n5, ZN =>
                           n93);
   U61 : INV_X1 port map( A => n96, ZN => Y(29));
   U62 : AOI22_X1 port map( A1 => A(29), A2 => n1, B1 => B(29), B2 => n4, ZN =>
                           n96);
   U63 : INV_X1 port map( A => n100, ZN => Y(3));
   U64 : AOI22_X1 port map( A1 => A(3), A2 => n1, B1 => B(3), B2 => n3, ZN => 
                           n100);
   U65 : INV_X1 port map( A => n104, ZN => Y(7));
   U66 : AOI22_X1 port map( A1 => A(7), A2 => SEL, B1 => B(7), B2 => n2, ZN => 
                           n104);
   U67 : INV_X1 port map( A => n105, ZN => Y(8));
   U68 : AOI22_X1 port map( A1 => A(8), A2 => n1, B1 => B(8), B2 => n2, ZN => 
                           n105);
   U69 : INV_X1 port map( A => n99, ZN => Y(31));
   U70 : AOI22_X1 port map( A1 => A(31), A2 => SEL, B1 => B(31), B2 => n3, ZN 
                           => n99);
   U71 : INV_X1 port map( A => n75, ZN => Y(0));
   U72 : INV_X1 port map( A => n86, ZN => Y(1));
   U73 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n7, ZN => 
                           n86);
   U74 : AOI22_X1 port map( A1 => A(0), A2 => n1, B1 => B(0), B2 => n9, ZN => 
                           n75);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => n1, Z => Y(0));
   U5 : MUX2_X1 port map( A => B(1), B => A(1), S => n1, Z => Y(1));
   U6 : MUX2_X1 port map( A => B(2), B => A(2), S => n1, Z => Y(2));
   U7 : MUX2_X1 port map( A => B(3), B => A(3), S => n1, Z => Y(3));
   U8 : MUX2_X1 port map( A => B(4), B => A(4), S => n1, Z => Y(4));
   U9 : MUX2_X1 port map( A => B(5), B => A(5), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => B(6), B => A(6), S => n1, Z => Y(6));
   U11 : MUX2_X1 port map( A => B(7), B => A(7), S => n1, Z => Y(7));
   U12 : MUX2_X1 port map( A => B(8), B => A(8), S => n1, Z => Y(8));
   U13 : MUX2_X1 port map( A => B(9), B => A(9), S => n1, Z => Y(9));
   U14 : MUX2_X1 port map( A => B(10), B => A(10), S => n1, Z => Y(10));
   U15 : MUX2_X1 port map( A => B(11), B => A(11), S => n1, Z => Y(11));
   U16 : MUX2_X1 port map( A => B(12), B => A(12), S => n2, Z => Y(12));
   U17 : MUX2_X1 port map( A => B(13), B => A(13), S => n2, Z => Y(13));
   U18 : MUX2_X1 port map( A => B(14), B => A(14), S => n2, Z => Y(14));
   U19 : MUX2_X1 port map( A => B(15), B => A(15), S => n2, Z => Y(15));
   U20 : MUX2_X1 port map( A => B(16), B => A(16), S => n2, Z => Y(16));
   U21 : MUX2_X1 port map( A => B(17), B => A(17), S => n2, Z => Y(17));
   U22 : MUX2_X1 port map( A => B(18), B => A(18), S => n2, Z => Y(18));
   U23 : MUX2_X1 port map( A => B(19), B => A(19), S => n2, Z => Y(19));
   U24 : MUX2_X1 port map( A => B(20), B => A(20), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => B(21), B => A(21), S => n2, Z => Y(21));
   U26 : MUX2_X1 port map( A => B(22), B => A(22), S => n2, Z => Y(22));
   U27 : MUX2_X1 port map( A => B(23), B => A(23), S => n2, Z => Y(23));
   U28 : MUX2_X1 port map( A => B(24), B => A(24), S => n3, Z => Y(24));
   U29 : MUX2_X1 port map( A => B(25), B => A(25), S => n3, Z => Y(25));
   U30 : MUX2_X1 port map( A => B(26), B => A(26), S => n3, Z => Y(26));
   U31 : MUX2_X1 port map( A => B(27), B => A(27), S => n3, Z => Y(27));
   U32 : MUX2_X1 port map( A => B(28), B => A(28), S => n3, Z => Y(28));
   U33 : MUX2_X1 port map( A => B(29), B => A(29), S => n3, Z => Y(29));
   U34 : MUX2_X1 port map( A => B(30), B => A(30), S => n3, Z => Y(30));
   U35 : MUX2_X1 port map( A => B(31), B => A(31), S => n3, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : MUX2_X1 port map( A => B(4), B => A(4), S => n1, Z => Y(4));
   U3 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U5 : MUX2_X1 port map( A => B(0), B => A(0), S => n1, Z => Y(0));
   U6 : MUX2_X1 port map( A => B(1), B => A(1), S => n1, Z => Y(1));
   U7 : MUX2_X1 port map( A => B(2), B => A(2), S => n1, Z => Y(2));
   U8 : MUX2_X1 port map( A => B(3), B => A(3), S => n1, Z => Y(3));
   U9 : MUX2_X1 port map( A => B(5), B => A(5), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => B(6), B => A(6), S => n1, Z => Y(6));
   U11 : MUX2_X1 port map( A => B(7), B => A(7), S => n1, Z => Y(7));
   U12 : MUX2_X1 port map( A => B(8), B => A(8), S => n1, Z => Y(8));
   U13 : MUX2_X1 port map( A => B(9), B => A(9), S => n1, Z => Y(9));
   U14 : MUX2_X1 port map( A => B(10), B => A(10), S => n1, Z => Y(10));
   U15 : MUX2_X1 port map( A => B(11), B => A(11), S => n1, Z => Y(11));
   U16 : MUX2_X1 port map( A => B(12), B => A(12), S => n2, Z => Y(12));
   U17 : MUX2_X1 port map( A => B(13), B => A(13), S => n2, Z => Y(13));
   U18 : MUX2_X1 port map( A => B(14), B => A(14), S => n2, Z => Y(14));
   U19 : MUX2_X1 port map( A => B(15), B => A(15), S => n2, Z => Y(15));
   U20 : MUX2_X1 port map( A => B(16), B => A(16), S => n2, Z => Y(16));
   U21 : MUX2_X1 port map( A => B(17), B => A(17), S => n2, Z => Y(17));
   U22 : MUX2_X1 port map( A => B(18), B => A(18), S => n2, Z => Y(18));
   U23 : MUX2_X1 port map( A => B(19), B => A(19), S => n2, Z => Y(19));
   U24 : MUX2_X1 port map( A => B(20), B => A(20), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => B(21), B => A(21), S => n2, Z => Y(21));
   U26 : MUX2_X1 port map( A => B(22), B => A(22), S => n2, Z => Y(22));
   U27 : MUX2_X1 port map( A => B(23), B => A(23), S => n2, Z => Y(23));
   U28 : MUX2_X1 port map( A => B(24), B => A(24), S => n3, Z => Y(24));
   U29 : MUX2_X1 port map( A => B(25), B => A(25), S => n3, Z => Y(25));
   U30 : MUX2_X1 port map( A => B(26), B => A(26), S => n3, Z => Y(26));
   U31 : MUX2_X1 port map( A => B(27), B => A(27), S => n3, Z => Y(27));
   U32 : MUX2_X1 port map( A => B(28), B => A(28), S => n3, Z => Y(28));
   U33 : MUX2_X1 port map( A => B(29), B => A(29), S => n3, Z => Y(29));
   U34 : MUX2_X1 port map( A => B(30), B => A(30), S => n3, Z => Y(30));
   U35 : MUX2_X1 port map( A => B(31), B => A(31), S => n3, Z => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => Y(1));
   U2 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n8);
   U3 : INV_X1 port map( A => n7, ZN => Y(2));
   U4 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n7);
   U5 : INV_X1 port map( A => n6, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n6);
   U7 : INV_X1 port map( A => n9, ZN => Y(0));
   U8 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n9);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity carry_select_block_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_block_N4_0;

architecture SYN_STRUCTURAL of carry_select_block_N4_0 is

   component MUX21_GENERIC_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1136, n_1137 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S0_3_port, 
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1136);
   RCA1 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1137);
   MUXSUM : MUX21_GENERIC_N4_0 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity BUFF_0 is

   port( IG, IP : in std_logic;  OG, OP : out std_logic);

end BUFF_0;

architecture SYN_BEHAVIORAL of BUFF_0 is

begin
   OG <= IG;
   OP <= IP;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity PG_0 is

   port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);

end PG_0;

architecture SYN_BEHAVIORAL of PG_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PB, A2 => PA, ZN => P);
   U2 : INV_X1 port map( A => n2, ZN => G);
   U3 : AOI21_X1 port map( B1 => GB, B2 => PA, A => GA, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity and_gate_0 is

   port( A, B : in std_logic;  O : out std_logic);

end and_gate_0;

architecture SYN_behavioral of and_gate_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity xor_gate_0 is

   port( A, B : in std_logic;  O : out std_logic);

end xor_gate_0;

architecture SYN_behavioral of xor_gate_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => O);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity G_0 is

   port( PA, GA, GB : in std_logic;  G : out std_logic);

end G_0;

architecture SYN_BEHAVIORAL of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => G);
   U2 : AOI21_X1 port map( B1 => PA, B2 => GB, A => GA, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (7 downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component carry_select_block_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   BLI_0 : carry_select_block_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), Ci => Cin(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   BLI_1 : carry_select_block_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), Ci => Cin(1), S(3) => 
                           S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   BLI_2 : carry_select_block_N4_6 port map( A(3) => A(11), A(2) => A(10), A(1)
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   BLI_3 : carry_select_block_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1)
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   BLI_4 : carry_select_block_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1)
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   BLI_5 : carry_select_block_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1)
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   BLI_6 : carry_select_block_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1)
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   BLI_7 : carry_select_block_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1)
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_STRUCTURAL of 
   CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_1
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component G_2
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component G_3
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component G_4
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component PG_1
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_2
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component BUFF_1
      port( IG, IP : in std_logic;  OG, OP : out std_logic);
   end component;
   
   component BUFF_2
      port( IG, IP : in std_logic;  OG, OP : out std_logic);
   end component;
   
   component G_5
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component G_6
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component PG_3
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component BUFF_3
      port( IG, IP : in std_logic;  OG, OP : out std_logic);
   end component;
   
   component PG_4
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component BUFF_4
      port( IG, IP : in std_logic;  OG, OP : out std_logic);
   end component;
   
   component PG_5
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component BUFF_0
      port( IG, IP : in std_logic;  OG, OP : out std_logic);
   end component;
   
   component G_7
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component PG_6
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_7
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_8
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_9
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_10
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_11
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_12
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component G_8
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component PG_13
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_14
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_15
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_16
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_17
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_18
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_19
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_20
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_21
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_22
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_23
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_24
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_25
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_26
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_0
      port( PA, PB, GA, GB : in std_logic;  P, G : out std_logic);
   end component;
   
   component G_9
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   component and_gate_1
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_1
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_2
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_2
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_3
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_3
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_4
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_4
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_5
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_5
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_6
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_6
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_7
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_7
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_8
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_8
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_9
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_9
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_10
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_10
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_11
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_11
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_12
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_12
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_13
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_13
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_14
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_14
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_15
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_15
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_16
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_16
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_17
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_17
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_18
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_18
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_19
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_19
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_20
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_20
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_21
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_21
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_22
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_22
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_23
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_23
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_24
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_24
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_25
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_25
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_26
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_26
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_27
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_27
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_28
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_28
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_29
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_29
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_30
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_30
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_31
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_31
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component and_gate_0
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component xor_gate_0
      port( A, B : in std_logic;  O : out std_logic);
   end component;
   
   component G_0
      port( PA, GA, GB : in std_logic;  G : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, n8, Co_2_port, n9, n10, 
      Psubtractor, Gsubtractor, matrixG_4_31_port, matrixG_4_27_port, 
      matrixG_4_23_port, matrixG_4_19_port, matrixG_3_31_port, 
      matrixG_3_27_port, matrixG_3_23_port, matrixG_3_19_port, 
      matrixG_3_15_port, matrixG_3_11_port, matrixG_2_31_port, 
      matrixG_2_27_port, matrixG_2_23_port, matrixG_2_19_port, 
      matrixG_2_15_port, matrixG_2_11_port, matrixG_2_7_port, matrixG_1_31_port
      , matrixG_1_29_port, matrixG_1_27_port, matrixG_1_25_port, 
      matrixG_1_23_port, matrixG_1_21_port, matrixG_1_19_port, 
      matrixG_1_17_port, matrixG_1_15_port, matrixG_1_13_port, 
      matrixG_1_11_port, matrixG_1_9_port, matrixG_1_7_port, matrixG_1_5_port, 
      matrixG_1_3_port, matrixG_1_1_port, matrixG_0_31_port, matrixG_0_30_port,
      matrixG_0_29_port, matrixG_0_28_port, matrixG_0_27_port, 
      matrixG_0_26_port, matrixG_0_25_port, matrixG_0_24_port, 
      matrixG_0_23_port, matrixG_0_22_port, matrixG_0_21_port, 
      matrixG_0_20_port, matrixG_0_19_port, matrixG_0_18_port, 
      matrixG_0_17_port, matrixG_0_16_port, matrixG_0_15_port, 
      matrixG_0_14_port, matrixG_0_13_port, matrixG_0_12_port, 
      matrixG_0_11_port, matrixG_0_10_port, matrixG_0_9_port, matrixG_0_8_port,
      matrixG_0_7_port, matrixG_0_6_port, matrixG_0_5_port, matrixG_0_4_port, 
      matrixG_0_3_port, matrixG_0_2_port, matrixG_0_1_port, matrixG_0_0_port, 
      matrixP_4_31_port, matrixP_4_27_port, matrixP_4_23_port, 
      matrixP_4_19_port, matrixP_3_31_port, matrixP_3_27_port, 
      matrixP_3_23_port, matrixP_3_19_port, matrixP_3_15_port, 
      matrixP_3_11_port, matrixP_2_31_port, matrixP_2_27_port, 
      matrixP_2_23_port, matrixP_2_19_port, matrixP_2_15_port, 
      matrixP_2_11_port, matrixP_2_7_port, matrixP_1_31_port, matrixP_1_29_port
      , matrixP_1_27_port, matrixP_1_25_port, matrixP_1_23_port, 
      matrixP_1_21_port, matrixP_1_19_port, matrixP_1_17_port, 
      matrixP_1_15_port, matrixP_1_13_port, matrixP_1_11_port, matrixP_1_9_port
      , matrixP_1_7_port, matrixP_1_5_port, matrixP_1_3_port, matrixP_0_31_port
      , matrixP_0_30_port, matrixP_0_29_port, matrixP_0_28_port, 
      matrixP_0_27_port, matrixP_0_26_port, matrixP_0_25_port, 
      matrixP_0_24_port, matrixP_0_23_port, matrixP_0_22_port, 
      matrixP_0_21_port, matrixP_0_20_port, matrixP_0_19_port, 
      matrixP_0_18_port, matrixP_0_17_port, matrixP_0_16_port, 
      matrixP_0_15_port, matrixP_0_14_port, matrixP_0_13_port, 
      matrixP_0_12_port, matrixP_0_11_port, matrixP_0_10_port, matrixP_0_9_port
      , matrixP_0_8_port, matrixP_0_7_port, matrixP_0_6_port, matrixP_0_5_port,
      matrixP_0_4_port, matrixP_0_3_port, matrixP_0_2_port, matrixP_0_1_port, 
      n1, n2, Co_0_port, Co_1_port, n5, Co_3_port, n7 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   Gsub : G_0 port map( PA => Psubtractor, GA => Gsubtractor, GB => Cin, G => 
                           matrixG_0_0_port);
   Xor_gsi_0_0 : xor_gate_0 port map( A => A(0), B => B(0), O => Psubtractor);
   and_gsi_0_0 : and_gate_0 port map( A => A(0), B => B(0), O => Gsubtractor);
   Xor_gsi_0_1 : xor_gate_31 port map( A => A(1), B => B(1), O => 
                           matrixP_0_1_port);
   and_gsi_0_1 : and_gate_31 port map( A => A(1), B => B(1), O => 
                           matrixG_0_1_port);
   Xor_gsi_0_2 : xor_gate_30 port map( A => A(2), B => B(2), O => 
                           matrixP_0_2_port);
   and_gsi_0_2 : and_gate_30 port map( A => A(2), B => B(2), O => 
                           matrixG_0_2_port);
   Xor_gsi_0_3 : xor_gate_29 port map( A => A(3), B => B(3), O => 
                           matrixP_0_3_port);
   and_gsi_0_3 : and_gate_29 port map( A => A(3), B => B(3), O => 
                           matrixG_0_3_port);
   Xor_gsi_0_4 : xor_gate_28 port map( A => A(4), B => B(4), O => 
                           matrixP_0_4_port);
   and_gsi_0_4 : and_gate_28 port map( A => A(4), B => B(4), O => 
                           matrixG_0_4_port);
   Xor_gsi_0_5 : xor_gate_27 port map( A => A(5), B => B(5), O => 
                           matrixP_0_5_port);
   and_gsi_0_5 : and_gate_27 port map( A => A(5), B => B(5), O => 
                           matrixG_0_5_port);
   Xor_gsi_0_6 : xor_gate_26 port map( A => A(6), B => B(6), O => 
                           matrixP_0_6_port);
   and_gsi_0_6 : and_gate_26 port map( A => A(6), B => B(6), O => 
                           matrixG_0_6_port);
   Xor_gsi_0_7 : xor_gate_25 port map( A => A(7), B => B(7), O => 
                           matrixP_0_7_port);
   and_gsi_0_7 : and_gate_25 port map( A => A(7), B => n1, O => 
                           matrixG_0_7_port);
   Xor_gsi_0_8 : xor_gate_24 port map( A => A(8), B => B(8), O => 
                           matrixP_0_8_port);
   and_gsi_0_8 : and_gate_24 port map( A => A(8), B => B(8), O => 
                           matrixG_0_8_port);
   Xor_gsi_0_9 : xor_gate_23 port map( A => A(9), B => B(9), O => 
                           matrixP_0_9_port);
   and_gsi_0_9 : and_gate_23 port map( A => A(9), B => B(9), O => 
                           matrixG_0_9_port);
   Xor_gsi_0_10 : xor_gate_22 port map( A => A(10), B => B(10), O => 
                           matrixP_0_10_port);
   and_gsi_0_10 : and_gate_22 port map( A => A(10), B => B(10), O => 
                           matrixG_0_10_port);
   Xor_gsi_0_11 : xor_gate_21 port map( A => A(11), B => B(11), O => 
                           matrixP_0_11_port);
   and_gsi_0_11 : and_gate_21 port map( A => A(11), B => B(11), O => 
                           matrixG_0_11_port);
   Xor_gsi_0_12 : xor_gate_20 port map( A => A(12), B => B(12), O => 
                           matrixP_0_12_port);
   and_gsi_0_12 : and_gate_20 port map( A => A(12), B => B(12), O => 
                           matrixG_0_12_port);
   Xor_gsi_0_13 : xor_gate_19 port map( A => A(13), B => B(13), O => 
                           matrixP_0_13_port);
   and_gsi_0_13 : and_gate_19 port map( A => A(13), B => B(13), O => 
                           matrixG_0_13_port);
   Xor_gsi_0_14 : xor_gate_18 port map( A => A(14), B => B(14), O => 
                           matrixP_0_14_port);
   and_gsi_0_14 : and_gate_18 port map( A => A(14), B => B(14), O => 
                           matrixG_0_14_port);
   Xor_gsi_0_15 : xor_gate_17 port map( A => A(15), B => B(15), O => 
                           matrixP_0_15_port);
   and_gsi_0_15 : and_gate_17 port map( A => A(15), B => B(15), O => 
                           matrixG_0_15_port);
   Xor_gsi_0_16 : xor_gate_16 port map( A => A(16), B => B(16), O => 
                           matrixP_0_16_port);
   and_gsi_0_16 : and_gate_16 port map( A => A(16), B => B(16), O => 
                           matrixG_0_16_port);
   Xor_gsi_0_17 : xor_gate_15 port map( A => A(17), B => B(17), O => 
                           matrixP_0_17_port);
   and_gsi_0_17 : and_gate_15 port map( A => A(17), B => B(17), O => 
                           matrixG_0_17_port);
   Xor_gsi_0_18 : xor_gate_14 port map( A => A(18), B => B(18), O => 
                           matrixP_0_18_port);
   and_gsi_0_18 : and_gate_14 port map( A => A(18), B => B(18), O => 
                           matrixG_0_18_port);
   Xor_gsi_0_19 : xor_gate_13 port map( A => A(19), B => B(19), O => 
                           matrixP_0_19_port);
   and_gsi_0_19 : and_gate_13 port map( A => A(19), B => B(19), O => 
                           matrixG_0_19_port);
   Xor_gsi_0_20 : xor_gate_12 port map( A => A(20), B => B(20), O => 
                           matrixP_0_20_port);
   and_gsi_0_20 : and_gate_12 port map( A => A(20), B => B(20), O => 
                           matrixG_0_20_port);
   Xor_gsi_0_21 : xor_gate_11 port map( A => A(21), B => B(21), O => 
                           matrixP_0_21_port);
   and_gsi_0_21 : and_gate_11 port map( A => A(21), B => B(21), O => 
                           matrixG_0_21_port);
   Xor_gsi_0_22 : xor_gate_10 port map( A => A(22), B => B(22), O => 
                           matrixP_0_22_port);
   and_gsi_0_22 : and_gate_10 port map( A => A(22), B => B(22), O => 
                           matrixG_0_22_port);
   Xor_gsi_0_23 : xor_gate_9 port map( A => A(23), B => B(23), O => 
                           matrixP_0_23_port);
   and_gsi_0_23 : and_gate_9 port map( A => A(23), B => B(23), O => 
                           matrixG_0_23_port);
   Xor_gsi_0_24 : xor_gate_8 port map( A => A(24), B => B(24), O => 
                           matrixP_0_24_port);
   and_gsi_0_24 : and_gate_8 port map( A => A(24), B => B(24), O => 
                           matrixG_0_24_port);
   Xor_gsi_0_25 : xor_gate_7 port map( A => A(25), B => B(25), O => 
                           matrixP_0_25_port);
   and_gsi_0_25 : and_gate_7 port map( A => A(25), B => B(25), O => 
                           matrixG_0_25_port);
   Xor_gsi_0_26 : xor_gate_6 port map( A => A(26), B => B(26), O => 
                           matrixP_0_26_port);
   and_gsi_0_26 : and_gate_6 port map( A => A(26), B => B(26), O => 
                           matrixG_0_26_port);
   Xor_gsi_0_27 : xor_gate_5 port map( A => A(27), B => B(27), O => 
                           matrixP_0_27_port);
   and_gsi_0_27 : and_gate_5 port map( A => A(27), B => B(27), O => 
                           matrixG_0_27_port);
   Xor_gsi_0_28 : xor_gate_4 port map( A => A(28), B => B(28), O => 
                           matrixP_0_28_port);
   and_gsi_0_28 : and_gate_4 port map( A => A(28), B => B(28), O => 
                           matrixG_0_28_port);
   Xor_gsi_0_29 : xor_gate_3 port map( A => A(29), B => B(29), O => 
                           matrixP_0_29_port);
   and_gsi_0_29 : and_gate_3 port map( A => A(29), B => B(29), O => 
                           matrixG_0_29_port);
   Xor_gsi_0_30 : xor_gate_2 port map( A => A(30), B => B(30), O => 
                           matrixP_0_30_port);
   and_gsi_0_30 : and_gate_2 port map( A => A(30), B => B(30), O => 
                           matrixG_0_30_port);
   Xor_gsi_0_31 : xor_gate_1 port map( A => A(31), B => B(31), O => 
                           matrixP_0_31_port);
   and_gsi_0_31 : and_gate_1 port map( A => A(31), B => B(31), O => 
                           matrixG_0_31_port);
   Gs_d_1_1 : G_9 port map( PA => matrixP_0_1_port, GA => matrixG_0_1_port, GB 
                           => matrixG_0_0_port, G => matrixG_1_1_port);
   PGsi_1_3 : PG_0 port map( PA => matrixP_0_3_port, PB => matrixP_0_2_port, GA
                           => matrixG_0_3_port, GB => matrixG_0_2_port, P => 
                           matrixP_1_3_port, G => matrixG_1_3_port);
   PGsi_1_5 : PG_26 port map( PA => matrixP_0_5_port, PB => matrixP_0_4_port, 
                           GA => matrixG_0_5_port, GB => matrixG_0_4_port, P =>
                           matrixP_1_5_port, G => matrixG_1_5_port);
   PGsi_1_7 : PG_25 port map( PA => matrixP_0_7_port, PB => matrixP_0_6_port, 
                           GA => matrixG_0_7_port, GB => matrixG_0_6_port, P =>
                           matrixP_1_7_port, G => matrixG_1_7_port);
   PGsi_1_9 : PG_24 port map( PA => matrixP_0_9_port, PB => matrixP_0_8_port, 
                           GA => matrixG_0_9_port, GB => matrixG_0_8_port, P =>
                           matrixP_1_9_port, G => matrixG_1_9_port);
   PGsi_1_11 : PG_23 port map( PA => matrixP_0_11_port, PB => matrixP_0_10_port
                           , GA => matrixG_0_11_port, GB => matrixG_0_10_port, 
                           P => matrixP_1_11_port, G => matrixG_1_11_port);
   PGsi_1_13 : PG_22 port map( PA => matrixP_0_13_port, PB => matrixP_0_12_port
                           , GA => matrixG_0_13_port, GB => matrixG_0_12_port, 
                           P => matrixP_1_13_port, G => matrixG_1_13_port);
   PGsi_1_15 : PG_21 port map( PA => matrixP_0_15_port, PB => matrixP_0_14_port
                           , GA => matrixG_0_15_port, GB => matrixG_0_14_port, 
                           P => matrixP_1_15_port, G => matrixG_1_15_port);
   PGsi_1_17 : PG_20 port map( PA => matrixP_0_17_port, PB => matrixP_0_16_port
                           , GA => matrixG_0_17_port, GB => matrixG_0_16_port, 
                           P => matrixP_1_17_port, G => matrixG_1_17_port);
   PGsi_1_19 : PG_19 port map( PA => matrixP_0_19_port, PB => matrixP_0_18_port
                           , GA => matrixG_0_19_port, GB => matrixG_0_18_port, 
                           P => matrixP_1_19_port, G => matrixG_1_19_port);
   PGsi_1_21 : PG_18 port map( PA => matrixP_0_21_port, PB => matrixP_0_20_port
                           , GA => matrixG_0_21_port, GB => matrixG_0_20_port, 
                           P => matrixP_1_21_port, G => matrixG_1_21_port);
   PGsi_1_23 : PG_17 port map( PA => matrixP_0_23_port, PB => matrixP_0_22_port
                           , GA => matrixG_0_23_port, GB => matrixG_0_22_port, 
                           P => matrixP_1_23_port, G => matrixG_1_23_port);
   PGsi_1_25 : PG_16 port map( PA => matrixP_0_25_port, PB => matrixP_0_24_port
                           , GA => matrixG_0_25_port, GB => matrixG_0_24_port, 
                           P => matrixP_1_25_port, G => matrixG_1_25_port);
   PGsi_1_27 : PG_15 port map( PA => matrixP_0_27_port, PB => matrixP_0_26_port
                           , GA => matrixG_0_27_port, GB => matrixG_0_26_port, 
                           P => matrixP_1_27_port, G => matrixG_1_27_port);
   PGsi_1_29 : PG_14 port map( PA => matrixP_0_29_port, PB => matrixP_0_28_port
                           , GA => matrixG_0_29_port, GB => matrixG_0_28_port, 
                           P => matrixP_1_29_port, G => matrixG_1_29_port);
   PGsi_1_31 : PG_13 port map( PA => matrixP_0_31_port, PB => matrixP_0_30_port
                           , GA => matrixG_0_31_port, GB => matrixG_0_30_port, 
                           P => matrixP_1_31_port, G => matrixG_1_31_port);
   Gs_d_2_3 : G_8 port map( PA => matrixP_1_3_port, GA => matrixG_1_3_port, GB 
                           => matrixG_1_1_port, G => n10);
   PGsi_2_7 : PG_12 port map( PA => matrixP_1_7_port, PB => matrixP_1_5_port, 
                           GA => matrixG_1_7_port, GB => matrixG_1_5_port, P =>
                           matrixP_2_7_port, G => matrixG_2_7_port);
   PGsi_2_11 : PG_11 port map( PA => matrixP_1_11_port, PB => matrixP_1_9_port,
                           GA => matrixG_1_11_port, GB => matrixG_1_9_port, P 
                           => matrixP_2_11_port, G => matrixG_2_11_port);
   PGsi_2_15 : PG_10 port map( PA => matrixP_1_15_port, PB => matrixP_1_13_port
                           , GA => matrixG_1_15_port, GB => matrixG_1_13_port, 
                           P => matrixP_2_15_port, G => matrixG_2_15_port);
   PGsi_2_19 : PG_9 port map( PA => matrixP_1_19_port, PB => matrixP_1_17_port,
                           GA => matrixG_1_19_port, GB => matrixG_1_17_port, P 
                           => matrixP_2_19_port, G => matrixG_2_19_port);
   PGsi_2_23 : PG_8 port map( PA => matrixP_1_23_port, PB => matrixP_1_21_port,
                           GA => matrixG_1_23_port, GB => matrixG_1_21_port, P 
                           => matrixP_2_23_port, G => matrixG_2_23_port);
   PGsi_2_27 : PG_7 port map( PA => matrixP_1_27_port, PB => matrixP_1_25_port,
                           GA => matrixG_1_27_port, GB => matrixG_1_25_port, P 
                           => matrixP_2_27_port, G => matrixG_2_27_port);
   PGsi_2_31 : PG_6 port map( PA => matrixP_1_31_port, PB => matrixP_1_29_port,
                           GA => matrixG_1_31_port, GB => matrixG_1_29_port, P 
                           => matrixP_2_31_port, G => matrixG_2_31_port);
   Gs_h_3_7 : G_7 port map( PA => matrixP_2_7_port, GA => matrixG_2_7_port, GB 
                           => n10, G => n9);
   Buf_h_3_11 : BUFF_0 port map( IG => matrixG_2_11_port, IP => 
                           matrixP_2_11_port, OG => matrixG_3_11_port, OP => 
                           matrixP_3_11_port);
   PGsi_3_15 : PG_5 port map( PA => matrixP_2_15_port, PB => matrixP_3_11_port,
                           GA => matrixG_2_15_port, GB => matrixG_2_11_port, P 
                           => matrixP_3_15_port, G => matrixG_3_15_port);
   Buf_h_3_19 : BUFF_4 port map( IG => n2, IP => matrixP_2_19_port, OG => 
                           matrixG_3_19_port, OP => matrixP_3_19_port);
   PGsi_3_23 : PG_4 port map( PA => matrixP_2_23_port, PB => matrixP_3_19_port,
                           GA => matrixG_2_23_port, GB => matrixG_2_19_port, P 
                           => matrixP_3_23_port, G => matrixG_3_23_port);
   Buf_h_3_27 : BUFF_3 port map( IG => matrixG_2_27_port, IP => 
                           matrixP_2_27_port, OG => matrixG_3_27_port, OP => 
                           matrixP_3_27_port);
   PGsi_3_31 : PG_3 port map( PA => matrixP_2_31_port, PB => matrixP_3_27_port,
                           GA => matrixG_2_31_port, GB => matrixG_2_27_port, P 
                           => matrixP_3_31_port, G => matrixG_3_31_port);
   Gs_h_4_11 : G_6 port map( PA => matrixP_3_11_port, GA => matrixG_3_11_port, 
                           GB => Co_1_port, G => Co_2_port);
   Gs_h_4_15 : G_5 port map( PA => matrixP_3_15_port, GA => matrixG_3_15_port, 
                           GB => n9, G => n8);
   Buf_h_4_19_0 : BUFF_2 port map( IG => matrixG_3_19_port, IP => 
                           matrixP_3_19_port, OG => matrixG_4_19_port, OP => 
                           matrixP_4_19_port);
   Buf_h_4_23_0 : BUFF_1 port map( IG => n7, IP => matrixP_3_23_port, OG => 
                           matrixG_4_23_port, OP => matrixP_4_23_port);
   PGsi_4_27_0 : PG_2 port map( PA => matrixP_3_27_port, PB => 
                           matrixP_3_23_port, GA => matrixG_3_27_port, GB => 
                           matrixG_3_23_port, P => matrixP_4_27_port, G => 
                           matrixG_4_27_port);
   PGsi_4_31_0 : PG_1 port map( PA => matrixP_3_31_port, PB => 
                           matrixP_3_23_port, GA => matrixG_3_31_port, GB => n7
                           , P => matrixP_4_31_port, G => matrixG_4_31_port);
   Gs_h_5_19 : G_4 port map( PA => matrixP_4_19_port, GA => matrixG_4_19_port, 
                           GB => n8, G => Co_4_port);
   Gs_h_5_23 : G_3 port map( PA => matrixP_4_23_port, GA => matrixG_4_23_port, 
                           GB => n8, G => Co_5_port);
   Gs_h_5_27 : G_2 port map( PA => matrixP_4_27_port, GA => matrixG_4_27_port, 
                           GB => n8, G => Co_6_port);
   Gs_h_5_31 : G_1 port map( PA => matrixP_4_31_port, GA => matrixG_4_31_port, 
                           GB => Co_3_port, G => Co_7_port);
   U1 : INV_X2 port map( A => n5, ZN => Co_3_port);
   U2 : CLKBUF_X1 port map( A => B(7), Z => n1);
   U3 : CLKBUF_X1 port map( A => matrixG_2_19_port, Z => n2);
   U4 : BUF_X1 port map( A => matrixG_3_23_port, Z => n7);
   U5 : CLKBUF_X1 port map( A => n9, Z => Co_1_port);
   U6 : CLKBUF_X1 port map( A => n10, Z => Co_0_port);
   U7 : INV_X1 port map( A => n8, ZN => n5);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity P4_ADDER_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4_ADDER_NBIT32;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (7 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal carryv_6_port, carryv_5_port, carryv_4_port, carryv_3_port, 
      carryv_2_port, carryv_1_port, carryv_0_port, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21 : 
      std_logic;

begin
   
   C_GEN : CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4 port map( A(31) =>
                           A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B(31), B(30) => B(30), B(29) => n1, B(28) 
                           => n5, B(27) => B(27), B(26) => B(26), B(25) => 
                           B(25), B(24) => B(24), B(23) => B(23), B(22) => 
                           B(22), B(21) => B(21), B(20) => B(20), B(19) => 
                           B(19), B(18) => B(18), B(17) => B(17), B(16) => 
                           B(16), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, Co(7) => Cout, Co(6) => carryv_6_port, Co(5)
                           => carryv_5_port, Co(4) => carryv_4_port, Co(3) => 
                           carryv_3_port, Co(2) => carryv_2_port, Co(1) => 
                           carryv_1_port, Co(0) => carryv_0_port);
   S_GEN : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => n12, B(26) => n21, B(25) => n18, B(24) => 
                           B(24), B(23) => n19, B(22) => n17, B(21) => n11, 
                           B(20) => n14, B(19) => n20, B(18) => n9, B(17) => 
                           n13, B(16) => B(16), B(15) => n16, B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => n6, B(10) 
                           => B(10), B(9) => n8, B(8) => B(8), B(7) => n15, 
                           B(6) => n4, B(5) => n2, B(4) => B(4), B(3) => n3, 
                           B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin(7) => 
                           carryv_6_port, Cin(6) => carryv_5_port, Cin(5) => 
                           carryv_4_port, Cin(4) => carryv_3_port, Cin(3) => 
                           carryv_2_port, Cin(2) => carryv_1_port, Cin(1) => 
                           carryv_0_port, Cin(0) => Cin, S(31) => S(31), S(30) 
                           => S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));
   U1 : BUF_X1 port map( A => B(20), Z => n14);
   U2 : CLKBUF_X1 port map( A => B(29), Z => n1);
   U3 : CLKBUF_X1 port map( A => B(5), Z => n2);
   U4 : CLKBUF_X1 port map( A => B(3), Z => n3);
   U5 : CLKBUF_X1 port map( A => B(6), Z => n4);
   U6 : CLKBUF_X1 port map( A => B(28), Z => n5);
   U7 : CLKBUF_X1 port map( A => B(25), Z => n18);
   U8 : CLKBUF_X1 port map( A => B(11), Z => n6);
   U9 : INV_X1 port map( A => B(9), ZN => n7);
   U10 : INV_X1 port map( A => n7, ZN => n8);
   U11 : CLKBUF_X1 port map( A => B(18), Z => n9);
   U12 : INV_X1 port map( A => B(21), ZN => n10);
   U13 : INV_X1 port map( A => n10, ZN => n11);
   U14 : CLKBUF_X1 port map( A => B(27), Z => n12);
   U15 : CLKBUF_X1 port map( A => B(17), Z => n13);
   U16 : CLKBUF_X1 port map( A => B(7), Z => n15);
   U17 : CLKBUF_X1 port map( A => B(15), Z => n16);
   U18 : CLKBUF_X1 port map( A => B(22), Z => n17);
   U19 : CLKBUF_X1 port map( A => B(23), Z => n19);
   U20 : CLKBUF_X1 port map( A => B(19), Z => n20);
   U21 : CLKBUF_X1 port map( A => B(26), Z => n21);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity add_sub_N32 is

   port( A : in std_logic_vector (31 downto 0);  SEL : in std_logic_vector (0 
         to 4);  O : out std_logic_vector (31 downto 0));

end add_sub_N32;

architecture SYN_Behavioral of add_sub_N32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component add_sub_N32_DW01_sub_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n3_port, n4_port, net29489, net29487, net29485, net37049, 
      net37424, net37956, net39102, net37839, net37838, n1, n2_port, n5_port, 
      n6_port, n7_port, n8_port, n9_port, n10_port, n11_port, n12_port, 
      n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, n19_port, 
      n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n_1138 : std_logic;

begin
   
   n3_port <= '0';
   n4_port <= '0';
   sub_20 : add_sub_N32_DW01_sub_2 port map( A(31) => n3_port, A(30) => n3_port
                           , A(29) => n3_port, A(28) => n3_port, A(27) => 
                           n3_port, A(26) => n3_port, A(25) => n3_port, A(24) 
                           => n3_port, A(23) => n3_port, A(22) => n3_port, 
                           A(21) => n3_port, A(20) => n3_port, A(19) => n3_port
                           , A(18) => n3_port, A(17) => n3_port, A(16) => 
                           n3_port, A(15) => n3_port, A(14) => n3_port, A(13) 
                           => n3_port, A(12) => n3_port, A(11) => n3_port, 
                           A(10) => n3_port, A(9) => n3_port, A(8) => n3_port, 
                           A(7) => n3_port, A(6) => n3_port, A(5) => n3_port, 
                           A(4) => n3_port, A(3) => n3_port, A(2) => n3_port, 
                           A(1) => n3_port, A(0) => n3_port, B(31) => A(31), 
                           B(30) => A(30), B(29) => A(29), B(28) => A(28), 
                           B(27) => A(27), B(26) => A(26), B(25) => A(25), 
                           B(24) => A(24), B(23) => A(23), B(22) => A(22), 
                           B(21) => A(21), B(20) => A(20), B(19) => A(19), 
                           B(18) => A(18), B(17) => A(17), B(16) => A(16), 
                           B(15) => A(15), B(14) => A(14), B(13) => A(13), 
                           B(12) => A(12), B(11) => A(11), B(10) => A(10), B(9)
                           => A(9), B(8) => A(8), B(7) => A(7), B(6) => A(6), 
                           B(5) => A(5), B(4) => A(4), B(3) => A(3), B(2) => 
                           A(2), B(1) => A(1), B(0) => A(0), CI => n4_port, 
                           DIFF(31) => N33, DIFF(30) => N32, DIFF(29) => N31, 
                           DIFF(28) => N30, DIFF(27) => N29, DIFF(26) => N28, 
                           DIFF(25) => N27, DIFF(24) => N26, DIFF(23) => N25, 
                           DIFF(22) => N24, DIFF(21) => N23, DIFF(20) => N22, 
                           DIFF(19) => N21, DIFF(18) => N20, DIFF(17) => N19, 
                           DIFF(16) => N18, DIFF(15) => N17, DIFF(14) => N16, 
                           DIFF(13) => N15, DIFF(12) => N14, DIFF(11) => N13, 
                           DIFF(10) => N12, DIFF(9) => N11, DIFF(8) => N10, 
                           DIFF(7) => N9, DIFF(6) => N8, DIFF(5) => N7, DIFF(4)
                           => N6, DIFF(3) => N5, DIFF(2) => N4, DIFF(1) => N3, 
                           DIFF(0) => N2, CO => n_1138);
   U4 : NAND2_X1 port map( A1 => N17, A2 => n1, ZN => n2_port);
   U5 : NAND2_X2 port map( A1 => n25_port, A2 => net37838, ZN => n5_port);
   U6 : NAND2_X1 port map( A1 => n2_port, A2 => n5_port, ZN => O(15));
   U7 : INV_X1 port map( A => net37838, ZN => n1);
   U8 : INV_X2 port map( A => net29487, ZN => net37838);
   U9 : NOR4_X1 port map( A1 => SEL(2), A2 => n13_port, A3 => SEL(0), A4 => 
                           SEL(1), ZN => n15_port);
   U10 : NAND2_X1 port map( A1 => A(17), A2 => net37956, ZN => n21_port);
   U11 : MUX2_X1 port map( A => A(13), B => N15, S => net29487, Z => O(13));
   U12 : MUX2_X1 port map( A => A(24), B => N26, S => net29489, Z => O(24));
   U13 : NAND2_X1 port map( A1 => A(19), A2 => net37838, ZN => net37839);
   U14 : CLKBUF_X1 port map( A => A(5), Z => n6_port);
   U15 : CLKBUF_X1 port map( A => A(10), Z => n7_port);
   U16 : CLKBUF_X1 port map( A => A(14), Z => n8_port);
   U17 : CLKBUF_X1 port map( A => A(0), Z => n9_port);
   U18 : INV_X1 port map( A => net29489, ZN => net37049);
   U19 : BUF_X1 port map( A => n15_port, Z => net29485);
   U20 : BUF_X1 port map( A => n15_port, Z => net29487);
   U21 : INV_X1 port map( A => net29489, ZN => net37424);
   U22 : NAND2_X1 port map( A1 => n28_port, A2 => n10_port, ZN => n11_port);
   U23 : NAND2_X1 port map( A1 => N8, A2 => net29485, ZN => n12_port);
   U24 : NAND2_X1 port map( A1 => n11_port, A2 => n12_port, ZN => O(6));
   U25 : INV_X1 port map( A => net29485, ZN => n10_port);
   U26 : MUX2_X2 port map( A => A(9), B => N11, S => net29485, Z => O(9));
   U27 : NAND2_X1 port map( A1 => N21, A2 => net29487, ZN => n16_port);
   U28 : NAND2_X1 port map( A1 => n16_port, A2 => net37839, ZN => O(19));
   U29 : CLKBUF_X1 port map( A => n15_port, Z => net29489);
   U30 : NAND2_X1 port map( A1 => SEL(3), A2 => n14_port, ZN => n13_port);
   U31 : INV_X1 port map( A => SEL(4), ZN => n14_port);
   U32 : NAND2_X1 port map( A1 => N20, A2 => net29489, ZN => n17_port);
   U33 : NAND2_X1 port map( A1 => A(18), A2 => net37424, ZN => n18_port);
   U34 : NAND2_X1 port map( A1 => n17_port, A2 => n18_port, ZN => O(18));
   U35 : NAND2_X1 port map( A1 => A(7), A2 => net39102, ZN => n19_port);
   U36 : NAND2_X1 port map( A1 => N9, A2 => net29485, ZN => n20_port);
   U37 : NAND2_X1 port map( A1 => n20_port, A2 => n19_port, ZN => O(7));
   U38 : INV_X1 port map( A => net29485, ZN => net39102);
   U39 : MUX2_X2 port map( A => A(8), B => N10, S => net29485, Z => O(8));
   U40 : MUX2_X1 port map( A => A(3), B => N5, S => net29485, Z => O(3));
   U41 : MUX2_X1 port map( A => A(25), B => N27, S => net29489, Z => O(25));
   U42 : NAND2_X1 port map( A1 => N19, A2 => net29487, ZN => n22_port);
   U43 : NAND2_X1 port map( A1 => n21_port, A2 => n22_port, ZN => O(17));
   U44 : INV_X1 port map( A => net29487, ZN => net37956);
   U45 : MUX2_X2 port map( A => A(22), B => N24, S => net29487, Z => O(22));
   U46 : NAND2_X1 port map( A1 => N29, A2 => net29489, ZN => n23_port);
   U47 : NAND2_X1 port map( A1 => A(27), A2 => net37049, ZN => n24_port);
   U48 : NAND2_X1 port map( A1 => n23_port, A2 => n24_port, ZN => O(27));
   U49 : MUX2_X2 port map( A => A(23), B => N25, S => net29487, Z => O(23));
   U50 : MUX2_X2 port map( A => n6_port, B => N7, S => net29485, Z => O(5));
   U51 : CLKBUF_X1 port map( A => A(15), Z => n25_port);
   U52 : MUX2_X2 port map( A => N22, B => A(20), S => net37956, Z => O(20));
   U53 : MUX2_X1 port map( A => A(21), B => N23, S => net29487, Z => O(21));
   U54 : NAND2_X1 port map( A1 => A(11), A2 => net37838, ZN => n26_port);
   U55 : NAND2_X1 port map( A1 => N13, A2 => net29485, ZN => n27_port);
   U56 : NAND2_X1 port map( A1 => n27_port, A2 => n26_port, ZN => O(11));
   U57 : MUX2_X2 port map( A => A(29), B => N31, S => net29489, Z => O(29));
   U58 : CLKBUF_X1 port map( A => A(6), Z => n28_port);
   U59 : NAND2_X1 port map( A1 => A(26), A2 => net37424, ZN => n29_port);
   U60 : NAND2_X1 port map( A1 => N28, A2 => net29489, ZN => n30_port);
   U61 : NAND2_X1 port map( A1 => n30_port, A2 => n29_port, ZN => O(26));
   U62 : MUX2_X2 port map( A => A(28), B => N30, S => net29489, Z => O(28));
   U63 : MUX2_X2 port map( A => n8_port, B => N16, S => net29487, Z => O(14));
   U64 : MUX2_X1 port map( A => n9_port, B => N2, S => net29485, Z => O(0));
   U65 : MUX2_X1 port map( A => A(1), B => N3, S => net29485, Z => O(1));
   U66 : MUX2_X1 port map( A => A(2), B => N4, S => net29485, Z => O(2));
   U67 : MUX2_X1 port map( A => A(4), B => N6, S => net29485, Z => O(4));
   U68 : MUX2_X1 port map( A => n7_port, B => N12, S => net29485, Z => O(10));
   U69 : MUX2_X1 port map( A => A(12), B => N14, S => net29487, Z => O(12));
   U70 : MUX2_X1 port map( A => A(16), B => N18, S => net29487, Z => O(16));
   U71 : MUX2_X1 port map( A => A(30), B => N32, S => net29489, Z => O(30));
   U72 : MUX2_X1 port map( A => A(31), B => N33, S => net29489, Z => O(31));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity mux4to1_N32 is

   port( inadd, inlog, insh, incom : in std_logic_vector (31 downto 0);  sel : 
         in std_logic_vector (0 to 4);  O : out std_logic_vector (31 downto 0)
         );

end mux4to1_N32;

architecture SYN_Behavioral of mux4to1_N32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n28, n29, n50, n51, n68, n69, n70, n71, net27574, net27576, net27607, 
      net29471, net29469, net29475, net29479, net29483, net29481, net38998, 
      net38995, net39329, net39295, net27572, net39337, net39325, net39320, 
      net39318, net39313, net39291, net39286, net39326, net39290, net27618, 
      net27616, net27611, net25507, n8, n1, n2, n3, n4, n5, n9, n10, n11, n24, 
      n25, n26, n27, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n72, n73, n74, n75, n76
      , n77 : std_logic;

begin
   
   U2 : NOR2_X1 port map( A1 => net39313, A2 => sel(2), ZN => net39320);
   U3 : INV_X1 port map( A => sel(1), ZN => net39313);
   U4 : INV_X1 port map( A => sel(0), ZN => n11);
   U5 : AOI21_X1 port map( B1 => net39326, B2 => net25507, A => sel(0), ZN => 
                           net39325);
   U6 : AOI21_X1 port map( B1 => n33, B2 => net39318, A => sel(2), ZN => n32);
   U7 : INV_X1 port map( A => sel(3), ZN => net39318);
   U8 : NOR2_X1 port map( A1 => sel(4), A2 => sel(0), ZN => n33);
   U9 : NAND2_X1 port map( A1 => sel(3), A2 => sel(4), ZN => net39326);
   U10 : NAND2_X1 port map( A1 => sel(1), A2 => net27611, ZN => net39290);
   U11 : OAI21_X1 port map( B1 => sel(3), B2 => sel(2), A => sel(0), ZN => n24)
                           ;
   U12 : NAND2_X1 port map( A1 => inlog(27), A2 => net29479, ZN => net38998);
   U13 : NAND2_X1 port map( A1 => net39286, A2 => n27, ZN => n26);
   U14 : NAND2_X1 port map( A1 => net39337, A2 => sel(3), ZN => n27);
   U15 : OAI21_X1 port map( B1 => net39320, B2 => net27611, A => n11, ZN => 
                           net39337);
   U16 : INV_X1 port map( A => inlog(28), ZN => net39329);
   U17 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => net39291);
   U18 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n30);
   U19 : NOR2_X1 port map( A1 => net27611, A2 => sel(2), ZN => n34);
   U20 : INV_X1 port map( A => sel(2), ZN => net25507);
   U21 : AND4_X1 port map( A1 => n11, A2 => sel(2), A3 => sel(3), A4 => 
                           net39290, ZN => n1);
   U22 : OR2_X1 port map( A1 => n37, A2 => net38995, ZN => n2);
   U23 : AND2_X1 port map( A1 => net39326, A2 => n11, ZN => n3);
   U24 : OR2_X1 port map( A1 => net39291, A2 => net39329, ZN => n4);
   U25 : AND2_X1 port map( A1 => net38998, A2 => n26, ZN => n5);
   U26 : AOI22_X1 port map( A1 => incom(0), A2 => net29471, B1 => insh(0), B2 
                           => net29483, ZN => n9);
   U27 : NAND2_X1 port map( A1 => n9, A2 => net27607, ZN => O(0));
   U28 : BUF_X1 port map( A => n1, Z => net29483);
   U29 : BUF_X1 port map( A => n1, Z => net29481);
   U30 : INV_X1 port map( A => sel(4), ZN => net27611);
   U31 : BUF_X1 port map( A => n8, Z => net29471);
   U32 : INV_X1 port map( A => net27616, ZN => n8);
   U33 : BUF_X1 port map( A => n8, Z => net29469);
   U34 : MUX2_X1 port map( A => n24, B => net27618, S => sel(1), Z => net27616)
                           ;
   U35 : OAI21_X1 port map( B1 => n3, B2 => n10, A => net25507, ZN => net27618)
                           ;
   U36 : NOR2_X1 port map( A1 => sel(4), A2 => sel(3), ZN => n10);
   U37 : AOI22_X1 port map( A1 => inlog(29), A2 => net29479, B1 => inadd(29), 
                           B2 => net29475, ZN => n25);
   U38 : NAND2_X1 port map( A1 => n25, A2 => net27572, ZN => O(29));
   U39 : INV_X2 port map( A => n26, ZN => net29475);
   U40 : INV_X2 port map( A => net39291, ZN => net29479);
   U41 : OAI211_X1 port map( C1 => n26, C2 => net39295, A => n4, B => net27574,
                           ZN => O(28));
   U42 : MUX2_X1 port map( A => n32, B => net39325, S => sel(1), Z => net39286)
                           ;
   U43 : MUX2_X1 port map( A => sel(2), B => n34, S => sel(3), Z => n31);
   U44 : AOI22_X1 port map( A1 => incom(29), A2 => net29471, B1 => insh(29), B2
                           => net29483, ZN => net27572);
   U45 : NOR2_X1 port map( A1 => inadd(27), A2 => n2, ZN => n36);
   U46 : INV_X1 port map( A => net27576, ZN => n37);
   U47 : INV_X1 port map( A => net38998, ZN => net38995);
   U48 : AND2_X1 port map( A1 => n5, A2 => net27576, ZN => n35);
   U49 : NOR2_X1 port map( A1 => n35, A2 => n36, ZN => O(27));
   U50 : INV_X1 port map( A => inadd(28), ZN => net39295);
   U51 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => O(9));
   U52 : AOI22_X1 port map( A1 => incom(9), A2 => net29469, B1 => insh(9), B2 
                           => net29481, ZN => n7);
   U53 : AOI22_X1 port map( A1 => inlog(9), A2 => net29479, B1 => inadd(9), B2 
                           => net29475, ZN => n6);
   U54 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => O(8));
   U55 : AOI22_X1 port map( A1 => incom(8), A2 => net29469, B1 => insh(8), B2 
                           => net29481, ZN => n13);
   U56 : AOI22_X1 port map( A1 => inlog(8), A2 => net29479, B1 => inadd(8), B2 
                           => net29475, ZN => n12);
   U57 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => O(10));
   U58 : AOI22_X1 port map( A1 => incom(10), A2 => net29469, B1 => insh(10), B2
                           => net29481, ZN => n71);
   U59 : AOI22_X1 port map( A1 => inlog(10), A2 => net29479, B1 => inadd(10), 
                           B2 => net29475, ZN => n70);
   U60 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => O(11));
   U61 : AOI22_X1 port map( A1 => incom(11), A2 => net29469, B1 => insh(11), B2
                           => net29481, ZN => n69);
   U62 : AOI22_X1 port map( A1 => inlog(11), A2 => net29479, B1 => inadd(11), 
                           B2 => net29475, ZN => n68);
   U63 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => O(7));
   U64 : AOI22_X1 port map( A1 => incom(7), A2 => net29469, B1 => insh(7), B2 
                           => net29481, ZN => n15);
   U65 : AOI22_X1 port map( A1 => inlog(7), A2 => net29479, B1 => inadd(7), B2 
                           => net29475, ZN => n14);
   U66 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => O(6));
   U67 : AOI22_X1 port map( A1 => incom(6), A2 => net29469, B1 => insh(6), B2 
                           => net29481, ZN => n17);
   U68 : AOI22_X1 port map( A1 => inlog(6), A2 => net29479, B1 => inadd(6), B2 
                           => net29475, ZN => n16);
   U69 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => O(4));
   U70 : AOI22_X1 port map( A1 => incom(4), A2 => net29469, B1 => insh(4), B2 
                           => net29481, ZN => n21);
   U71 : AOI22_X1 port map( A1 => inlog(4), A2 => net29479, B1 => inadd(4), B2 
                           => net29475, ZN => n20);
   U72 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => O(5));
   U73 : AOI22_X1 port map( A1 => incom(5), A2 => net29469, B1 => insh(5), B2 
                           => net29481, ZN => n19);
   U74 : AOI22_X1 port map( A1 => inlog(5), A2 => net29479, B1 => inadd(5), B2 
                           => net29475, ZN => n18);
   U75 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => O(1));
   U76 : AOI22_X1 port map( A1 => inlog(1), A2 => net29479, B1 => inadd(1), B2 
                           => net29475, ZN => n50);
   U77 : AOI22_X1 port map( A1 => incom(1), A2 => net29469, B1 => insh(1), B2 
                           => net29481, ZN => n51);
   U78 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => O(2));
   U79 : AOI22_X1 port map( A1 => inlog(2), A2 => net29479, B1 => inadd(2), B2 
                           => net29475, ZN => n28);
   U80 : AOI22_X1 port map( A1 => incom(2), A2 => net29469, B1 => insh(2), B2 
                           => net29481, ZN => n29);
   U81 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => O(3));
   U82 : AOI22_X1 port map( A1 => inlog(3), A2 => net29479, B1 => inadd(3), B2 
                           => net29475, ZN => n22);
   U83 : AOI22_X1 port map( A1 => incom(3), A2 => net29469, B1 => insh(3), B2 
                           => net29481, ZN => n23);
   U84 : AOI22_X1 port map( A1 => inlog(0), A2 => net29479, B1 => inadd(0), B2 
                           => net29475, ZN => net27607);
   U85 : AOI22_X1 port map( A1 => inlog(12), A2 => net29479, B1 => inadd(12), 
                           B2 => net29475, ZN => n39);
   U86 : AOI22_X1 port map( A1 => incom(12), A2 => net29471, B1 => insh(12), B2
                           => net29483, ZN => n38);
   U87 : NAND2_X1 port map( A1 => n39, A2 => n38, ZN => O(12));
   U88 : AOI22_X1 port map( A1 => inlog(13), A2 => net29479, B1 => inadd(13), 
                           B2 => net29475, ZN => n41);
   U89 : AOI22_X1 port map( A1 => incom(13), A2 => net29471, B1 => insh(13), B2
                           => net29483, ZN => n40);
   U90 : NAND2_X1 port map( A1 => n41, A2 => n40, ZN => O(13));
   U91 : AOI22_X1 port map( A1 => inlog(14), A2 => net29479, B1 => inadd(14), 
                           B2 => net29475, ZN => n43);
   U92 : AOI22_X1 port map( A1 => incom(14), A2 => net29471, B1 => insh(14), B2
                           => net29483, ZN => n42);
   U93 : NAND2_X1 port map( A1 => n43, A2 => n42, ZN => O(14));
   U94 : AOI22_X1 port map( A1 => inlog(15), A2 => net29479, B1 => inadd(15), 
                           B2 => net29475, ZN => n45);
   U95 : AOI22_X1 port map( A1 => incom(15), A2 => net29471, B1 => insh(15), B2
                           => net29483, ZN => n44);
   U96 : NAND2_X1 port map( A1 => n45, A2 => n44, ZN => O(15));
   U97 : AOI22_X1 port map( A1 => inlog(16), A2 => net29479, B1 => inadd(16), 
                           B2 => net29475, ZN => n47);
   U98 : AOI22_X1 port map( A1 => incom(16), A2 => net29471, B1 => insh(16), B2
                           => net29483, ZN => n46);
   U99 : NAND2_X1 port map( A1 => n47, A2 => n46, ZN => O(16));
   U100 : AOI22_X1 port map( A1 => inlog(17), A2 => net29479, B1 => inadd(17), 
                           B2 => net29475, ZN => n49);
   U101 : AOI22_X1 port map( A1 => incom(17), A2 => net29471, B1 => insh(17), 
                           B2 => net29483, ZN => n48);
   U102 : NAND2_X1 port map( A1 => n49, A2 => n48, ZN => O(17));
   U103 : AOI22_X1 port map( A1 => inlog(18), A2 => net29479, B1 => inadd(18), 
                           B2 => net29475, ZN => n53);
   U104 : AOI22_X1 port map( A1 => incom(18), A2 => net29471, B1 => insh(18), 
                           B2 => net29483, ZN => n52);
   U105 : NAND2_X1 port map( A1 => n53, A2 => n52, ZN => O(18));
   U106 : AOI22_X1 port map( A1 => inlog(19), A2 => net29479, B1 => inadd(19), 
                           B2 => net29475, ZN => n55);
   U107 : AOI22_X1 port map( A1 => incom(19), A2 => net29471, B1 => insh(19), 
                           B2 => net29483, ZN => n54);
   U108 : NAND2_X1 port map( A1 => n55, A2 => n54, ZN => O(19));
   U109 : AOI22_X1 port map( A1 => inlog(20), A2 => net29479, B1 => inadd(20), 
                           B2 => net29475, ZN => n57);
   U110 : AOI22_X1 port map( A1 => incom(20), A2 => net29471, B1 => insh(20), 
                           B2 => net29483, ZN => n56);
   U111 : NAND2_X1 port map( A1 => n57, A2 => n56, ZN => O(20));
   U112 : AOI22_X1 port map( A1 => inlog(21), A2 => net29479, B1 => inadd(21), 
                           B2 => net29475, ZN => n59);
   U113 : AOI22_X1 port map( A1 => incom(21), A2 => net29471, B1 => insh(21), 
                           B2 => net29483, ZN => n58);
   U114 : NAND2_X1 port map( A1 => n59, A2 => n58, ZN => O(21));
   U115 : AOI22_X1 port map( A1 => inlog(22), A2 => net29479, B1 => inadd(22), 
                           B2 => net29475, ZN => n61);
   U116 : AOI22_X1 port map( A1 => incom(22), A2 => net29471, B1 => insh(22), 
                           B2 => net29483, ZN => n60);
   U117 : NAND2_X1 port map( A1 => n61, A2 => n60, ZN => O(22));
   U118 : AOI22_X1 port map( A1 => inlog(23), A2 => net29479, B1 => inadd(23), 
                           B2 => net29475, ZN => n63);
   U119 : AOI22_X1 port map( A1 => incom(23), A2 => net29471, B1 => insh(23), 
                           B2 => net29483, ZN => n62);
   U120 : NAND2_X1 port map( A1 => n63, A2 => n62, ZN => O(23));
   U121 : AOI22_X1 port map( A1 => inlog(24), A2 => net29479, B1 => inadd(24), 
                           B2 => net29475, ZN => n65);
   U122 : AOI22_X1 port map( A1 => incom(24), A2 => net29471, B1 => insh(24), 
                           B2 => net29483, ZN => n64);
   U123 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => O(24));
   U124 : AOI22_X1 port map( A1 => inlog(25), A2 => net29479, B1 => inadd(25), 
                           B2 => net29475, ZN => n67);
   U125 : AOI22_X1 port map( A1 => incom(25), A2 => net29471, B1 => insh(25), 
                           B2 => net29483, ZN => n66);
   U126 : NAND2_X1 port map( A1 => n67, A2 => n66, ZN => O(25));
   U127 : AOI22_X1 port map( A1 => inlog(26), A2 => net29479, B1 => inadd(26), 
                           B2 => net29475, ZN => n73);
   U128 : AOI22_X1 port map( A1 => incom(26), A2 => net29471, B1 => insh(26), 
                           B2 => net29483, ZN => n72);
   U129 : NAND2_X1 port map( A1 => n73, A2 => n72, ZN => O(26));
   U130 : AOI22_X1 port map( A1 => incom(27), A2 => net29471, B1 => insh(27), 
                           B2 => net29483, ZN => net27576);
   U131 : AOI22_X1 port map( A1 => incom(28), A2 => net29471, B1 => insh(28), 
                           B2 => net29483, ZN => net27574);
   U132 : AOI22_X1 port map( A1 => inlog(30), A2 => net29479, B1 => inadd(30), 
                           B2 => net29475, ZN => n75);
   U133 : AOI22_X1 port map( A1 => incom(30), A2 => net29471, B1 => insh(30), 
                           B2 => net29483, ZN => n74);
   U134 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => O(30));
   U135 : AOI22_X1 port map( A1 => inlog(31), A2 => net29479, B1 => inadd(31), 
                           B2 => net29475, ZN => n77);
   U136 : AOI22_X1 port map( A1 => incom(31), A2 => net29469, B1 => insh(31), 
                           B2 => net29481, ZN => n76);
   U137 : NAND2_X1 port map( A1 => n77, A2 => n76, ZN => O(31));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity comparator_N32 is

   port( inA, inB : in std_logic_vector (31 downto 0);  op : in 
         std_logic_vector (0 to 4);  res : out std_logic_vector (31 downto 0));

end comparator_N32;

architecture SYN_Behavioral of comparator_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_N32_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   signal X_Logic0_port, res_0_port, N8, n13, net27627, net27642, net27652, 
      net27653, net27661, net27665, net27668, net27736, net27753, net36280, 
      net36538, net36884, net36937, net36956, net36967, net36976, net37153, 
      net37179, net37323, net37334, net37410, net37531, net37588, net37593, 
      net37592, net37658, net37657, net37746, net37745, net38175, net38169, 
      net38153, net27641, net27636, net27650, net27647, net27646, net27644, 
      net37765, net37406, net36906, net27658, net27657, net27655, net35853, 
      net35852, net29761, net27659, net27651, net27649, net27648, net27645, 
      net27643, net27640, net27639, net27637, net27635, net27632, net27631, 
      net27630, net27629, net27628, net38080, n1, n2, n3, n4, n5, n6, n7, 
      n8_port, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n_1139,
      n_1140, n_1141, n_1142, n_1143 : std_logic;

begin
   res <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, res_0_port 
      );
   
   X_Logic0_port <= '0';
   n13 <= '0';
   r57 : comparator_N32_DW01_cmp6_0 port map( A(31) => inA(31), A(30) => 
                           inA(30), A(29) => inA(29), A(28) => inA(28), A(27) 
                           => inA(27), A(26) => inA(26), A(25) => inA(25), 
                           A(24) => inA(24), A(23) => inA(23), A(22) => inA(22)
                           , A(21) => inA(21), A(20) => inA(20), A(19) => 
                           inA(19), A(18) => inA(18), A(17) => inA(17), A(16) 
                           => inA(16), A(15) => inA(15), A(14) => inA(14), 
                           A(13) => inA(13), A(12) => inA(12), A(11) => inA(11)
                           , A(10) => inA(10), A(9) => inA(9), A(8) => inA(8), 
                           A(7) => inA(7), A(6) => inA(6), A(5) => inA(5), A(4)
                           => inA(4), A(3) => inA(3), A(2) => inA(2), A(1) => 
                           inA(1), A(0) => inA(0), B(31) => inB(31), B(30) => 
                           inB(30), B(29) => inB(29), B(28) => inB(28), B(27) 
                           => inB(27), B(26) => inB(26), B(25) => inB(25), 
                           B(24) => inB(24), B(23) => inB(23), B(22) => inB(22)
                           , B(21) => inB(21), B(20) => inB(20), B(19) => 
                           inB(19), B(18) => inB(18), B(17) => inB(17), B(16) 
                           => inB(16), B(15) => inB(15), B(14) => inB(14), 
                           B(13) => inB(13), B(12) => inB(12), B(11) => inB(11)
                           , B(10) => inB(10), B(9) => inB(9), B(8) => inB(8), 
                           B(7) => inB(7), B(6) => inB(6), B(5) => inB(5), B(4)
                           => inB(4), B(3) => inB(3), B(2) => inB(2), B(1) => 
                           inB(1), B(0) => net36956, TC => n13, LT => n_1139, 
                           GT => n_1140, EQ => N8, LE => n_1141, GE => n_1142, 
                           NE => n_1143);
   U2 : OR2_X2 port map( A1 => net37593, A2 => net37334, ZN => net37592);
   U3 : INV_X1 port map( A => inB(5), ZN => n41);
   U4 : OR2_X1 port map( A1 => n23, A2 => n108, ZN => net36976);
   U5 : NAND2_X1 port map( A1 => net37153, A2 => net36976, ZN => n22);
   U6 : INV_X1 port map( A => net36976, ZN => net37593);
   U7 : NAND2_X1 port map( A1 => n16, A2 => n27, ZN => net37746);
   U8 : INV_X1 port map( A => net37153, ZN => n16);
   U10 : INV_X1 port map( A => inB(30), ZN => n25);
   U11 : INV_X1 port map( A => inB(2), ZN => net38175);
   U12 : INV_X1 port map( A => inB(4), ZN => n42);
   U13 : NAND2_X1 port map( A1 => n41, A2 => inA(5), ZN => net36937);
   U14 : NAND2_X1 port map( A1 => inB(28), A2 => net27668, ZN => n24);
   U15 : INV_X1 port map( A => inB(29), ZN => n21);
   U16 : INV_X1 port map( A => n22, ZN => net37531);
   U17 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => net37765);
   U18 : NAND2_X1 port map( A1 => net37588, A2 => n4, ZN => net37406);
   U19 : OAI21_X1 port map( B1 => net37765, B2 => net27659, A => net27658, ZN 
                           => net27639);
   U20 : NAND2_X1 port map( A1 => net37323, A2 => n4, ZN => net36906);
   U21 : AND2_X1 port map( A1 => n127, A2 => n128, ZN => n1);
   U22 : AND2_X1 port map( A1 => n125, A2 => n126, ZN => n2);
   U23 : AND2_X1 port map( A1 => n89, A2 => n90, ZN => n3);
   U24 : AND2_X1 port map( A1 => n19, A2 => n20, ZN => n4);
   U25 : AND2_X1 port map( A1 => n102, A2 => n103, ZN => n5);
   U26 : AND2_X1 port map( A1 => net27643, A2 => op(3), ZN => n6);
   U27 : AND2_X1 port map( A1 => net27643, A2 => op(4), ZN => n7);
   U28 : INV_X1 port map( A => n23, ZN => net36280);
   U29 : OAI211_X1 port map( C1 => inA(29), C2 => n21, A => n24, B => net27665,
                           ZN => n23);
   U30 : AND2_X1 port map( A1 => n129, A2 => n130, ZN => n8_port);
   U31 : AND2_X1 port map( A1 => n69, A2 => n68, ZN => n9);
   U32 : AND2_X1 port map( A1 => n105, A2 => n104, ZN => n10);
   U33 : AND2_X1 port map( A1 => n78, A2 => n79, ZN => n11);
   U34 : AND2_X1 port map( A1 => n100, A2 => n101, ZN => n12);
   U35 : AND2_X1 port map( A1 => n120, A2 => n119, ZN => n14);
   U36 : AND2_X1 port map( A1 => n99, A2 => n98, ZN => n15);
   U37 : NAND3_X1 port map( A1 => net37410, A2 => n27, A3 => net37179, ZN => 
                           net37745);
   U38 : NAND3_X1 port map( A1 => inA(29), A2 => n21, A3 => net27665, ZN => n20
                           );
   U39 : NAND3_X1 port map( A1 => net37410, A2 => net37592, A3 => net37179, ZN 
                           => n18);
   U40 : NAND2_X1 port map( A1 => inA(30), A2 => n25, ZN => n19);
   U41 : INV_X1 port map( A => inA(30), ZN => net27661);
   U42 : BUF_X1 port map( A => net37334, Z => n27);
   U43 : AND2_X1 port map( A1 => net37592, A2 => net37410, ZN => net37658);
   U44 : NAND2_X1 port map( A1 => net37592, A2 => n22, ZN => n26);
   U45 : AND2_X1 port map( A1 => n4, A2 => n26, ZN => n17);
   U46 : AOI21_X1 port map( B1 => n31, B2 => net38080, A => inB(1), ZN => n28);
   U47 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => net38153);
   U48 : INV_X1 port map( A => inA(1), ZN => net38080);
   U49 : OAI22_X1 port map( A1 => n32, A2 => net38080, B1 => inB(2), B2 => 
                           net38169, ZN => n29);
   U50 : NOR2_X1 port map( A1 => inA(0), A2 => n30, ZN => n31);
   U51 : INV_X1 port map( A => inB(0), ZN => n30);
   U52 : NOR2_X1 port map( A1 => inA(0), A2 => n30, ZN => n32);
   U53 : OAI211_X1 port map( C1 => net27627, C2 => net27628, A => net27630, B 
                           => net27629, ZN => res_0_port);
   U54 : OAI211_X1 port map( C1 => op(4), C2 => net27643, A => net27648, B => 
                           net27649, ZN => net27629);
   U55 : NAND2_X1 port map( A1 => net36967, A2 => n7, ZN => net27649);
   U56 : INV_X1 port map( A => N8, ZN => net27643);
   U57 : NAND2_X1 port map( A1 => net36884, A2 => net27643, ZN => net27632);
   U58 : NOR4_X1 port map( A1 => op(3), A2 => op(2), A3 => op(0), A4 => 
                           net27651, ZN => net27648);
   U59 : INV_X1 port map( A => op(1), ZN => net27651);
   U60 : NAND2_X1 port map( A1 => op(0), A2 => net27651, ZN => net27627);
   U61 : NOR3_X1 port map( A1 => n34, A2 => net27635, A3 => net29761, ZN => 
                           net27630);
   U62 : NOR2_X1 port map( A1 => net35852, A2 => net35853, ZN => net29761);
   U63 : OR3_X1 port map( A1 => net27644, A2 => op(0), A3 => net27640, ZN => 
                           net35853);
   U64 : INV_X1 port map( A => op(3), ZN => net27640);
   U65 : NAND2_X1 port map( A1 => op(4), A2 => net27640, ZN => net27637);
   U66 : NOR2_X1 port map( A1 => net27650, A2 => N8, ZN => net35852);
   U67 : OAI33_X1 port map( A1 => net27636, A2 => net27637, A3 => net27632, B1 
                           => n33, B2 => op(4), B3 => net27636, ZN => net27635)
                           ;
   U68 : AOI21_X1 port map( B1 => net27639, B2 => op(3), A => N8, ZN => n33);
   U69 : INV_X1 port map( A => net27657, ZN => net27659);
   U70 : OAI21_X1 port map( B1 => net36906, B2 => net27659, A => net27658, ZN 
                           => net36884);
   U71 : AND2_X1 port map( A1 => net27632, A2 => net27631, ZN => n34);
   U72 : NOR3_X1 port map( A1 => net27644, A2 => op(3), A3 => net27645, ZN => 
                           net27631);
   U73 : INV_X1 port map( A => op(0), ZN => net27645);
   U74 : NAND3_X1 port map( A1 => net27652, A2 => net27653, A3 => n6, ZN => 
                           net27628);
   U75 : NAND2_X1 port map( A1 => inB(31), A2 => n35, ZN => net27658);
   U76 : INV_X1 port map( A => net27658, ZN => net27655);
   U77 : INV_X1 port map( A => inA(31), ZN => n35);
   U78 : NAND2_X1 port map( A1 => inA(31), A2 => n36, ZN => net27657);
   U79 : OAI21_X1 port map( B1 => net37406, B2 => net27655, A => net27657, ZN 
                           => net27650);
   U80 : OAI21_X1 port map( B1 => net27655, B2 => net37765, A => net27657, ZN 
                           => net36967);
   U81 : INV_X1 port map( A => inB(31), ZN => n36);
   U82 : NAND3_X1 port map( A1 => op(1), A2 => net27646, A3 => net27647, ZN => 
                           net27644);
   U83 : INV_X1 port map( A => op(2), ZN => net27647);
   U84 : INV_X1 port map( A => op(4), ZN => net27646);
   U85 : NOR2_X1 port map( A1 => op(2), A2 => net27646, ZN => n37);
   U86 : OAI21_X1 port map( B1 => op(2), B2 => net27642, A => net27646, ZN => 
                           net27653);
   U87 : AOI22_X1 port map( A1 => op(2), A2 => net36884, B1 => net27650, B2 => 
                           n37, ZN => net27652);
   U88 : NAND2_X1 port map( A1 => op(2), A2 => net27641, ZN => net27636);
   U89 : INV_X1 port map( A => net27627, ZN => net27641);
   U90 : NOR2_X1 port map( A1 => n38, A2 => net37593, ZN => net37588);
   U91 : NAND2_X1 port map( A1 => net37745, A2 => net37746, ZN => n38);
   U92 : NAND2_X1 port map( A1 => n57, A2 => n55, ZN => n39);
   U93 : NAND2_X1 port map( A1 => n1, A2 => n40, ZN => n84);
   U94 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => n40);
   U95 : NAND2_X1 port map( A1 => inA(3), A2 => n48, ZN => n50);
   U96 : INV_X1 port map( A => inB(3), ZN => n48);
   U97 : NAND2_X1 port map( A1 => inB(5), A2 => n47, ZN => n43);
   U98 : OAI21_X1 port map( B1 => inA(4), B2 => n42, A => n43, ZN => n51);
   U99 : OAI22_X1 port map( A1 => inA(2), A2 => net38175, B1 => inA(3), B2 => 
                           n48, ZN => n49);
   U100 : OAI21_X1 port map( B1 => net38153, B2 => n49, A => n50, ZN => n44);
   U101 : NOR2_X1 port map( A1 => n51, A2 => net36538, ZN => n46);
   U102 : AOI21_X1 port map( B1 => n44, B2 => n45, A => n46, ZN => net27736);
   U103 : INV_X1 port map( A => n51, ZN => n45);
   U104 : INV_X1 port map( A => inA(5), ZN => n47);
   U105 : INV_X1 port map( A => inA(4), ZN => net27753);
   U106 : INV_X1 port map( A => inA(2), ZN => net38169);
   U107 : INV_X1 port map( A => n30, ZN => net36956);
   U108 : NAND2_X1 port map( A1 => n39, A2 => n5, ZN => n52);
   U109 : AND2_X1 port map( A1 => n83, A2 => n75, ZN => n53);
   U110 : NOR2_X1 port map( A1 => n53, A2 => n54, ZN => net37410);
   U111 : NOR2_X1 port map( A1 => n82, A2 => n85, ZN => n54);
   U112 : AND2_X1 port map( A1 => n58, A2 => n9, ZN => n55);
   U113 : NAND2_X1 port map( A1 => n52, A2 => n70, ZN => n56);
   U114 : AND2_X1 port map( A1 => n109, A2 => n84, ZN => n83);
   U115 : NAND2_X1 port map( A1 => n72, A2 => n59, ZN => n57);
   U116 : OR2_X1 port map( A1 => n62, A2 => n3, ZN => n58);
   U117 : AND2_X1 port map( A1 => n64, A2 => n63, ZN => n59);
   U118 : NAND2_X1 port map( A1 => n56, A2 => net37658, ZN => n60);
   U119 : AND2_X1 port map( A1 => n60, A2 => n61, ZN => net37323);
   U120 : OR2_X1 port map( A1 => net37657, A2 => net37531, ZN => n61);
   U121 : INV_X1 port map( A => net37592, ZN => net37657);
   U122 : NAND2_X1 port map( A1 => n81, A2 => n80, ZN => n62);
   U123 : INV_X1 port map( A => n62, ZN => n63);
   U124 : AND2_X1 port map( A1 => n71, A2 => n86, ZN => net37334);
   U125 : AND2_X1 port map( A1 => n73, A2 => n10, ZN => n64);
   U126 : NOR2_X1 port map( A1 => n66, A2 => n67, ZN => n65);
   U127 : NOR2_X1 port map( A1 => inA(6), A2 => n133, ZN => n66);
   U128 : NOR2_X1 port map( A1 => inA(7), A2 => n134, ZN => n67);
   U129 : OR2_X1 port map( A1 => inB(16), A2 => n155, ZN => n68);
   U130 : OR2_X1 port map( A1 => inB(15), A2 => n154, ZN => n69);
   U131 : NAND2_X1 port map( A1 => n52, A2 => n70, ZN => net37179);
   U132 : AND2_X1 port map( A1 => n106, A2 => n83, ZN => n70);
   U133 : OR2_X1 port map( A1 => n76, A2 => n2, ZN => n71);
   U134 : AND2_X1 port map( A1 => n11, A2 => n77, ZN => net37153);
   U135 : NAND2_X1 port map( A1 => n141, A2 => n74, ZN => n72);
   U136 : OR2_X1 port map( A1 => n110, A2 => n87, ZN => n73);
   U137 : AND2_X1 port map( A1 => n14, A2 => n88, ZN => n74);
   U138 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => n75);
   U139 : NAND2_X1 port map( A1 => n138, A2 => n8_port, ZN => n141);
   U140 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => n76);
   U141 : INV_X1 port map( A => n76, ZN => n77);
   U142 : OR2_X1 port map( A1 => inB(26), A2 => n175, ZN => n91);
   U143 : OR2_X1 port map( A1 => inB(14), A2 => n151, ZN => n89);
   U144 : OR2_X1 port map( A1 => inB(24), A2 => n171, ZN => n78);
   U145 : OR2_X1 port map( A1 => inB(23), A2 => n170, ZN => n79);
   U146 : OR2_X1 port map( A1 => inA(15), A2 => n153, ZN => n80);
   U147 : OR2_X1 port map( A1 => inA(14), A2 => n152, ZN => n81);
   U148 : INV_X1 port map( A => n84, ZN => n82);
   U149 : NAND2_X1 port map( A1 => n132, A2 => n65, ZN => n135);
   U150 : AND2_X1 port map( A1 => n12, A2 => n1, ZN => n85);
   U151 : AND2_X1 port map( A1 => n15, A2 => net36280, ZN => n86);
   U152 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => n87);
   U153 : INV_X1 port map( A => n87, ZN => n88);
   U154 : OR2_X1 port map( A1 => inB(12), A2 => n147, ZN => n94);
   U155 : OR2_X1 port map( A1 => inB(13), A2 => n150, ZN => n90);
   U156 : OR2_X1 port map( A1 => inB(25), A2 => n174, ZN => n92);
   U157 : OR2_X1 port map( A1 => inB(6), A2 => n131, ZN => n93);
   U158 : NAND3_X1 port map( A1 => net27736, A2 => net36937, A3 => n93, ZN => 
                           n132);
   U159 : OR2_X1 port map( A1 => inB(11), A2 => n146, ZN => n95);
   U160 : OR2_X1 port map( A1 => inA(19), A2 => n161, ZN => n96);
   U161 : OR2_X1 port map( A1 => inA(18), A2 => n160, ZN => n97);
   U162 : OR2_X1 port map( A1 => inA(27), A2 => n177, ZN => n98);
   U163 : OR2_X1 port map( A1 => inA(26), A2 => n176, ZN => n99);
   U164 : OR2_X1 port map( A1 => inA(21), A2 => n165, ZN => n100);
   U165 : OR2_X1 port map( A1 => inA(20), A2 => n164, ZN => n101);
   U166 : OR2_X1 port map( A1 => inA(17), A2 => n157, ZN => n102);
   U167 : OR2_X1 port map( A1 => inA(16), A2 => n156, ZN => n103);
   U168 : OR2_X1 port map( A1 => inA(13), A2 => n149, ZN => n104);
   U169 : OR2_X1 port map( A1 => inA(12), A2 => n148, ZN => n105);
   U170 : OR2_X1 port map( A1 => inB(4), A2 => net27753, ZN => net36538);
   U171 : AND2_X1 port map( A1 => n114, A2 => n113, ZN => n106);
   U172 : AND2_X1 port map( A1 => n116, A2 => n115, ZN => n107);
   U173 : AND2_X1 port map( A1 => n121, A2 => n122, ZN => n108);
   U174 : AND2_X1 port map( A1 => n118, A2 => n117, ZN => n109);
   U175 : NOR2_X1 port map( A1 => n111, A2 => n112, ZN => n110);
   U176 : NOR2_X1 port map( A1 => n144, A2 => inA(10), ZN => n111);
   U177 : NOR2_X1 port map( A1 => inA(11), A2 => n145, ZN => n112);
   U178 : NAND2_X1 port map( A1 => n135, A2 => n107, ZN => n138);
   U179 : OR2_X1 port map( A1 => inB(18), A2 => n159, ZN => n113);
   U180 : OR2_X1 port map( A1 => inB(17), A2 => n158, ZN => n114);
   U181 : OR2_X1 port map( A1 => inB(8), A2 => n137, ZN => n115);
   U182 : OR2_X1 port map( A1 => inB(7), A2 => n136, ZN => n116);
   U183 : OR2_X1 port map( A1 => inB(20), A2 => n163, ZN => n117);
   U184 : OR2_X1 port map( A1 => inB(19), A2 => n162, ZN => n118);
   U185 : OR2_X1 port map( A1 => inB(10), A2 => n143, ZN => n119);
   U186 : OR2_X1 port map( A1 => inB(9), A2 => n142, ZN => n120);
   U187 : OR2_X1 port map( A1 => inB(28), A2 => net27668, ZN => n121);
   U188 : OR2_X1 port map( A1 => inB(27), A2 => n178, ZN => n122);
   U189 : OR2_X1 port map( A1 => inB(22), A2 => n167, ZN => n123);
   U190 : OR2_X1 port map( A1 => inB(21), A2 => n166, ZN => n124);
   U191 : OR2_X1 port map( A1 => inA(25), A2 => n173, ZN => n125);
   U192 : OR2_X1 port map( A1 => inA(24), A2 => n172, ZN => n126);
   U193 : OR2_X1 port map( A1 => inA(23), A2 => n169, ZN => n127);
   U194 : OR2_X1 port map( A1 => inA(22), A2 => n168, ZN => n128);
   U195 : OR2_X1 port map( A1 => inA(9), A2 => n140, ZN => n129);
   U196 : OR2_X1 port map( A1 => inA(8), A2 => n139, ZN => n130);
   U197 : NAND2_X1 port map( A1 => inB(30), A2 => net27661, ZN => net27665);
   U198 : INV_X1 port map( A => inA(28), ZN => net27668);
   U199 : INV_X1 port map( A => inA(27), ZN => n178);
   U200 : INV_X1 port map( A => inB(27), ZN => n177);
   U201 : INV_X1 port map( A => inB(26), ZN => n176);
   U202 : INV_X1 port map( A => inA(26), ZN => n175);
   U203 : INV_X1 port map( A => inA(25), ZN => n174);
   U204 : INV_X1 port map( A => inB(25), ZN => n173);
   U205 : INV_X1 port map( A => inB(24), ZN => n172);
   U206 : INV_X1 port map( A => inA(24), ZN => n171);
   U207 : INV_X1 port map( A => inA(23), ZN => n170);
   U208 : INV_X1 port map( A => inB(23), ZN => n169);
   U209 : INV_X1 port map( A => inB(22), ZN => n168);
   U210 : INV_X1 port map( A => inA(22), ZN => n167);
   U211 : INV_X1 port map( A => inA(21), ZN => n166);
   U212 : INV_X1 port map( A => inB(21), ZN => n165);
   U213 : INV_X1 port map( A => inB(20), ZN => n164);
   U214 : INV_X1 port map( A => inA(20), ZN => n163);
   U215 : INV_X1 port map( A => inA(19), ZN => n162);
   U216 : INV_X1 port map( A => inB(19), ZN => n161);
   U217 : INV_X1 port map( A => inB(18), ZN => n160);
   U218 : INV_X1 port map( A => inA(18), ZN => n159);
   U219 : INV_X1 port map( A => inA(17), ZN => n158);
   U220 : INV_X1 port map( A => inB(17), ZN => n157);
   U221 : INV_X1 port map( A => inB(16), ZN => n156);
   U222 : INV_X1 port map( A => inA(16), ZN => n155);
   U223 : INV_X1 port map( A => inA(15), ZN => n154);
   U224 : INV_X1 port map( A => inB(15), ZN => n153);
   U225 : INV_X1 port map( A => inB(14), ZN => n152);
   U226 : INV_X1 port map( A => inA(14), ZN => n151);
   U227 : INV_X1 port map( A => inA(13), ZN => n150);
   U228 : INV_X1 port map( A => inB(13), ZN => n149);
   U229 : INV_X1 port map( A => inB(12), ZN => n148);
   U230 : INV_X1 port map( A => inA(12), ZN => n147);
   U231 : INV_X1 port map( A => inA(11), ZN => n146);
   U232 : INV_X1 port map( A => inB(11), ZN => n145);
   U233 : INV_X1 port map( A => inB(10), ZN => n144);
   U234 : INV_X1 port map( A => inA(10), ZN => n143);
   U235 : INV_X1 port map( A => inA(9), ZN => n142);
   U236 : INV_X1 port map( A => inB(9), ZN => n140);
   U237 : INV_X1 port map( A => inB(8), ZN => n139);
   U238 : INV_X1 port map( A => inA(8), ZN => n137);
   U239 : INV_X1 port map( A => inA(7), ZN => n136);
   U240 : INV_X1 port map( A => inB(7), ZN => n134);
   U241 : INV_X1 port map( A => inB(6), ZN => n133);
   U242 : INV_X1 port map( A => inA(6), ZN => n131);
   U243 : INV_X1 port map( A => net36967, ZN => net27642);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SHIFTER_GENERIC_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (0 to 4);  OUTPUT : out std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32;

architecture SYN_BEHAVIORAL of SHIFTER_GENERIC_N32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
      N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46
      , N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, 
      N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75
      , N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, 
      N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
      N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, n7, n8, n9, 
      n13, n14, n15, n16, n17, n18_port, n19_port, n20_port, n21_port, n22_port
      , n23_port, n24_port, n25_port, n26_port, n27_port, n28_port, n29_port, 
      n30_port, n31_port, n32_port, n33_port, n34_port, n35_port, n36_port, 
      n37_port, n38_port, n39_port, n40_port, n41_port, n42_port, n43_port, 
      n44_port, n45_port, n46_port, n47_port, n48_port, n49_port, n50_port, 
      n51_port, n52_port, n53_port, n54_port, n55_port, n56_port, n57_port, 
      n58_port, n59_port, n60_port, n61_port, n62_port, n63_port, n64_port, 
      n65_port, n66_port, n67_port, n68_port, n69_port, n70_port, n71_port, 
      n72_port, n73_port, n74_port, n75_port, n76_port, n77_port, n78_port, 
      n79_port, n80_port, n81_port, n1, n2, n3, n4, n5, n6, n10, n11, n12, 
      n82_port, n83_port, n84_port, n85_port, n86_port, n87_port, n88_port : 
      std_logic;

begin
   
   n7 <= '0';
   n8 <= '0';
   n9 <= '0';
   U110 : NAND3_X1 port map( A1 => sel(3), A2 => n87_port, A3 => sel(2), ZN => 
                           n81_port);
   sra_28 : SHIFTER_GENERIC_N32_DW_sra_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n85_port, SH(3) => 
                           B(3), SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), 
                           SH_TC => n7, B(31) => N113, B(30) => N112, B(29) => 
                           N111, B(28) => N110, B(27) => N109, B(26) => N108, 
                           B(25) => N107, B(24) => N106, B(23) => N105, B(22) 
                           => N104, B(21) => N103, B(20) => N102, B(19) => N101
                           , B(18) => N100, B(17) => N99, B(16) => N98, B(15) 
                           => N97, B(14) => N96, B(13) => N95, B(12) => N94, 
                           B(11) => N93, B(10) => N92, B(9) => N91, B(8) => N90
                           , B(7) => N89, B(6) => N88, B(5) => N87, B(4) => N86
                           , B(3) => N85, B(2) => N84, B(1) => N83, B(0) => N82
                           );
   srl_26 : SHIFTER_GENERIC_N32_DW_rash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n8, SH(4) => 
                           n85_port, SH(3) => B(3), SH(2) => B(2), SH(1) => 
                           B(1), SH(0) => B(0), SH_TC => n8, B(31) => N81, 
                           B(30) => N80, B(29) => N79, B(28) => N78, B(27) => 
                           N77, B(26) => N76, B(25) => N75, B(24) => N74, B(23)
                           => N73, B(22) => N72, B(21) => N71, B(20) => N70, 
                           B(19) => N69, B(18) => N68, B(17) => N67, B(16) => 
                           N66, B(15) => N65, B(14) => N64, B(13) => N63, B(12)
                           => N62, B(11) => N61, B(10) => N60, B(9) => N59, 
                           B(8) => N58, B(7) => N57, B(6) => N56, B(5) => N55, 
                           B(4) => N54, B(3) => N53, B(2) => N52, B(1) => N51, 
                           B(0) => N50);
   sll_27 : SHIFTER_GENERIC_N32_DW01_ash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n9, SH(4) => 
                           n85_port, SH(3) => B(3), SH(2) => B(2), SH(1) => 
                           B(1), SH(0) => B(0), SH_TC => n9, B(31) => N49, 
                           B(30) => N48, B(29) => N47, B(28) => N46, B(27) => 
                           N45, B(26) => N44, B(25) => N43, B(24) => N42, B(23)
                           => N41, B(22) => N40, B(21) => N39, B(20) => N38, 
                           B(19) => N37, B(18) => N36, B(17) => N35, B(16) => 
                           N34, B(15) => N33, B(14) => N32, B(13) => N31, B(12)
                           => N30, B(11) => N29, B(10) => N28, B(9) => N27, 
                           B(8) => N26, B(7) => N25, B(6) => N24, B(5) => N23, 
                           B(4) => N22, B(3) => N21, B(2) => N20, B(1) => N19, 
                           B(0) => N18);
   U3 : BUF_X4 port map( A => B(4), Z => n85_port);
   U4 : AOI22_X1 port map( A1 => N87, A2 => n84_port, B1 => N55, B2 => n12, ZN 
                           => n26_port);
   U5 : AOI22_X1 port map( A1 => N86, A2 => n84_port, B1 => N54, B2 => n12, ZN 
                           => n28_port);
   U7 : AOI22_X1 port map( A1 => N88, A2 => n84_port, B1 => N56, B2 => n12, ZN 
                           => n24_port);
   U8 : AOI22_X1 port map( A1 => N91, A2 => n84_port, B1 => N59, B2 => n12, ZN 
                           => n14);
   U9 : AOI22_X1 port map( A1 => N90, A2 => n84_port, B1 => N58, B2 => n12, ZN 
                           => n20_port);
   U10 : AOI22_X1 port map( A1 => N89, A2 => n84_port, B1 => N57, B2 => n12, ZN
                           => n22_port);
   U11 : AOI22_X1 port map( A1 => N110, A2 => n83_port, B1 => N78, B2 => n11, 
                           ZN => n40_port);
   U12 : AOI22_X1 port map( A1 => N111, A2 => n83_port, B1 => N79, B2 => n11, 
                           ZN => n38_port);
   U13 : AOI22_X1 port map( A1 => N112, A2 => n83_port, B1 => N80, B2 => n11, 
                           ZN => n34_port);
   U14 : AOI22_X1 port map( A1 => N104, A2 => n83_port, B1 => N72, B2 => n11, 
                           ZN => n52_port);
   U15 : AOI22_X1 port map( A1 => N105, A2 => n83_port, B1 => N73, B2 => n11, 
                           ZN => n50_port);
   U16 : AOI22_X1 port map( A1 => N106, A2 => n83_port, B1 => N74, B2 => n11, 
                           ZN => n48_port);
   U17 : AOI22_X1 port map( A1 => N107, A2 => n83_port, B1 => N75, B2 => n11, 
                           ZN => n46_port);
   U18 : AOI22_X1 port map( A1 => N108, A2 => n83_port, B1 => N76, B2 => n11, 
                           ZN => n44_port);
   U19 : AOI22_X1 port map( A1 => N95, A2 => n82_port, B1 => N63, B2 => n10, ZN
                           => n72_port);
   U20 : AOI22_X1 port map( A1 => N96, A2 => n82_port, B1 => N64, B2 => n10, ZN
                           => n70_port);
   U21 : AOI22_X1 port map( A1 => N97, A2 => n82_port, B1 => N65, B2 => n10, ZN
                           => n68_port);
   U22 : AOI22_X1 port map( A1 => N93, A2 => n82_port, B1 => N61, B2 => n10, ZN
                           => n76_port);
   U23 : AOI22_X1 port map( A1 => N92, A2 => n82_port, B1 => N60, B2 => n10, ZN
                           => n78_port);
   U24 : AOI22_X1 port map( A1 => N94, A2 => n82_port, B1 => N62, B2 => n10, ZN
                           => n74_port);
   U25 : AOI22_X1 port map( A1 => N99, A2 => n82_port, B1 => N67, B2 => n10, ZN
                           => n64_port);
   U26 : AOI22_X1 port map( A1 => N98, A2 => n82_port, B1 => N66, B2 => n10, ZN
                           => n66_port);
   U27 : AOI22_X1 port map( A1 => N100, A2 => n82_port, B1 => N68, B2 => n10, 
                           ZN => n62_port);
   U28 : AOI22_X1 port map( A1 => N102, A2 => n83_port, B1 => N70, B2 => n11, 
                           ZN => n56_port);
   U29 : AOI22_X1 port map( A1 => N101, A2 => n82_port, B1 => N69, B2 => n10, 
                           ZN => n60_port);
   U30 : AOI22_X1 port map( A1 => N103, A2 => n83_port, B1 => N71, B2 => n11, 
                           ZN => n54_port);
   U31 : NAND2_X1 port map( A1 => n57_port, A2 => n58_port, ZN => OUTPUT(1));
   U32 : AOI22_X1 port map( A1 => N83, A2 => n82_port, B1 => N51, B2 => n10, ZN
                           => n58_port);
   U33 : NAND2_X1 port map( A1 => n29_port, A2 => n30_port, ZN => OUTPUT(3));
   U34 : AOI22_X1 port map( A1 => N21, A2 => n6, B1 => A(3), B2 => n3, ZN => 
                           n29_port);
   U35 : AOI22_X1 port map( A1 => N85, A2 => n84_port, B1 => N53, B2 => n12, ZN
                           => n30_port);
   U36 : NAND2_X1 port map( A1 => n79_port, A2 => n80_port, ZN => OUTPUT(0));
   U37 : AOI22_X1 port map( A1 => N18, A2 => n4, B1 => A(0), B2 => n1, ZN => 
                           n79_port);
   U38 : AOI22_X1 port map( A1 => N82, A2 => n82_port, B1 => N50, B2 => n10, ZN
                           => n80_port);
   U39 : AOI22_X1 port map( A1 => N25, A2 => n6, B1 => A(7), B2 => n3, ZN => 
                           n21_port);
   U40 : AOI22_X1 port map( A1 => N24, A2 => n6, B1 => A(6), B2 => n3, ZN => 
                           n23_port);
   U41 : AOI22_X1 port map( A1 => N30, A2 => n4, B1 => A(12), B2 => n1, ZN => 
                           n73_port);
   U42 : AOI22_X1 port map( A1 => N32, A2 => n4, B1 => A(14), B2 => n1, ZN => 
                           n69_port);
   U43 : AOI22_X1 port map( A1 => N35, A2 => n4, B1 => A(17), B2 => n1, ZN => 
                           n63_port);
   U44 : AOI22_X1 port map( A1 => N31, A2 => n4, B1 => A(13), B2 => n1, ZN => 
                           n71_port);
   U45 : AOI22_X1 port map( A1 => N33, A2 => n4, B1 => A(15), B2 => n1, ZN => 
                           n67_port);
   U46 : AOI22_X1 port map( A1 => N34, A2 => n4, B1 => A(16), B2 => n1, ZN => 
                           n65_port);
   U47 : AOI22_X1 port map( A1 => N45, A2 => n5, B1 => A(27), B2 => n2, ZN => 
                           n41_port);
   U48 : AOI22_X1 port map( A1 => N44, A2 => n5, B1 => A(26), B2 => n2, ZN => 
                           n43_port);
   U49 : AOI22_X1 port map( A1 => N49, A2 => n6, B1 => A(31), B2 => n3, ZN => 
                           n31_port);
   U50 : AOI22_X1 port map( A1 => N46, A2 => n5, B1 => A(28), B2 => n2, ZN => 
                           n39_port);
   U51 : AOI22_X1 port map( A1 => N36, A2 => n4, B1 => A(18), B2 => n1, ZN => 
                           n61_port);
   U52 : AOI22_X1 port map( A1 => N113, A2 => n84_port, B1 => N81, B2 => n12, 
                           ZN => n32_port);
   U53 : AOI22_X1 port map( A1 => N47, A2 => n5, B1 => A(29), B2 => n2, ZN => 
                           n37_port);
   U54 : BUF_X1 port map( A => n15, Z => n82_port);
   U55 : BUF_X1 port map( A => n15, Z => n83_port);
   U56 : BUF_X1 port map( A => n16, Z => n10);
   U57 : BUF_X1 port map( A => n16, Z => n11);
   U58 : AOI22_X1 port map( A1 => N37, A2 => n4, B1 => A(19), B2 => n1, ZN => 
                           n59_port);
   U59 : BUF_X1 port map( A => n17, Z => n4);
   U60 : BUF_X1 port map( A => n17, Z => n5);
   U61 : BUF_X1 port map( A => n18_port, Z => n1);
   U62 : BUF_X1 port map( A => n18_port, Z => n2);
   U63 : AOI22_X1 port map( A1 => N48, A2 => n5, B1 => A(30), B2 => n2, ZN => 
                           n33_port);
   U64 : BUF_X1 port map( A => n15, Z => n84_port);
   U65 : BUF_X1 port map( A => n16, Z => n12);
   U66 : AOI22_X1 port map( A1 => N109, A2 => n83_port, B1 => N77, B2 => n11, 
                           ZN => n42_port);
   U67 : BUF_X1 port map( A => n17, Z => n6);
   U68 : AOI22_X1 port map( A1 => N26, A2 => n6, B1 => A(8), B2 => n3, ZN => 
                           n19_port);
   U69 : AOI22_X1 port map( A1 => N27, A2 => n6, B1 => A(9), B2 => n3, ZN => 
                           n13);
   U70 : BUF_X1 port map( A => n18_port, Z => n3);
   U71 : AOI22_X1 port map( A1 => N28, A2 => n4, B1 => A(10), B2 => n1, ZN => 
                           n77_port);
   U72 : AOI22_X1 port map( A1 => N42, A2 => n5, B1 => A(24), B2 => n2, ZN => 
                           n47_port);
   U73 : AOI22_X1 port map( A1 => N43, A2 => n5, B1 => A(25), B2 => n2, ZN => 
                           n45_port);
   U74 : AOI22_X1 port map( A1 => N29, A2 => n4, B1 => A(11), B2 => n1, ZN => 
                           n75_port);
   U75 : INV_X1 port map( A => n81_port, ZN => n86_port);
   U76 : NAND2_X1 port map( A1 => n35_port, A2 => n36_port, ZN => OUTPUT(2));
   U77 : AOI22_X1 port map( A1 => N84, A2 => n83_port, B1 => N52, B2 => n11, ZN
                           => n36_port);
   U78 : AOI22_X1 port map( A1 => N39, A2 => n5, B1 => A(21), B2 => n2, ZN => 
                           n53_port);
   U79 : AOI22_X1 port map( A1 => N38, A2 => n5, B1 => A(20), B2 => n2, ZN => 
                           n55_port);
   U80 : AOI22_X1 port map( A1 => N40, A2 => n5, B1 => A(22), B2 => n2, ZN => 
                           n51_port);
   U81 : AOI22_X1 port map( A1 => N41, A2 => n5, B1 => A(23), B2 => n2, ZN => 
                           n49_port);
   U82 : NOR3_X1 port map( A1 => sel(4), A2 => sel(1), A3 => n81_port, ZN => 
                           n17);
   U83 : INV_X1 port map( A => sel(0), ZN => n87_port);
   U84 : OAI21_X1 port map( B1 => sel(4), B2 => n88_port, A => n86_port, ZN => 
                           n18_port);
   U85 : INV_X1 port map( A => sel(1), ZN => n88_port);
   U86 : AND3_X1 port map( A1 => sel(4), A2 => n86_port, A3 => sel(1), ZN => 
                           n15);
   U87 : AND3_X1 port map( A1 => n86_port, A2 => n88_port, A3 => sel(4), ZN => 
                           n16);
   U88 : NAND2_X1 port map( A1 => n39_port, A2 => n40_port, ZN => OUTPUT(28));
   U89 : NAND2_X1 port map( A1 => n37_port, A2 => n38_port, ZN => OUTPUT(29));
   U90 : NAND2_X1 port map( A1 => n33_port, A2 => n34_port, ZN => OUTPUT(30));
   U91 : NAND2_X1 port map( A1 => n55_port, A2 => n56_port, ZN => OUTPUT(20));
   U92 : NAND2_X1 port map( A1 => n53_port, A2 => n54_port, ZN => OUTPUT(21));
   U93 : NAND2_X1 port map( A1 => n51_port, A2 => n52_port, ZN => OUTPUT(22));
   U94 : NAND2_X1 port map( A1 => n49_port, A2 => n50_port, ZN => OUTPUT(23));
   U95 : NAND2_X1 port map( A1 => n47_port, A2 => n48_port, ZN => OUTPUT(24));
   U96 : NAND2_X1 port map( A1 => n45_port, A2 => n46_port, ZN => OUTPUT(25));
   U97 : NAND2_X1 port map( A1 => n43_port, A2 => n44_port, ZN => OUTPUT(26));
   U98 : NAND2_X1 port map( A1 => n41_port, A2 => n42_port, ZN => OUTPUT(27));
   U99 : NAND2_X1 port map( A1 => n63_port, A2 => n64_port, ZN => OUTPUT(17));
   U100 : NAND2_X1 port map( A1 => n61_port, A2 => n62_port, ZN => OUTPUT(18));
   U101 : NAND2_X1 port map( A1 => n59_port, A2 => n60_port, ZN => OUTPUT(19));
   U102 : NAND2_X1 port map( A1 => n65_port, A2 => n66_port, ZN => OUTPUT(16));
   U103 : NAND2_X1 port map( A1 => n73_port, A2 => n74_port, ZN => OUTPUT(12));
   U104 : NAND2_X1 port map( A1 => n71_port, A2 => n72_port, ZN => OUTPUT(13));
   U105 : NAND2_X1 port map( A1 => n69_port, A2 => n70_port, ZN => OUTPUT(14));
   U106 : NAND2_X1 port map( A1 => n67_port, A2 => n68_port, ZN => OUTPUT(15));
   U107 : NAND2_X1 port map( A1 => n31_port, A2 => n32_port, ZN => OUTPUT(31));
   U108 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => OUTPUT(9));
   U109 : NAND2_X1 port map( A1 => n19_port, A2 => n20_port, ZN => OUTPUT(8));
   U111 : NAND2_X1 port map( A1 => n77_port, A2 => n78_port, ZN => OUTPUT(10));
   U112 : NAND2_X1 port map( A1 => n75_port, A2 => n76_port, ZN => OUTPUT(11));
   U113 : NAND2_X1 port map( A1 => n21_port, A2 => n22_port, ZN => OUTPUT(7));
   U114 : NAND2_X1 port map( A1 => n23_port, A2 => n24_port, ZN => OUTPUT(6));
   U115 : NAND2_X1 port map( A1 => n27_port, A2 => n28_port, ZN => OUTPUT(4));
   U116 : NAND2_X1 port map( A1 => n25_port, A2 => n26_port, ZN => OUTPUT(5));
   U117 : AOI22_X1 port map( A1 => N20, A2 => n5, B1 => A(2), B2 => n2, ZN => 
                           n35_port);
   U118 : AOI22_X1 port map( A1 => N23, A2 => n6, B1 => A(5), B2 => n3, ZN => 
                           n25_port);
   U119 : AOI22_X1 port map( A1 => N22, A2 => n6, B1 => A(4), B2 => n3, ZN => 
                           n27_port);
   U120 : AOI22_X1 port map( A1 => N19, A2 => n4, B1 => A(1), B2 => n1, ZN => 
                           n57_port);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity logic_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic_vector 
         (0 to 4);  O : out std_logic_vector (31 downto 0));

end logic_N32;

architecture SYN_Behavioral of logic_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n69, n135, n136, n137, n138, 
      n139, n140, n141, n142 : std_logic;

begin
   
   U2 : INV_X1 port map( A => SEL(2), ZN => n142);
   U3 : AOI22_X1 port map( A1 => n8, A2 => n16, B1 => A(0), B2 => n2, ZN => 
                           n132);
   U4 : AOI22_X1 port map( A1 => n9, A2 => n41, B1 => A(3), B2 => n4, ZN => n82
                           );
   U5 : AOI21_X1 port map( B1 => n10, B2 => n11, A => n5, ZN => n133);
   U6 : AOI21_X1 port map( B1 => n10, B2 => n12, A => n5, ZN => n111);
   U7 : AOI21_X1 port map( B1 => n9, B2 => n13, A => n6, ZN => n89);
   U8 : AOI21_X1 port map( B1 => n8, B2 => n14, A => n7, ZN => n83);
   U9 : INV_X1 port map( A => A(3), ZN => n41);
   U10 : INV_X1 port map( A => A(0), ZN => n16);
   U11 : INV_X1 port map( A => n1, ZN => n10);
   U12 : BUF_X1 port map( A => n70, Z => n5);
   U13 : BUF_X1 port map( A => n70, Z => n6);
   U14 : OAI22_X1 port map( A1 => n116, A2 => n55, B1 => n117, B2 => n24, ZN =>
                           O(17));
   U15 : AOI21_X1 port map( B1 => n10, B2 => n55, A => n5, ZN => n117);
   U16 : AOI22_X1 port map( A1 => n9, A2 => n24, B1 => A(17), B2 => n2, ZN => 
                           n116);
   U17 : INV_X1 port map( A => B(17), ZN => n55);
   U18 : OAI22_X1 port map( A1 => n106, A2 => n59, B1 => n107, B2 => n29, ZN =>
                           O(21));
   U19 : AOI21_X1 port map( B1 => n10, B2 => n59, A => n6, ZN => n107);
   U20 : AOI22_X1 port map( A1 => n9, A2 => n29, B1 => A(21), B2 => n3, ZN => 
                           n106);
   U21 : INV_X1 port map( A => B(21), ZN => n59);
   U22 : OAI22_X1 port map( A1 => n80, A2 => n15, B1 => n81, B2 => n42, ZN => 
                           O(4));
   U23 : AOI21_X1 port map( B1 => n9, B2 => n15, A => n7, ZN => n81);
   U24 : OAI22_X1 port map( A1 => n78, A2 => n137, B1 => n79, B2 => n43, ZN => 
                           O(5));
   U25 : AOI21_X1 port map( B1 => n8, B2 => n137, A => n7, ZN => n79);
   U26 : INV_X1 port map( A => B(5), ZN => n137);
   U27 : OAI22_X1 port map( A1 => n74, A2 => n139, B1 => n75, B2 => n45, ZN => 
                           O(7));
   U28 : AOI21_X1 port map( B1 => n8, B2 => n139, A => n7, ZN => n75);
   U29 : AOI22_X1 port map( A1 => n8, A2 => n45, B1 => A(7), B2 => n4, ZN => 
                           n74);
   U30 : INV_X1 port map( A => B(7), ZN => n139);
   U31 : OAI22_X1 port map( A1 => n76, A2 => n138, B1 => n77, B2 => n44, ZN => 
                           O(6));
   U32 : AOI21_X1 port map( B1 => n8, B2 => n138, A => n7, ZN => n77);
   U33 : AOI22_X1 port map( A1 => n8, A2 => n44, B1 => A(6), B2 => n4, ZN => 
                           n76);
   U34 : INV_X1 port map( A => B(6), ZN => n138);
   U35 : OAI22_X1 port map( A1 => n67, A2 => n141, B1 => n68, B2 => n47, ZN => 
                           O(9));
   U36 : AOI21_X1 port map( B1 => n9, B2 => n141, A => n7, ZN => n68);
   U37 : AOI22_X1 port map( A1 => n8, A2 => n47, B1 => n4, B2 => A(9), ZN => 
                           n67);
   U38 : INV_X1 port map( A => B(9), ZN => n141);
   U39 : OAI22_X1 port map( A1 => n72, A2 => n140, B1 => n73, B2 => n46, ZN => 
                           O(8));
   U40 : AOI21_X1 port map( B1 => n8, B2 => n140, A => n7, ZN => n73);
   U41 : AOI22_X1 port map( A1 => n8, A2 => n46, B1 => A(8), B2 => n4, ZN => 
                           n72);
   U42 : INV_X1 port map( A => B(8), ZN => n140);
   U43 : OAI22_X1 port map( A1 => n130, A2 => n48, B1 => n131, B2 => n17, ZN =>
                           O(10));
   U44 : AOI21_X1 port map( B1 => n8, B2 => n48, A => n5, ZN => n131);
   U45 : AOI22_X1 port map( A1 => n8, A2 => n17, B1 => A(10), B2 => n2, ZN => 
                           n130);
   U46 : INV_X1 port map( A => B(10), ZN => n48);
   U47 : OAI22_X1 port map( A1 => n128, A2 => n49, B1 => n129, B2 => n18, ZN =>
                           O(11));
   U48 : AOI21_X1 port map( B1 => n9, B2 => n49, A => n5, ZN => n129);
   U49 : AOI22_X1 port map( A1 => n8, A2 => n18, B1 => A(11), B2 => n2, ZN => 
                           n128);
   U50 : INV_X1 port map( A => B(11), ZN => n49);
   U51 : OAI22_X1 port map( A1 => n112, A2 => n57, B1 => n113, B2 => n26, ZN =>
                           O(19));
   U52 : AOI21_X1 port map( B1 => n10, B2 => n57, A => n5, ZN => n113);
   U53 : AOI22_X1 port map( A1 => n9, A2 => n26, B1 => A(19), B2 => n2, ZN => 
                           n112);
   U54 : INV_X1 port map( A => B(19), ZN => n57);
   U55 : OAI22_X1 port map( A1 => n108, A2 => n58, B1 => n109, B2 => n28, ZN =>
                           O(20));
   U56 : AOI21_X1 port map( B1 => n10, B2 => n58, A => n6, ZN => n109);
   U57 : AOI22_X1 port map( A1 => n9, A2 => n28, B1 => A(20), B2 => n3, ZN => 
                           n108);
   U58 : INV_X1 port map( A => B(20), ZN => n58);
   U59 : BUF_X1 port map( A => n71, Z => n2);
   U60 : BUF_X1 port map( A => n71, Z => n3);
   U61 : OAI22_X1 port map( A1 => n86, A2 => n135, B1 => n87, B2 => n39, ZN => 
                           O(30));
   U62 : AOI21_X1 port map( B1 => n8, B2 => n135, A => n6, ZN => n87);
   U63 : AOI22_X1 port map( A1 => n9, A2 => n39, B1 => A(30), B2 => n3, ZN => 
                           n86);
   U64 : INV_X1 port map( A => B(30), ZN => n135);
   U65 : INV_X1 port map( A => A(7), ZN => n45);
   U66 : OAI22_X1 port map( A1 => n102, A2 => n61, B1 => n103, B2 => n31, ZN =>
                           O(23));
   U67 : AOI21_X1 port map( B1 => n10, B2 => n61, A => n6, ZN => n103);
   U68 : AOI22_X1 port map( A1 => n9, A2 => n31, B1 => A(23), B2 => n3, ZN => 
                           n102);
   U69 : INV_X1 port map( A => B(23), ZN => n61);
   U70 : OAI22_X1 port map( A1 => n126, A2 => n50, B1 => n127, B2 => n19, ZN =>
                           O(12));
   U71 : AOI21_X1 port map( B1 => n10, B2 => n50, A => n5, ZN => n127);
   U72 : AOI22_X1 port map( A1 => n8, A2 => n19, B1 => A(12), B2 => n2, ZN => 
                           n126);
   U73 : INV_X1 port map( A => B(12), ZN => n50);
   U74 : OAI22_X1 port map( A1 => n122, A2 => n52, B1 => n123, B2 => n21, ZN =>
                           O(14));
   U75 : AOI21_X1 port map( B1 => n10, B2 => n52, A => n5, ZN => n123);
   U76 : AOI22_X1 port map( A1 => n8, A2 => n21, B1 => A(14), B2 => n2, ZN => 
                           n122);
   U77 : INV_X1 port map( A => B(14), ZN => n52);
   U78 : OAI22_X1 port map( A1 => n124, A2 => n51, B1 => n125, B2 => n20, ZN =>
                           O(13));
   U79 : AOI21_X1 port map( B1 => n8, B2 => n51, A => n5, ZN => n125);
   U80 : AOI22_X1 port map( A1 => n8, A2 => n20, B1 => A(13), B2 => n2, ZN => 
                           n124);
   U81 : INV_X1 port map( A => B(13), ZN => n51);
   U82 : OAI22_X1 port map( A1 => n120, A2 => n53, B1 => n121, B2 => n22, ZN =>
                           O(15));
   U83 : AOI21_X1 port map( B1 => n10, B2 => n53, A => n5, ZN => n121);
   U84 : AOI22_X1 port map( A1 => n8, A2 => n22, B1 => A(15), B2 => n2, ZN => 
                           n120);
   U85 : INV_X1 port map( A => B(15), ZN => n53);
   U86 : OAI22_X1 port map( A1 => n118, A2 => n54, B1 => n119, B2 => n23, ZN =>
                           O(16));
   U87 : AOI21_X1 port map( B1 => n10, B2 => n54, A => n5, ZN => n119);
   U88 : AOI22_X1 port map( A1 => n8, A2 => n23, B1 => A(16), B2 => n2, ZN => 
                           n118);
   U89 : INV_X1 port map( A => B(16), ZN => n54);
   U90 : OAI22_X1 port map( A1 => n94, A2 => n65, B1 => n95, B2 => n35, ZN => 
                           O(27));
   U91 : AOI21_X1 port map( B1 => n10, B2 => n65, A => n6, ZN => n95);
   U92 : AOI22_X1 port map( A1 => n10, A2 => n35, B1 => A(27), B2 => n3, ZN => 
                           n94);
   U93 : INV_X1 port map( A => B(27), ZN => n65);
   U94 : OAI22_X1 port map( A1 => n96, A2 => n64, B1 => n97, B2 => n34, ZN => 
                           O(26));
   U95 : AOI21_X1 port map( B1 => n8, B2 => n64, A => n6, ZN => n97);
   U96 : AOI22_X1 port map( A1 => n9, A2 => n34, B1 => A(26), B2 => n3, ZN => 
                           n96);
   U97 : INV_X1 port map( A => B(26), ZN => n64);
   U98 : OAI22_X1 port map( A1 => n84, A2 => n136, B1 => n85, B2 => n40, ZN => 
                           O(31));
   U99 : AOI21_X1 port map( B1 => n9, B2 => n136, A => n7, ZN => n85);
   U100 : AOI22_X1 port map( A1 => n8, A2 => n40, B1 => A(31), B2 => n4, ZN => 
                           n84);
   U101 : INV_X1 port map( A => B(31), ZN => n136);
   U102 : OAI22_X1 port map( A1 => n92, A2 => n66, B1 => n93, B2 => n36, ZN => 
                           O(28));
   U103 : AOI21_X1 port map( B1 => n10, B2 => n66, A => n6, ZN => n93);
   U104 : AOI22_X1 port map( A1 => n9, A2 => n36, B1 => A(28), B2 => n3, ZN => 
                           n92);
   U105 : INV_X1 port map( A => B(28), ZN => n66);
   U106 : OAI22_X1 port map( A1 => n114, A2 => n56, B1 => n115, B2 => n25, ZN 
                           => O(18));
   U107 : AOI21_X1 port map( B1 => n10, B2 => n56, A => n5, ZN => n115);
   U108 : AOI22_X1 port map( A1 => n9, A2 => n25, B1 => A(18), B2 => n2, ZN => 
                           n114);
   U109 : INV_X1 port map( A => B(18), ZN => n56);
   U110 : OAI22_X1 port map( A1 => n90, A2 => n69, B1 => n91, B2 => n37, ZN => 
                           O(29));
   U111 : AOI21_X1 port map( B1 => n8, B2 => n69, A => n6, ZN => n91);
   U112 : AOI22_X1 port map( A1 => n8, A2 => n37, B1 => A(29), B2 => n3, ZN => 
                           n90);
   U113 : INV_X1 port map( A => B(29), ZN => n69);
   U114 : INV_X1 port map( A => A(6), ZN => n44);
   U115 : OAI22_X1 port map( A1 => n104, A2 => n60, B1 => n105, B2 => n30, ZN 
                           => O(22));
   U116 : AOI21_X1 port map( B1 => n10, B2 => n60, A => n6, ZN => n105);
   U117 : AOI22_X1 port map( A1 => n9, A2 => n30, B1 => A(22), B2 => n3, ZN => 
                           n104);
   U118 : INV_X1 port map( A => B(22), ZN => n60);
   U119 : OAI22_X1 port map( A1 => n100, A2 => n62, B1 => n101, B2 => n32, ZN 
                           => O(24));
   U120 : AOI21_X1 port map( B1 => n10, B2 => n62, A => n6, ZN => n101);
   U121 : AOI22_X1 port map( A1 => n9, A2 => n32, B1 => A(24), B2 => n3, ZN => 
                           n100);
   U122 : INV_X1 port map( A => B(24), ZN => n62);
   U123 : OAI22_X1 port map( A1 => n98, A2 => n63, B1 => n99, B2 => n33, ZN => 
                           O(25));
   U124 : AOI21_X1 port map( B1 => n9, B2 => n63, A => n6, ZN => n99);
   U125 : AOI22_X1 port map( A1 => n9, A2 => n33, B1 => A(25), B2 => n3, ZN => 
                           n98);
   U126 : INV_X1 port map( A => B(25), ZN => n63);
   U127 : INV_X1 port map( A => A(12), ZN => n19);
   U128 : INV_X1 port map( A => A(14), ZN => n21);
   U129 : BUF_X1 port map( A => n70, Z => n7);
   U130 : INV_X1 port map( A => A(17), ZN => n24);
   U131 : INV_X1 port map( A => A(21), ZN => n29);
   U132 : INV_X1 port map( A => A(13), ZN => n20);
   U133 : INV_X1 port map( A => A(15), ZN => n22);
   U134 : INV_X1 port map( A => A(16), ZN => n23);
   U135 : INV_X1 port map( A => A(27), ZN => n35);
   U136 : INV_X1 port map( A => A(26), ZN => n34);
   U137 : INV_X1 port map( A => A(31), ZN => n40);
   U138 : BUF_X1 port map( A => n71, Z => n4);
   U139 : INV_X1 port map( A => A(28), ZN => n36);
   U140 : INV_X1 port map( A => A(18), ZN => n25);
   U141 : INV_X1 port map( A => A(29), ZN => n37);
   U142 : INV_X1 port map( A => A(19), ZN => n26);
   U143 : INV_X1 port map( A => A(20), ZN => n28);
   U144 : INV_X1 port map( A => A(30), ZN => n39);
   U145 : INV_X1 port map( A => A(9), ZN => n47);
   U146 : INV_X1 port map( A => A(8), ZN => n46);
   U147 : INV_X1 port map( A => A(10), ZN => n17);
   U148 : INV_X1 port map( A => A(11), ZN => n18);
   U149 : INV_X1 port map( A => A(23), ZN => n31);
   U150 : INV_X1 port map( A => A(22), ZN => n30);
   U151 : INV_X1 port map( A => A(24), ZN => n32);
   U152 : INV_X1 port map( A => A(25), ZN => n33);
   U153 : OAI22_X1 port map( A1 => n132, A2 => n11, B1 => n133, B2 => n16, ZN 
                           => O(0));
   U154 : NOR2_X1 port map( A1 => n1, A2 => SEL(4), ZN => n70);
   U155 : AND3_X1 port map( A1 => SEL(3), A2 => SEL(4), A3 => n134, ZN => n71);
   U156 : NOR3_X1 port map( A1 => SEL(2), A2 => SEL(0), A3 => SEL(1), ZN => 
                           n134);
   U157 : OR4_X1 port map( A1 => n142, A2 => SEL(3), A3 => SEL(1), A4 => SEL(0)
                           , ZN => n1);
   U158 : OAI22_X1 port map( A1 => n110, A2 => n12, B1 => n111, B2 => n27, ZN 
                           => O(1));
   U159 : OAI22_X1 port map( A1 => n88, A2 => n13, B1 => n89, B2 => n38, ZN => 
                           O(2));
   U160 : OAI22_X1 port map( A1 => n82, A2 => n14, B1 => n83, B2 => n41, ZN => 
                           O(3));
   U161 : AOI22_X1 port map( A1 => n8, A2 => n38, B1 => A(2), B2 => n3, ZN => 
                           n88);
   U162 : INV_X1 port map( A => A(2), ZN => n38);
   U163 : AOI22_X1 port map( A1 => n9, A2 => n43, B1 => A(5), B2 => n4, ZN => 
                           n78);
   U164 : INV_X1 port map( A => A(5), ZN => n43);
   U165 : AOI22_X1 port map( A1 => n9, A2 => n42, B1 => A(4), B2 => n4, ZN => 
                           n80);
   U166 : INV_X1 port map( A => A(4), ZN => n42);
   U167 : AOI22_X1 port map( A1 => n9, A2 => n27, B1 => A(1), B2 => n2, ZN => 
                           n110);
   U168 : INV_X1 port map( A => A(1), ZN => n27);
   U169 : INV_X1 port map( A => n1, ZN => n8);
   U170 : INV_X1 port map( A => n1, ZN => n9);
   U171 : INV_X1 port map( A => B(0), ZN => n11);
   U172 : INV_X1 port map( A => B(1), ZN => n12);
   U173 : INV_X1 port map( A => B(2), ZN => n13);
   U174 : INV_X1 port map( A => B(3), ZN => n14);
   U175 : INV_X1 port map( A => B(4), ZN => n15);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity add_wrapper_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic_vector 
         (0 to 4);  O : out std_logic_vector (31 downto 0));

end add_wrapper_N32;

architecture SYN_Behavioral of add_wrapper_N32 is

   component P4_ADDER_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component add_sub_N32
      port( A : in std_logic_vector (31 downto 0);  SEL : in std_logic_vector 
            (0 to 4);  O : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, outp_31_port, outp_30_port, outp_29_port, outp_28_port
      , outp_27_port, outp_26_port, outp_25_port, outp_24_port, outp_23_port, 
      outp_22_port, outp_21_port, outp_20_port, outp_19_port, outp_18_port, 
      outp_17_port, outp_16_port, outp_15_port, outp_14_port, outp_13_port, 
      outp_12_port, outp_11_port, outp_10_port, outp_9_port, outp_8_port, 
      outp_7_port, outp_6_port, outp_5_port, outp_4_port, outp_3_port, 
      outp_2_port, outp_1_port, outp_0_port, n_1144 : std_logic;

begin
   
   X_Logic0_port <= '0';
   sign : add_sub_N32 port map( A(31) => B(31), A(30) => B(30), A(29) => B(29),
                           A(28) => B(28), A(27) => B(27), A(26) => B(26), 
                           A(25) => B(25), A(24) => B(24), A(23) => B(23), 
                           A(22) => B(22), A(21) => B(21), A(20) => B(20), 
                           A(19) => B(19), A(18) => B(18), A(17) => B(17), 
                           A(16) => B(16), A(15) => B(15), A(14) => B(14), 
                           A(13) => B(13), A(12) => B(12), A(11) => B(11), 
                           A(10) => B(10), A(9) => B(9), A(8) => B(8), A(7) => 
                           B(7), A(6) => B(6), A(5) => B(5), A(4) => B(4), A(3)
                           => B(3), A(2) => B(2), A(1) => B(1), A(0) => B(0), 
                           SEL(0) => SEL(0), SEL(1) => SEL(1), SEL(2) => SEL(2)
                           , SEL(3) => SEL(3), SEL(4) => SEL(4), O(31) => 
                           outp_31_port, O(30) => outp_30_port, O(29) => 
                           outp_29_port, O(28) => outp_28_port, O(27) => 
                           outp_27_port, O(26) => outp_26_port, O(25) => 
                           outp_25_port, O(24) => outp_24_port, O(23) => 
                           outp_23_port, O(22) => outp_22_port, O(21) => 
                           outp_21_port, O(20) => outp_20_port, O(19) => 
                           outp_19_port, O(18) => outp_18_port, O(17) => 
                           outp_17_port, O(16) => outp_16_port, O(15) => 
                           outp_15_port, O(14) => outp_14_port, O(13) => 
                           outp_13_port, O(12) => outp_12_port, O(11) => 
                           outp_11_port, O(10) => outp_10_port, O(9) => 
                           outp_9_port, O(8) => outp_8_port, O(7) => 
                           outp_7_port, O(6) => outp_6_port, O(5) => 
                           outp_5_port, O(4) => outp_4_port, O(3) => 
                           outp_3_port, O(2) => outp_2_port, O(1) => 
                           outp_1_port, O(0) => outp_0_port);
   adder : P4_ADDER_NBIT32 port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => outp_31_port, B(30) => 
                           outp_30_port, B(29) => outp_29_port, B(28) => 
                           outp_28_port, B(27) => outp_27_port, B(26) => 
                           outp_26_port, B(25) => outp_25_port, B(24) => 
                           outp_24_port, B(23) => outp_23_port, B(22) => 
                           outp_22_port, B(21) => outp_21_port, B(20) => 
                           outp_20_port, B(19) => outp_19_port, B(18) => 
                           outp_18_port, B(17) => outp_17_port, B(16) => 
                           outp_16_port, B(15) => outp_15_port, B(14) => 
                           outp_14_port, B(13) => outp_13_port, B(12) => 
                           outp_12_port, B(11) => outp_11_port, B(10) => 
                           outp_10_port, B(9) => outp_9_port, B(8) => 
                           outp_8_port, B(7) => outp_7_port, B(6) => 
                           outp_6_port, B(5) => outp_5_port, B(4) => 
                           outp_4_port, B(3) => outp_3_port, B(2) => 
                           outp_2_port, B(1) => outp_1_port, B(0) => 
                           outp_0_port, Cin => X_Logic0_port, S(31) => O(31), 
                           S(30) => O(30), S(29) => O(29), S(28) => O(28), 
                           S(27) => O(27), S(26) => O(26), S(25) => O(25), 
                           S(24) => O(24), S(23) => O(23), S(22) => O(22), 
                           S(21) => O(21), S(20) => O(20), S(19) => O(19), 
                           S(18) => O(18), S(17) => O(17), S(16) => O(16), 
                           S(15) => O(15), S(14) => O(14), S(13) => O(13), 
                           S(12) => O(12), S(11) => O(11), S(10) => O(10), S(9)
                           => O(9), S(8) => O(8), S(7) => O(7), S(6) => O(6), 
                           S(5) => O(5), S(4) => O(4), S(3) => O(3), S(2) => 
                           O(2), S(1) => O(1), S(0) => O(0), Cout => n_1144);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FWD_CAM_0 is

   port( RST : in std_logic;  DATA_IN_1, DATA_IN_2, DATA_IN_3 : in 
         std_logic_vector (5 downto 0);  MATCH_1, MATCH_2, MATCH_3 : out 
         std_logic);

end FWD_CAM_0;

architecture SYN_Behavioral of FWD_CAM_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net35857, net28092, net28091, net28089, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => n29, A2 => RST, ZN => MATCH_2);
   U4 : AND2_X1 port map( A1 => DATA_IN_1(3), A2 => DATA_IN_1(4), ZN => n1);
   U5 : AND2_X1 port map( A1 => DATA_IN_2(3), A2 => DATA_IN_2(4), ZN => n2);
   U6 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n6, B2 => n8, ZN => n3);
   U7 : OAI21_X1 port map( B1 => n3, B2 => DATA_IN_3(5), A => net28091, ZN => 
                           net28089);
   U8 : CLKBUF_X1 port map( A => DATA_IN_3(3), Z => n8);
   U9 : AND2_X1 port map( A1 => DATA_IN_3(4), A2 => n8, ZN => net35857);
   U10 : OAI211_X1 port map( C1 => DATA_IN_3(0), C2 => DATA_IN_3(4), A => 
                           DATA_IN_3(1), B => DATA_IN_3(2), ZN => n6);
   U11 : AND2_X1 port map( A1 => DATA_IN_3(4), A2 => DATA_IN_3(2), ZN => n4);
   U12 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n5);
   U13 : NAND2_X1 port map( A1 => n7, A2 => DATA_IN_3(1), ZN => n10);
   U14 : INV_X1 port map( A => DATA_IN_3(3), ZN => n7);
   U15 : OR2_X1 port map( A1 => DATA_IN_3(0), A2 => DATA_IN_3(1), ZN => n9);
   U16 : XOR2_X1 port map( A => DATA_IN_3(1), B => DATA_IN_3(2), Z => net28092)
                           ;
   U17 : OR2_X1 port map( A1 => DATA_IN_1(1), A2 => DATA_IN_1(0), ZN => n16);
   U18 : AND2_X1 port map( A1 => net28089, A2 => RST, ZN => MATCH_3);
   U19 : NAND2_X1 port map( A1 => net28092, A2 => net35857, ZN => net28091);
   U20 : NAND2_X1 port map( A1 => n26, A2 => n2, ZN => n27);
   U21 : NAND2_X1 port map( A1 => DATA_IN_2(1), A2 => n12, ZN => n13);
   U22 : NAND2_X1 port map( A1 => n11, A2 => DATA_IN_2(2), ZN => n14);
   U23 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n26);
   U24 : INV_X1 port map( A => DATA_IN_2(1), ZN => n11);
   U25 : INV_X1 port map( A => DATA_IN_2(2), ZN => n12);
   U26 : AND2_X1 port map( A1 => DATA_IN_1(4), A2 => DATA_IN_1(2), ZN => n33);
   U27 : NAND2_X1 port map( A1 => n30, A2 => DATA_IN_1(1), ZN => n17);
   U28 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n32);
   U29 : INV_X1 port map( A => DATA_IN_1(1), ZN => n15);
   U30 : NAND2_X1 port map( A1 => n34, A2 => n1, ZN => n35);
   U31 : AND2_X1 port map( A1 => DATA_IN_2(4), A2 => DATA_IN_2(2), ZN => n25);
   U32 : NAND2_X1 port map( A1 => DATA_IN_1(1), A2 => n18, ZN => n19);
   U33 : NAND2_X1 port map( A1 => n15, A2 => DATA_IN_1(2), ZN => n20);
   U34 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => n34);
   U35 : INV_X1 port map( A => DATA_IN_1(2), ZN => n18);
   U36 : INV_X1 port map( A => DATA_IN_2(0), ZN => n22);
   U37 : INV_X1 port map( A => DATA_IN_2(3), ZN => n21);
   U38 : MUX2_X1 port map( A => n22, B => n21, S => DATA_IN_2(1), Z => n24);
   U39 : OAI211_X1 port map( C1 => DATA_IN_2(0), C2 => DATA_IN_2(4), A => 
                           DATA_IN_2(1), B => DATA_IN_2(2), ZN => n23);
   U40 : AOI22_X1 port map( A1 => n24, A2 => n25, B1 => n23, B2 => DATA_IN_2(3)
                           , ZN => n28);
   U41 : OAI21_X1 port map( B1 => n28, B2 => DATA_IN_2(5), A => n27, ZN => n29)
                           ;
   U42 : INV_X1 port map( A => DATA_IN_1(3), ZN => n30);
   U43 : OAI211_X1 port map( C1 => DATA_IN_1(0), C2 => DATA_IN_1(4), A => 
                           DATA_IN_1(1), B => DATA_IN_1(2), ZN => n31);
   U44 : AOI22_X1 port map( A1 => n33, A2 => n32, B1 => DATA_IN_1(3), B2 => n31
                           , ZN => n36);
   U45 : OAI21_X1 port map( B1 => n36, B2 => DATA_IN_1(5), A => n35, ZN => n37)
                           ;
   U46 : AND2_X1 port map( A1 => n37, A2 => RST, ZN => MATCH_1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity SNPS_CLOCK_GATE_HIGH_IF_ID is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic;  TE : in std_logic);

end SNPS_CLOCK_GATE_HIGH_IF_ID;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_IF_ID is

   component CLKGATETST_X1
      port( CK, E, SE : in std_logic;  GCK : out std_logic);
   end component;

begin
   
   latch : CLKGATETST_X1 port map( CK => CLK, E => EN, SE => TE, GCK => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MEM_WB is

   port( CLK, RST : in std_logic;  NPC_L_IN, ALU_IN, LMD_IN : in 
         std_logic_vector (31 downto 0);  RD_IN : in std_logic_vector (4 downto
         0);  OPCODE_IN : in std_logic_vector (5 downto 0);  NPC_L_OUT, ALU_OUT
         , LMD_OUT : out std_logic_vector (31 downto 0);  RD_OUT : out 
         std_logic_vector (4 downto 0);  OPCODE_OUT : out std_logic_vector (5 
         downto 0));

end MEM_WB;

architecture SYN_Behavioral of MEM_WB is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n3, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, 
      n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, 
      n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, 
      n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, 
      n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, 
      n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, 
      n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251 : 
      std_logic;

begin
   
   OPCODE_OUT_reg_5_inst : DFFR_X1 port map( D => OPCODE_IN(5), CK => CLK, RN 
                           => n12, Q => OPCODE_OUT(5), QN => n_1145);
   OPCODE_OUT_reg_4_inst : DFFR_X1 port map( D => OPCODE_IN(4), CK => CLK, RN 
                           => n12, Q => OPCODE_OUT(4), QN => n_1146);
   OPCODE_OUT_reg_3_inst : DFFR_X1 port map( D => OPCODE_IN(3), CK => CLK, RN 
                           => n12, Q => n_1147, QN => n7);
   OPCODE_OUT_reg_1_inst : DFFR_X1 port map( D => OPCODE_IN(1), CK => CLK, RN 
                           => n12, Q => n_1148, QN => n1);
   OPCODE_OUT_reg_0_inst : DFFR_X1 port map( D => OPCODE_IN(0), CK => CLK, RN 
                           => n12, Q => n_1149, QN => n3);
   ALU_OUT_reg_31_inst : DFFR_X1 port map( D => ALU_IN(31), CK => CLK, RN => 
                           n12, Q => ALU_OUT(31), QN => n_1150);
   ALU_OUT_reg_30_inst : DFFR_X1 port map( D => ALU_IN(30), CK => CLK, RN => 
                           n12, Q => ALU_OUT(30), QN => n_1151);
   ALU_OUT_reg_29_inst : DFFR_X1 port map( D => ALU_IN(29), CK => CLK, RN => 
                           n12, Q => ALU_OUT(29), QN => n_1152);
   ALU_OUT_reg_28_inst : DFFR_X1 port map( D => ALU_IN(28), CK => CLK, RN => 
                           n12, Q => ALU_OUT(28), QN => n_1153);
   ALU_OUT_reg_27_inst : DFFR_X1 port map( D => ALU_IN(27), CK => CLK, RN => 
                           n12, Q => ALU_OUT(27), QN => n_1154);
   ALU_OUT_reg_26_inst : DFFR_X1 port map( D => ALU_IN(26), CK => CLK, RN => 
                           n12, Q => ALU_OUT(26), QN => n_1155);
   ALU_OUT_reg_25_inst : DFFR_X1 port map( D => ALU_IN(25), CK => CLK, RN => 
                           n13, Q => ALU_OUT(25), QN => n_1156);
   ALU_OUT_reg_24_inst : DFFR_X1 port map( D => ALU_IN(24), CK => CLK, RN => 
                           n13, Q => ALU_OUT(24), QN => n_1157);
   ALU_OUT_reg_23_inst : DFFR_X1 port map( D => ALU_IN(23), CK => CLK, RN => 
                           n13, Q => ALU_OUT(23), QN => n_1158);
   ALU_OUT_reg_22_inst : DFFR_X1 port map( D => ALU_IN(22), CK => CLK, RN => 
                           n13, Q => ALU_OUT(22), QN => n_1159);
   ALU_OUT_reg_21_inst : DFFR_X1 port map( D => ALU_IN(21), CK => CLK, RN => 
                           n13, Q => ALU_OUT(21), QN => n_1160);
   ALU_OUT_reg_20_inst : DFFR_X1 port map( D => ALU_IN(20), CK => CLK, RN => 
                           n13, Q => ALU_OUT(20), QN => n_1161);
   ALU_OUT_reg_19_inst : DFFR_X1 port map( D => ALU_IN(19), CK => CLK, RN => 
                           n13, Q => ALU_OUT(19), QN => n_1162);
   ALU_OUT_reg_18_inst : DFFR_X1 port map( D => ALU_IN(18), CK => CLK, RN => 
                           n13, Q => ALU_OUT(18), QN => n_1163);
   ALU_OUT_reg_17_inst : DFFR_X1 port map( D => ALU_IN(17), CK => CLK, RN => 
                           n13, Q => ALU_OUT(17), QN => n_1164);
   ALU_OUT_reg_16_inst : DFFR_X1 port map( D => ALU_IN(16), CK => CLK, RN => 
                           n13, Q => ALU_OUT(16), QN => n_1165);
   ALU_OUT_reg_15_inst : DFFR_X1 port map( D => ALU_IN(15), CK => CLK, RN => 
                           n13, Q => ALU_OUT(15), QN => n_1166);
   ALU_OUT_reg_14_inst : DFFR_X1 port map( D => ALU_IN(14), CK => CLK, RN => 
                           n13, Q => ALU_OUT(14), QN => n_1167);
   ALU_OUT_reg_13_inst : DFFR_X1 port map( D => ALU_IN(13), CK => CLK, RN => 
                           n14, Q => ALU_OUT(13), QN => n_1168);
   ALU_OUT_reg_12_inst : DFFR_X1 port map( D => ALU_IN(12), CK => CLK, RN => 
                           n14, Q => ALU_OUT(12), QN => n_1169);
   ALU_OUT_reg_11_inst : DFFR_X1 port map( D => ALU_IN(11), CK => CLK, RN => 
                           n14, Q => ALU_OUT(11), QN => n_1170);
   ALU_OUT_reg_10_inst : DFFR_X1 port map( D => ALU_IN(10), CK => CLK, RN => 
                           n14, Q => ALU_OUT(10), QN => n_1171);
   ALU_OUT_reg_9_inst : DFFR_X1 port map( D => ALU_IN(9), CK => CLK, RN => n14,
                           Q => ALU_OUT(9), QN => n_1172);
   ALU_OUT_reg_8_inst : DFFR_X1 port map( D => ALU_IN(8), CK => CLK, RN => n14,
                           Q => ALU_OUT(8), QN => n_1173);
   ALU_OUT_reg_7_inst : DFFR_X1 port map( D => ALU_IN(7), CK => CLK, RN => n14,
                           Q => ALU_OUT(7), QN => n_1174);
   ALU_OUT_reg_6_inst : DFFR_X1 port map( D => ALU_IN(6), CK => CLK, RN => n14,
                           Q => ALU_OUT(6), QN => n_1175);
   ALU_OUT_reg_5_inst : DFFR_X1 port map( D => ALU_IN(5), CK => CLK, RN => n14,
                           Q => ALU_OUT(5), QN => n_1176);
   ALU_OUT_reg_4_inst : DFFR_X1 port map( D => ALU_IN(4), CK => CLK, RN => n14,
                           Q => ALU_OUT(4), QN => n_1177);
   ALU_OUT_reg_3_inst : DFFR_X1 port map( D => ALU_IN(3), CK => CLK, RN => n14,
                           Q => ALU_OUT(3), QN => n_1178);
   ALU_OUT_reg_2_inst : DFFR_X1 port map( D => ALU_IN(2), CK => CLK, RN => n14,
                           Q => ALU_OUT(2), QN => n_1179);
   ALU_OUT_reg_1_inst : DFFR_X1 port map( D => ALU_IN(1), CK => CLK, RN => n15,
                           Q => ALU_OUT(1), QN => n_1180);
   ALU_OUT_reg_0_inst : DFFR_X1 port map( D => ALU_IN(0), CK => CLK, RN => n15,
                           Q => ALU_OUT(0), QN => n_1181);
   LMD_OUT_reg_31_inst : DFFR_X1 port map( D => LMD_IN(31), CK => CLK, RN => 
                           n15, Q => LMD_OUT(31), QN => n_1182);
   LMD_OUT_reg_30_inst : DFFR_X1 port map( D => LMD_IN(30), CK => CLK, RN => 
                           n15, Q => LMD_OUT(30), QN => n_1183);
   LMD_OUT_reg_29_inst : DFFR_X1 port map( D => LMD_IN(29), CK => CLK, RN => 
                           n15, Q => LMD_OUT(29), QN => n_1184);
   LMD_OUT_reg_28_inst : DFFR_X1 port map( D => LMD_IN(28), CK => CLK, RN => 
                           n15, Q => LMD_OUT(28), QN => n_1185);
   LMD_OUT_reg_27_inst : DFFR_X1 port map( D => LMD_IN(27), CK => CLK, RN => 
                           n15, Q => LMD_OUT(27), QN => n_1186);
   LMD_OUT_reg_26_inst : DFFR_X1 port map( D => LMD_IN(26), CK => CLK, RN => 
                           n15, Q => LMD_OUT(26), QN => n_1187);
   LMD_OUT_reg_25_inst : DFFR_X1 port map( D => LMD_IN(25), CK => CLK, RN => 
                           n15, Q => LMD_OUT(25), QN => n_1188);
   LMD_OUT_reg_24_inst : DFFR_X1 port map( D => LMD_IN(24), CK => CLK, RN => 
                           n15, Q => LMD_OUT(24), QN => n_1189);
   LMD_OUT_reg_23_inst : DFFR_X1 port map( D => LMD_IN(23), CK => CLK, RN => 
                           n15, Q => LMD_OUT(23), QN => n_1190);
   LMD_OUT_reg_22_inst : DFFR_X1 port map( D => LMD_IN(22), CK => CLK, RN => 
                           n15, Q => LMD_OUT(22), QN => n_1191);
   LMD_OUT_reg_21_inst : DFFR_X1 port map( D => LMD_IN(21), CK => CLK, RN => 
                           n16, Q => LMD_OUT(21), QN => n_1192);
   LMD_OUT_reg_20_inst : DFFR_X1 port map( D => LMD_IN(20), CK => CLK, RN => 
                           n16, Q => LMD_OUT(20), QN => n_1193);
   LMD_OUT_reg_19_inst : DFFR_X1 port map( D => LMD_IN(19), CK => CLK, RN => 
                           n16, Q => LMD_OUT(19), QN => n_1194);
   LMD_OUT_reg_18_inst : DFFR_X1 port map( D => LMD_IN(18), CK => CLK, RN => 
                           n16, Q => LMD_OUT(18), QN => n_1195);
   LMD_OUT_reg_17_inst : DFFR_X1 port map( D => LMD_IN(17), CK => CLK, RN => 
                           n16, Q => LMD_OUT(17), QN => n_1196);
   LMD_OUT_reg_16_inst : DFFR_X1 port map( D => LMD_IN(16), CK => CLK, RN => 
                           n16, Q => LMD_OUT(16), QN => n_1197);
   LMD_OUT_reg_15_inst : DFFR_X1 port map( D => LMD_IN(15), CK => CLK, RN => 
                           n16, Q => LMD_OUT(15), QN => n_1198);
   LMD_OUT_reg_14_inst : DFFR_X1 port map( D => LMD_IN(14), CK => CLK, RN => 
                           n16, Q => LMD_OUT(14), QN => n_1199);
   LMD_OUT_reg_13_inst : DFFR_X1 port map( D => LMD_IN(13), CK => CLK, RN => 
                           n16, Q => LMD_OUT(13), QN => n_1200);
   LMD_OUT_reg_12_inst : DFFR_X1 port map( D => LMD_IN(12), CK => CLK, RN => 
                           n16, Q => LMD_OUT(12), QN => n_1201);
   LMD_OUT_reg_11_inst : DFFR_X1 port map( D => LMD_IN(11), CK => CLK, RN => 
                           n16, Q => LMD_OUT(11), QN => n_1202);
   LMD_OUT_reg_10_inst : DFFR_X1 port map( D => LMD_IN(10), CK => CLK, RN => 
                           n16, Q => LMD_OUT(10), QN => n_1203);
   LMD_OUT_reg_9_inst : DFFR_X1 port map( D => LMD_IN(9), CK => CLK, RN => n17,
                           Q => LMD_OUT(9), QN => n_1204);
   LMD_OUT_reg_8_inst : DFFR_X1 port map( D => LMD_IN(8), CK => CLK, RN => n17,
                           Q => LMD_OUT(8), QN => n_1205);
   LMD_OUT_reg_7_inst : DFFR_X1 port map( D => LMD_IN(7), CK => CLK, RN => n17,
                           Q => LMD_OUT(7), QN => n_1206);
   LMD_OUT_reg_6_inst : DFFR_X1 port map( D => LMD_IN(6), CK => CLK, RN => n17,
                           Q => LMD_OUT(6), QN => n_1207);
   LMD_OUT_reg_5_inst : DFFR_X1 port map( D => LMD_IN(5), CK => CLK, RN => n17,
                           Q => LMD_OUT(5), QN => n_1208);
   LMD_OUT_reg_4_inst : DFFR_X1 port map( D => LMD_IN(4), CK => CLK, RN => n17,
                           Q => LMD_OUT(4), QN => n_1209);
   LMD_OUT_reg_3_inst : DFFR_X1 port map( D => LMD_IN(3), CK => CLK, RN => n17,
                           Q => LMD_OUT(3), QN => n_1210);
   LMD_OUT_reg_2_inst : DFFR_X1 port map( D => LMD_IN(2), CK => CLK, RN => n17,
                           Q => LMD_OUT(2), QN => n_1211);
   LMD_OUT_reg_1_inst : DFFR_X1 port map( D => LMD_IN(1), CK => CLK, RN => n17,
                           Q => LMD_OUT(1), QN => n_1212);
   LMD_OUT_reg_0_inst : DFFR_X1 port map( D => LMD_IN(0), CK => CLK, RN => n17,
                           Q => LMD_OUT(0), QN => n_1213);
   NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => NPC_L_IN(31), CK => CLK, RN 
                           => n17, Q => NPC_L_OUT(31), QN => n_1214);
   NPC_L_OUT_reg_30_inst : DFFR_X1 port map( D => NPC_L_IN(30), CK => CLK, RN 
                           => n17, Q => NPC_L_OUT(30), QN => n_1215);
   NPC_L_OUT_reg_29_inst : DFFR_X1 port map( D => NPC_L_IN(29), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(29), QN => n_1216);
   NPC_L_OUT_reg_28_inst : DFFR_X1 port map( D => NPC_L_IN(28), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(28), QN => n_1217);
   NPC_L_OUT_reg_27_inst : DFFR_X1 port map( D => NPC_L_IN(27), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(27), QN => n_1218);
   NPC_L_OUT_reg_26_inst : DFFR_X1 port map( D => NPC_L_IN(26), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(26), QN => n_1219);
   NPC_L_OUT_reg_25_inst : DFFR_X1 port map( D => NPC_L_IN(25), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(25), QN => n_1220);
   NPC_L_OUT_reg_24_inst : DFFR_X1 port map( D => NPC_L_IN(24), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(24), QN => n_1221);
   NPC_L_OUT_reg_23_inst : DFFR_X1 port map( D => NPC_L_IN(23), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(23), QN => n_1222);
   NPC_L_OUT_reg_22_inst : DFFR_X1 port map( D => NPC_L_IN(22), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(22), QN => n_1223);
   NPC_L_OUT_reg_21_inst : DFFR_X1 port map( D => NPC_L_IN(21), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(21), QN => n_1224);
   NPC_L_OUT_reg_20_inst : DFFR_X1 port map( D => NPC_L_IN(20), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(20), QN => n_1225);
   NPC_L_OUT_reg_19_inst : DFFR_X1 port map( D => NPC_L_IN(19), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(19), QN => n_1226);
   NPC_L_OUT_reg_18_inst : DFFR_X1 port map( D => NPC_L_IN(18), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(18), QN => n_1227);
   NPC_L_OUT_reg_17_inst : DFFR_X1 port map( D => NPC_L_IN(17), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(17), QN => n_1228);
   NPC_L_OUT_reg_16_inst : DFFR_X1 port map( D => NPC_L_IN(16), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(16), QN => n_1229);
   NPC_L_OUT_reg_15_inst : DFFR_X1 port map( D => NPC_L_IN(15), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(15), QN => n_1230);
   NPC_L_OUT_reg_14_inst : DFFR_X1 port map( D => NPC_L_IN(14), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(14), QN => n_1231);
   NPC_L_OUT_reg_13_inst : DFFR_X1 port map( D => NPC_L_IN(13), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(13), QN => n_1232);
   NPC_L_OUT_reg_12_inst : DFFR_X1 port map( D => NPC_L_IN(12), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(12), QN => n_1233);
   NPC_L_OUT_reg_11_inst : DFFR_X1 port map( D => NPC_L_IN(11), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(11), QN => n_1234);
   NPC_L_OUT_reg_10_inst : DFFR_X1 port map( D => NPC_L_IN(10), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(10), QN => n_1235);
   NPC_L_OUT_reg_9_inst : DFFR_X1 port map( D => NPC_L_IN(9), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(9), QN => n_1236);
   NPC_L_OUT_reg_8_inst : DFFR_X1 port map( D => NPC_L_IN(8), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(8), QN => n_1237);
   NPC_L_OUT_reg_7_inst : DFFR_X1 port map( D => NPC_L_IN(7), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(7), QN => n_1238);
   NPC_L_OUT_reg_6_inst : DFFR_X1 port map( D => NPC_L_IN(6), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(6), QN => n_1239);
   NPC_L_OUT_reg_5_inst : DFFR_X1 port map( D => NPC_L_IN(5), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(5), QN => n_1240);
   NPC_L_OUT_reg_4_inst : DFFR_X1 port map( D => NPC_L_IN(4), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(4), QN => n_1241);
   NPC_L_OUT_reg_3_inst : DFFR_X1 port map( D => NPC_L_IN(3), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(3), QN => n_1242);
   NPC_L_OUT_reg_2_inst : DFFR_X1 port map( D => NPC_L_IN(2), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(2), QN => n_1243);
   NPC_L_OUT_reg_1_inst : DFFR_X1 port map( D => NPC_L_IN(1), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(1), QN => n_1244);
   NPC_L_OUT_reg_0_inst : DFFR_X1 port map( D => NPC_L_IN(0), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(0), QN => n_1245);
   RD_OUT_reg_3_inst : DFFR_X1 port map( D => RD_IN(3), CK => CLK, RN => n20, Q
                           => RD_OUT(3), QN => n_1246);
   RD_OUT_reg_2_inst : DFFR_X1 port map( D => RD_IN(2), CK => CLK, RN => n20, Q
                           => RD_OUT(2), QN => n_1247);
   RD_OUT_reg_0_inst : DFFR_X1 port map( D => RD_IN(0), CK => CLK, RN => n20, Q
                           => RD_OUT(0), QN => n_1248);
   OPCODE_OUT_reg_2_inst : DFFR_X1 port map( D => OPCODE_IN(2), CK => CLK, RN 
                           => n12, Q => n_1249, QN => n5);
   RD_OUT_reg_1_inst : DFFR_X2 port map( D => RD_IN(1), CK => CLK, RN => n20, Q
                           => RD_OUT(1), QN => n_1250);
   RD_OUT_reg_4_inst : DFFR_X2 port map( D => RD_IN(4), CK => CLK, RN => n20, Q
                           => RD_OUT(4), QN => n_1251);
   U3 : INV_X1 port map( A => n3, ZN => OPCODE_OUT(0));
   U4 : INV_X1 port map( A => n5, ZN => OPCODE_OUT(2));
   U5 : INV_X1 port map( A => n1, ZN => OPCODE_OUT(1));
   U6 : INV_X1 port map( A => n7, ZN => OPCODE_OUT(3));
   U7 : CLKBUF_X1 port map( A => RST, Z => n9);
   U8 : CLKBUF_X1 port map( A => RST, Z => n10);
   U9 : CLKBUF_X1 port map( A => RST, Z => n11);
   U10 : CLKBUF_X1 port map( A => n9, Z => n12);
   U11 : CLKBUF_X1 port map( A => n9, Z => n13);
   U12 : CLKBUF_X1 port map( A => n9, Z => n14);
   U13 : CLKBUF_X1 port map( A => n10, Z => n15);
   U14 : CLKBUF_X1 port map( A => n10, Z => n16);
   U15 : CLKBUF_X1 port map( A => n10, Z => n17);
   U16 : CLKBUF_X1 port map( A => n11, Z => n18);
   U17 : CLKBUF_X1 port map( A => n11, Z => n19);
   U18 : CLKBUF_X1 port map( A => n11, Z => n20);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity EX_MEM is

   port( CLK, RST : in std_logic;  NPC_IN, NPC_L_IN, ALU_IN, B_IN : in 
         std_logic_vector (31 downto 0);  RD_IN : in std_logic_vector (4 downto
         0);  OPCODE_IN : in std_logic_vector (5 downto 0);  NPC_OUT, NPC_L_OUT
         , ALU_OUT, B_OUT : out std_logic_vector (31 downto 0);  RD_OUT : out 
         std_logic_vector (4 downto 0);  OPCODE_OUT : out std_logic_vector (5 
         downto 0));

end EX_MEM;

architecture SYN_Behavioral of EX_MEM is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n5, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21
      , n22, n23, n24, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390 : std_logic;

begin
   
   OPCODE_OUT_reg_5_inst : DFFR_X1 port map( D => OPCODE_IN(5), CK => CLK, RN 
                           => n13, Q => OPCODE_OUT(5), QN => n_1252);
   OPCODE_OUT_reg_4_inst : DFFR_X1 port map( D => OPCODE_IN(4), CK => CLK, RN 
                           => n13, Q => n_1253, QN => n3);
   OPCODE_OUT_reg_3_inst : DFFR_X1 port map( D => OPCODE_IN(3), CK => CLK, RN 
                           => n13, Q => n_1254, QN => n7);
   OPCODE_OUT_reg_0_inst : DFFR_X1 port map( D => OPCODE_IN(0), CK => CLK, RN 
                           => n13, Q => OPCODE_OUT(0), QN => n_1255);
   ALU_OUT_reg_31_inst : DFFR_X1 port map( D => ALU_IN(31), CK => CLK, RN => 
                           n13, Q => ALU_OUT(31), QN => n_1256);
   ALU_OUT_reg_30_inst : DFFR_X1 port map( D => ALU_IN(30), CK => CLK, RN => 
                           n13, Q => ALU_OUT(30), QN => n_1257);
   ALU_OUT_reg_29_inst : DFFR_X1 port map( D => ALU_IN(29), CK => CLK, RN => 
                           n13, Q => ALU_OUT(29), QN => n_1258);
   ALU_OUT_reg_28_inst : DFFR_X1 port map( D => ALU_IN(28), CK => CLK, RN => 
                           n13, Q => ALU_OUT(28), QN => n_1259);
   ALU_OUT_reg_27_inst : DFFR_X1 port map( D => ALU_IN(27), CK => CLK, RN => 
                           n13, Q => ALU_OUT(27), QN => n_1260);
   ALU_OUT_reg_26_inst : DFFR_X1 port map( D => ALU_IN(26), CK => CLK, RN => 
                           n13, Q => ALU_OUT(26), QN => n_1261);
   ALU_OUT_reg_25_inst : DFFR_X1 port map( D => ALU_IN(25), CK => CLK, RN => 
                           n14, Q => ALU_OUT(25), QN => n_1262);
   ALU_OUT_reg_24_inst : DFFR_X1 port map( D => ALU_IN(24), CK => CLK, RN => 
                           n14, Q => ALU_OUT(24), QN => n_1263);
   ALU_OUT_reg_23_inst : DFFR_X1 port map( D => ALU_IN(23), CK => CLK, RN => 
                           n14, Q => ALU_OUT(23), QN => n_1264);
   ALU_OUT_reg_22_inst : DFFR_X1 port map( D => ALU_IN(22), CK => CLK, RN => 
                           n14, Q => ALU_OUT(22), QN => n_1265);
   ALU_OUT_reg_21_inst : DFFR_X1 port map( D => ALU_IN(21), CK => CLK, RN => 
                           n14, Q => ALU_OUT(21), QN => n_1266);
   ALU_OUT_reg_20_inst : DFFR_X1 port map( D => ALU_IN(20), CK => CLK, RN => 
                           n14, Q => ALU_OUT(20), QN => n_1267);
   ALU_OUT_reg_19_inst : DFFR_X1 port map( D => ALU_IN(19), CK => CLK, RN => 
                           n14, Q => ALU_OUT(19), QN => n_1268);
   ALU_OUT_reg_18_inst : DFFR_X1 port map( D => ALU_IN(18), CK => CLK, RN => 
                           n14, Q => ALU_OUT(18), QN => n_1269);
   ALU_OUT_reg_17_inst : DFFR_X1 port map( D => ALU_IN(17), CK => CLK, RN => 
                           n14, Q => ALU_OUT(17), QN => n_1270);
   ALU_OUT_reg_16_inst : DFFR_X1 port map( D => ALU_IN(16), CK => CLK, RN => 
                           n14, Q => ALU_OUT(16), QN => n_1271);
   ALU_OUT_reg_15_inst : DFFR_X1 port map( D => ALU_IN(15), CK => CLK, RN => 
                           n14, Q => ALU_OUT(15), QN => n_1272);
   ALU_OUT_reg_14_inst : DFFR_X1 port map( D => ALU_IN(14), CK => CLK, RN => 
                           n14, Q => ALU_OUT(14), QN => n_1273);
   ALU_OUT_reg_13_inst : DFFR_X1 port map( D => ALU_IN(13), CK => CLK, RN => 
                           n15, Q => ALU_OUT(13), QN => n_1274);
   ALU_OUT_reg_12_inst : DFFR_X1 port map( D => ALU_IN(12), CK => CLK, RN => 
                           n15, Q => ALU_OUT(12), QN => n_1275);
   ALU_OUT_reg_11_inst : DFFR_X1 port map( D => ALU_IN(11), CK => CLK, RN => 
                           n15, Q => ALU_OUT(11), QN => n_1276);
   ALU_OUT_reg_10_inst : DFFR_X1 port map( D => ALU_IN(10), CK => CLK, RN => 
                           n15, Q => ALU_OUT(10), QN => n_1277);
   ALU_OUT_reg_9_inst : DFFR_X1 port map( D => ALU_IN(9), CK => CLK, RN => n15,
                           Q => ALU_OUT(9), QN => n_1278);
   ALU_OUT_reg_8_inst : DFFR_X1 port map( D => ALU_IN(8), CK => CLK, RN => n15,
                           Q => ALU_OUT(8), QN => n_1279);
   ALU_OUT_reg_7_inst : DFFR_X1 port map( D => ALU_IN(7), CK => CLK, RN => n15,
                           Q => ALU_OUT(7), QN => n_1280);
   ALU_OUT_reg_6_inst : DFFR_X1 port map( D => ALU_IN(6), CK => CLK, RN => n15,
                           Q => ALU_OUT(6), QN => n_1281);
   ALU_OUT_reg_5_inst : DFFR_X1 port map( D => ALU_IN(5), CK => CLK, RN => n15,
                           Q => ALU_OUT(5), QN => n_1282);
   ALU_OUT_reg_4_inst : DFFR_X1 port map( D => ALU_IN(4), CK => CLK, RN => n15,
                           Q => ALU_OUT(4), QN => n_1283);
   ALU_OUT_reg_3_inst : DFFR_X1 port map( D => ALU_IN(3), CK => CLK, RN => n15,
                           Q => ALU_OUT(3), QN => n_1284);
   ALU_OUT_reg_2_inst : DFFR_X1 port map( D => ALU_IN(2), CK => CLK, RN => n15,
                           Q => ALU_OUT(2), QN => n_1285);
   ALU_OUT_reg_1_inst : DFFR_X1 port map( D => ALU_IN(1), CK => CLK, RN => n16,
                           Q => ALU_OUT(1), QN => n_1286);
   ALU_OUT_reg_0_inst : DFFR_X1 port map( D => ALU_IN(0), CK => CLK, RN => n16,
                           Q => ALU_OUT(0), QN => n_1287);
   B_OUT_reg_31_inst : DFFR_X1 port map( D => B_IN(31), CK => CLK, RN => n16, Q
                           => B_OUT(31), QN => n_1288);
   B_OUT_reg_30_inst : DFFR_X1 port map( D => B_IN(30), CK => CLK, RN => n16, Q
                           => B_OUT(30), QN => n_1289);
   B_OUT_reg_29_inst : DFFR_X1 port map( D => B_IN(29), CK => CLK, RN => n16, Q
                           => B_OUT(29), QN => n_1290);
   B_OUT_reg_28_inst : DFFR_X1 port map( D => B_IN(28), CK => CLK, RN => n16, Q
                           => B_OUT(28), QN => n_1291);
   B_OUT_reg_27_inst : DFFR_X1 port map( D => B_IN(27), CK => CLK, RN => n16, Q
                           => B_OUT(27), QN => n_1292);
   B_OUT_reg_26_inst : DFFR_X1 port map( D => B_IN(26), CK => CLK, RN => n16, Q
                           => B_OUT(26), QN => n_1293);
   B_OUT_reg_25_inst : DFFR_X1 port map( D => B_IN(25), CK => CLK, RN => n16, Q
                           => B_OUT(25), QN => n_1294);
   B_OUT_reg_24_inst : DFFR_X1 port map( D => B_IN(24), CK => CLK, RN => n16, Q
                           => B_OUT(24), QN => n_1295);
   B_OUT_reg_23_inst : DFFR_X1 port map( D => B_IN(23), CK => CLK, RN => n16, Q
                           => B_OUT(23), QN => n_1296);
   B_OUT_reg_22_inst : DFFR_X1 port map( D => B_IN(22), CK => CLK, RN => n16, Q
                           => B_OUT(22), QN => n_1297);
   B_OUT_reg_21_inst : DFFR_X1 port map( D => B_IN(21), CK => CLK, RN => n17, Q
                           => B_OUT(21), QN => n_1298);
   B_OUT_reg_20_inst : DFFR_X1 port map( D => B_IN(20), CK => CLK, RN => n17, Q
                           => B_OUT(20), QN => n_1299);
   B_OUT_reg_19_inst : DFFR_X1 port map( D => B_IN(19), CK => CLK, RN => n17, Q
                           => B_OUT(19), QN => n_1300);
   B_OUT_reg_18_inst : DFFR_X1 port map( D => B_IN(18), CK => CLK, RN => n17, Q
                           => B_OUT(18), QN => n_1301);
   B_OUT_reg_17_inst : DFFR_X1 port map( D => B_IN(17), CK => CLK, RN => n17, Q
                           => B_OUT(17), QN => n_1302);
   B_OUT_reg_16_inst : DFFR_X1 port map( D => B_IN(16), CK => CLK, RN => n17, Q
                           => B_OUT(16), QN => n_1303);
   B_OUT_reg_15_inst : DFFR_X1 port map( D => B_IN(15), CK => CLK, RN => n17, Q
                           => B_OUT(15), QN => n_1304);
   B_OUT_reg_14_inst : DFFR_X1 port map( D => B_IN(14), CK => CLK, RN => n17, Q
                           => B_OUT(14), QN => n_1305);
   B_OUT_reg_13_inst : DFFR_X1 port map( D => B_IN(13), CK => CLK, RN => n17, Q
                           => B_OUT(13), QN => n_1306);
   B_OUT_reg_12_inst : DFFR_X1 port map( D => B_IN(12), CK => CLK, RN => n17, Q
                           => B_OUT(12), QN => n_1307);
   B_OUT_reg_11_inst : DFFR_X1 port map( D => B_IN(11), CK => CLK, RN => n17, Q
                           => B_OUT(11), QN => n_1308);
   B_OUT_reg_10_inst : DFFR_X1 port map( D => B_IN(10), CK => CLK, RN => n17, Q
                           => B_OUT(10), QN => n_1309);
   B_OUT_reg_9_inst : DFFR_X1 port map( D => B_IN(9), CK => CLK, RN => n18, Q 
                           => B_OUT(9), QN => n_1310);
   B_OUT_reg_8_inst : DFFR_X1 port map( D => B_IN(8), CK => CLK, RN => n18, Q 
                           => B_OUT(8), QN => n_1311);
   B_OUT_reg_7_inst : DFFR_X1 port map( D => B_IN(7), CK => CLK, RN => n18, Q 
                           => B_OUT(7), QN => n_1312);
   B_OUT_reg_6_inst : DFFR_X1 port map( D => B_IN(6), CK => CLK, RN => n18, Q 
                           => B_OUT(6), QN => n_1313);
   B_OUT_reg_5_inst : DFFR_X1 port map( D => B_IN(5), CK => CLK, RN => n18, Q 
                           => B_OUT(5), QN => n_1314);
   B_OUT_reg_4_inst : DFFR_X1 port map( D => B_IN(4), CK => CLK, RN => n18, Q 
                           => B_OUT(4), QN => n_1315);
   B_OUT_reg_3_inst : DFFR_X1 port map( D => B_IN(3), CK => CLK, RN => n18, Q 
                           => B_OUT(3), QN => n_1316);
   B_OUT_reg_2_inst : DFFR_X1 port map( D => B_IN(2), CK => CLK, RN => n18, Q 
                           => B_OUT(2), QN => n_1317);
   B_OUT_reg_1_inst : DFFR_X1 port map( D => B_IN(1), CK => CLK, RN => n18, Q 
                           => B_OUT(1), QN => n_1318);
   B_OUT_reg_0_inst : DFFR_X1 port map( D => B_IN(0), CK => CLK, RN => n18, Q 
                           => B_OUT(0), QN => n_1319);
   NPC_OUT_reg_31_inst : DFFR_X1 port map( D => NPC_IN(31), CK => CLK, RN => 
                           n18, Q => NPC_OUT(31), QN => n_1320);
   NPC_OUT_reg_30_inst : DFFR_X1 port map( D => NPC_IN(30), CK => CLK, RN => 
                           n18, Q => NPC_OUT(30), QN => n_1321);
   NPC_OUT_reg_29_inst : DFFR_X1 port map( D => NPC_IN(29), CK => CLK, RN => 
                           n19, Q => NPC_OUT(29), QN => n_1322);
   NPC_OUT_reg_28_inst : DFFR_X1 port map( D => NPC_IN(28), CK => CLK, RN => 
                           n19, Q => NPC_OUT(28), QN => n_1323);
   NPC_OUT_reg_27_inst : DFFR_X1 port map( D => NPC_IN(27), CK => CLK, RN => 
                           n19, Q => NPC_OUT(27), QN => n_1324);
   NPC_OUT_reg_26_inst : DFFR_X1 port map( D => NPC_IN(26), CK => CLK, RN => 
                           n19, Q => NPC_OUT(26), QN => n_1325);
   NPC_OUT_reg_25_inst : DFFR_X1 port map( D => NPC_IN(25), CK => CLK, RN => 
                           n19, Q => NPC_OUT(25), QN => n_1326);
   NPC_OUT_reg_24_inst : DFFR_X1 port map( D => NPC_IN(24), CK => CLK, RN => 
                           n19, Q => NPC_OUT(24), QN => n_1327);
   NPC_OUT_reg_23_inst : DFFR_X1 port map( D => NPC_IN(23), CK => CLK, RN => 
                           n19, Q => NPC_OUT(23), QN => n_1328);
   NPC_OUT_reg_22_inst : DFFR_X1 port map( D => NPC_IN(22), CK => CLK, RN => 
                           n19, Q => NPC_OUT(22), QN => n_1329);
   NPC_OUT_reg_21_inst : DFFR_X1 port map( D => NPC_IN(21), CK => CLK, RN => 
                           n19, Q => NPC_OUT(21), QN => n_1330);
   NPC_OUT_reg_20_inst : DFFR_X1 port map( D => NPC_IN(20), CK => CLK, RN => 
                           n19, Q => NPC_OUT(20), QN => n_1331);
   NPC_OUT_reg_19_inst : DFFR_X1 port map( D => NPC_IN(19), CK => CLK, RN => 
                           n19, Q => NPC_OUT(19), QN => n_1332);
   NPC_OUT_reg_18_inst : DFFR_X1 port map( D => NPC_IN(18), CK => CLK, RN => 
                           n19, Q => NPC_OUT(18), QN => n_1333);
   NPC_OUT_reg_17_inst : DFFR_X1 port map( D => NPC_IN(17), CK => CLK, RN => 
                           n20, Q => NPC_OUT(17), QN => n_1334);
   NPC_OUT_reg_16_inst : DFFR_X1 port map( D => NPC_IN(16), CK => CLK, RN => 
                           n20, Q => NPC_OUT(16), QN => n_1335);
   NPC_OUT_reg_15_inst : DFFR_X1 port map( D => NPC_IN(15), CK => CLK, RN => 
                           n20, Q => NPC_OUT(15), QN => n_1336);
   NPC_OUT_reg_14_inst : DFFR_X1 port map( D => NPC_IN(14), CK => CLK, RN => 
                           n20, Q => NPC_OUT(14), QN => n_1337);
   NPC_OUT_reg_13_inst : DFFR_X1 port map( D => NPC_IN(13), CK => CLK, RN => 
                           n20, Q => NPC_OUT(13), QN => n_1338);
   NPC_OUT_reg_12_inst : DFFR_X1 port map( D => NPC_IN(12), CK => CLK, RN => 
                           n20, Q => NPC_OUT(12), QN => n_1339);
   NPC_OUT_reg_11_inst : DFFR_X1 port map( D => NPC_IN(11), CK => CLK, RN => 
                           n20, Q => NPC_OUT(11), QN => n_1340);
   NPC_OUT_reg_10_inst : DFFR_X1 port map( D => NPC_IN(10), CK => CLK, RN => 
                           n20, Q => NPC_OUT(10), QN => n_1341);
   NPC_OUT_reg_9_inst : DFFR_X1 port map( D => NPC_IN(9), CK => CLK, RN => n20,
                           Q => NPC_OUT(9), QN => n_1342);
   NPC_OUT_reg_8_inst : DFFR_X1 port map( D => NPC_IN(8), CK => CLK, RN => n20,
                           Q => NPC_OUT(8), QN => n_1343);
   NPC_OUT_reg_7_inst : DFFR_X1 port map( D => NPC_IN(7), CK => CLK, RN => n20,
                           Q => NPC_OUT(7), QN => n_1344);
   NPC_OUT_reg_6_inst : DFFR_X1 port map( D => NPC_IN(6), CK => CLK, RN => n20,
                           Q => NPC_OUT(6), QN => n_1345);
   NPC_OUT_reg_5_inst : DFFR_X1 port map( D => NPC_IN(5), CK => CLK, RN => n21,
                           Q => NPC_OUT(5), QN => n_1346);
   NPC_OUT_reg_4_inst : DFFR_X1 port map( D => NPC_IN(4), CK => CLK, RN => n21,
                           Q => NPC_OUT(4), QN => n_1347);
   NPC_OUT_reg_3_inst : DFFR_X1 port map( D => NPC_IN(3), CK => CLK, RN => n21,
                           Q => NPC_OUT(3), QN => n_1348);
   NPC_OUT_reg_2_inst : DFFR_X1 port map( D => NPC_IN(2), CK => CLK, RN => n21,
                           Q => NPC_OUT(2), QN => n_1349);
   NPC_OUT_reg_1_inst : DFFR_X1 port map( D => NPC_IN(1), CK => CLK, RN => n21,
                           Q => NPC_OUT(1), QN => n_1350);
   NPC_OUT_reg_0_inst : DFFR_X1 port map( D => NPC_IN(0), CK => CLK, RN => n21,
                           Q => NPC_OUT(0), QN => n_1351);
   NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => NPC_L_IN(31), CK => CLK, RN 
                           => n21, Q => NPC_L_OUT(31), QN => n_1352);
   NPC_L_OUT_reg_30_inst : DFFR_X1 port map( D => NPC_L_IN(30), CK => CLK, RN 
                           => n21, Q => NPC_L_OUT(30), QN => n_1353);
   NPC_L_OUT_reg_29_inst : DFFR_X1 port map( D => NPC_L_IN(29), CK => CLK, RN 
                           => n21, Q => NPC_L_OUT(29), QN => n_1354);
   NPC_L_OUT_reg_28_inst : DFFR_X1 port map( D => NPC_L_IN(28), CK => CLK, RN 
                           => n21, Q => NPC_L_OUT(28), QN => n_1355);
   NPC_L_OUT_reg_27_inst : DFFR_X1 port map( D => NPC_L_IN(27), CK => CLK, RN 
                           => n21, Q => NPC_L_OUT(27), QN => n_1356);
   NPC_L_OUT_reg_26_inst : DFFR_X1 port map( D => NPC_L_IN(26), CK => CLK, RN 
                           => n21, Q => NPC_L_OUT(26), QN => n_1357);
   NPC_L_OUT_reg_25_inst : DFFR_X1 port map( D => NPC_L_IN(25), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(25), QN => n_1358);
   NPC_L_OUT_reg_24_inst : DFFR_X1 port map( D => NPC_L_IN(24), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(24), QN => n_1359);
   NPC_L_OUT_reg_23_inst : DFFR_X1 port map( D => NPC_L_IN(23), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(23), QN => n_1360);
   NPC_L_OUT_reg_22_inst : DFFR_X1 port map( D => NPC_L_IN(22), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(22), QN => n_1361);
   NPC_L_OUT_reg_21_inst : DFFR_X1 port map( D => NPC_L_IN(21), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(21), QN => n_1362);
   NPC_L_OUT_reg_20_inst : DFFR_X1 port map( D => NPC_L_IN(20), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(20), QN => n_1363);
   NPC_L_OUT_reg_19_inst : DFFR_X1 port map( D => NPC_L_IN(19), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(19), QN => n_1364);
   NPC_L_OUT_reg_18_inst : DFFR_X1 port map( D => NPC_L_IN(18), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(18), QN => n_1365);
   NPC_L_OUT_reg_17_inst : DFFR_X1 port map( D => NPC_L_IN(17), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(17), QN => n_1366);
   NPC_L_OUT_reg_16_inst : DFFR_X1 port map( D => NPC_L_IN(16), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(16), QN => n_1367);
   NPC_L_OUT_reg_15_inst : DFFR_X1 port map( D => NPC_L_IN(15), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(15), QN => n_1368);
   NPC_L_OUT_reg_14_inst : DFFR_X1 port map( D => NPC_L_IN(14), CK => CLK, RN 
                           => n22, Q => NPC_L_OUT(14), QN => n_1369);
   NPC_L_OUT_reg_13_inst : DFFR_X1 port map( D => NPC_L_IN(13), CK => CLK, RN 
                           => n23, Q => NPC_L_OUT(13), QN => n_1370);
   NPC_L_OUT_reg_12_inst : DFFR_X1 port map( D => NPC_L_IN(12), CK => CLK, RN 
                           => n23, Q => NPC_L_OUT(12), QN => n_1371);
   NPC_L_OUT_reg_11_inst : DFFR_X1 port map( D => NPC_L_IN(11), CK => CLK, RN 
                           => n23, Q => NPC_L_OUT(11), QN => n_1372);
   NPC_L_OUT_reg_10_inst : DFFR_X1 port map( D => NPC_L_IN(10), CK => CLK, RN 
                           => n23, Q => NPC_L_OUT(10), QN => n_1373);
   NPC_L_OUT_reg_9_inst : DFFR_X1 port map( D => NPC_L_IN(9), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(9), QN => n_1374);
   NPC_L_OUT_reg_8_inst : DFFR_X1 port map( D => NPC_L_IN(8), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(8), QN => n_1375);
   NPC_L_OUT_reg_7_inst : DFFR_X1 port map( D => NPC_L_IN(7), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(7), QN => n_1376);
   NPC_L_OUT_reg_6_inst : DFFR_X1 port map( D => NPC_L_IN(6), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(6), QN => n_1377);
   NPC_L_OUT_reg_5_inst : DFFR_X1 port map( D => NPC_L_IN(5), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(5), QN => n_1378);
   NPC_L_OUT_reg_4_inst : DFFR_X1 port map( D => NPC_L_IN(4), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(4), QN => n_1379);
   NPC_L_OUT_reg_3_inst : DFFR_X1 port map( D => NPC_L_IN(3), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(3), QN => n_1380);
   NPC_L_OUT_reg_2_inst : DFFR_X1 port map( D => NPC_L_IN(2), CK => CLK, RN => 
                           n23, Q => NPC_L_OUT(2), QN => n_1381);
   NPC_L_OUT_reg_1_inst : DFFR_X1 port map( D => NPC_L_IN(1), CK => CLK, RN => 
                           n24, Q => NPC_L_OUT(1), QN => n_1382);
   NPC_L_OUT_reg_0_inst : DFFR_X1 port map( D => NPC_L_IN(0), CK => CLK, RN => 
                           n24, Q => NPC_L_OUT(0), QN => n_1383);
   RD_OUT_reg_4_inst : DFFR_X1 port map( D => RD_IN(4), CK => CLK, RN => n24, Q
                           => RD_OUT(4), QN => n_1384);
   RD_OUT_reg_3_inst : DFFR_X1 port map( D => RD_IN(3), CK => CLK, RN => n24, Q
                           => RD_OUT(3), QN => n_1385);
   RD_OUT_reg_1_inst : DFFR_X1 port map( D => RD_IN(1), CK => CLK, RN => n24, Q
                           => RD_OUT(1), QN => n_1386);
   RD_OUT_reg_0_inst : DFFR_X1 port map( D => RD_IN(0), CK => CLK, RN => n24, Q
                           => RD_OUT(0), QN => n_1387);
   OPCODE_OUT_reg_1_inst : DFFR_X1 port map( D => OPCODE_IN(1), CK => CLK, RN 
                           => n13, Q => n_1388, QN => n5);
   OPCODE_OUT_reg_2_inst : DFFR_X1 port map( D => OPCODE_IN(2), CK => CLK, RN 
                           => n13, Q => n_1389, QN => n9);
   RD_OUT_reg_2_inst : DFFR_X1 port map( D => RD_IN(2), CK => CLK, RN => RST, Q
                           => RD_OUT(2), QN => n_1390);
   U3 : INV_X1 port map( A => n3, ZN => OPCODE_OUT(4));
   U4 : INV_X1 port map( A => n5, ZN => OPCODE_OUT(1));
   U5 : INV_X1 port map( A => n9, ZN => OPCODE_OUT(2));
   U6 : INV_X1 port map( A => n7, ZN => OPCODE_OUT(3));
   U7 : BUF_X1 port map( A => RST, Z => n12);
   U8 : BUF_X1 port map( A => RST, Z => n11);
   U9 : CLKBUF_X1 port map( A => n11, Z => n13);
   U10 : CLKBUF_X1 port map( A => n11, Z => n14);
   U11 : CLKBUF_X1 port map( A => n11, Z => n15);
   U12 : CLKBUF_X1 port map( A => n11, Z => n16);
   U13 : CLKBUF_X1 port map( A => n11, Z => n17);
   U14 : CLKBUF_X1 port map( A => n11, Z => n18);
   U15 : CLKBUF_X1 port map( A => n12, Z => n19);
   U16 : CLKBUF_X1 port map( A => n12, Z => n20);
   U17 : CLKBUF_X1 port map( A => n12, Z => n21);
   U18 : CLKBUF_X1 port map( A => n12, Z => n22);
   U19 : CLKBUF_X1 port map( A => n12, Z => n23);
   U20 : CLKBUF_X1 port map( A => n12, Z => n24);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_cond_N32 is

   port( A : in std_logic_vector (31 downto 0);  EN : in std_logic;  OP : in 
         std_logic_vector (0 to 4);  PRE : in std_logic;  DISCARD, WRONG, RIGHT
         , SEL : out std_logic);

end branch_cond_N32;

architecture SYN_Behavioral of branch_cond_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal WRONG_port, SEL_port, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n1, n2, n3, n4, n5 : std_logic;

begin
   WRONG <= WRONG_port;
   SEL <= SEL_port;
   
   U29 : NAND3_X1 port map( A1 => OP(2), A2 => n2, A3 => OP(1), ZN => n12);
   U3 : NOR2_X1 port map( A1 => n5, A2 => n11, ZN => WRONG_port);
   U4 : AOI22_X1 port map( A1 => n1, A2 => n8, B1 => n9, B2 => n7, ZN => n11);
   U5 : NOR4_X1 port map( A1 => A(23), A2 => A(22), A3 => A(21), A4 => A(20), 
                           ZN => n19);
   U6 : NOR4_X1 port map( A1 => A(9), A2 => A(8), A3 => A(7), A4 => A(6), ZN =>
                           n23);
   U7 : NOR4_X1 port map( A1 => A(1), A2 => A(19), A3 => A(18), A4 => A(17), ZN
                           => n18);
   U8 : NOR4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(3), A4 => A(31), ZN 
                           => n22);
   U9 : NOR4_X1 port map( A1 => A(16), A2 => A(15), A3 => A(14), A4 => A(13), 
                           ZN => n17);
   U10 : NOR4_X1 port map( A1 => A(30), A2 => A(2), A3 => A(29), A4 => A(28), 
                           ZN => n21);
   U11 : NOR4_X1 port map( A1 => A(12), A2 => A(11), A3 => A(10), A4 => A(0), 
                           ZN => n16);
   U12 : NOR4_X1 port map( A1 => A(27), A2 => A(26), A3 => A(25), A4 => A(24), 
                           ZN => n20);
   U13 : INV_X1 port map( A => n9, ZN => n1);
   U14 : OR2_X1 port map( A1 => WRONG_port, A2 => SEL_port, ZN => DISCARD);
   U15 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => RIGHT);
   U16 : AOI22_X1 port map( A1 => n7, A2 => n1, B1 => n8, B2 => n9, ZN => n6);
   U17 : NOR3_X1 port map( A1 => n12, A2 => OP(4), A3 => n3, ZN => n7);
   U18 : INV_X1 port map( A => OP(0), ZN => n2);
   U19 : XNOR2_X1 port map( A => PRE, B => n13, ZN => n9);
   U20 : NOR2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U21 : NAND4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => 
                           n14);
   U22 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           n15);
   U23 : INV_X1 port map( A => OP(3), ZN => n3);
   U24 : NOR3_X1 port map( A1 => n12, A2 => OP(3), A3 => n4, ZN => n8);
   U25 : INV_X1 port map( A => OP(4), ZN => n4);
   U26 : AND4_X1 port map( A1 => OP(0), A2 => EN, A3 => n10, A4 => n3, ZN => 
                           SEL_port);
   U27 : NOR2_X1 port map( A1 => OP(1), A2 => OP(2), ZN => n10);
   U28 : INV_X1 port map( A => EN, ZN => n5);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FWD_UNIT_BRANCH is

   port( Rst : in std_logic;  Rs1, Rd_M, Rd_W : in std_logic_vector (4 downto 
         0);  ICODE, ICODE_M, ICODE_W : in std_logic_vector (5 downto 0);  SEL 
         : out std_logic_vector (1 downto 0));

end FWD_UNIT_BRANCH;

architecture SYN_Behavioral of FWD_UNIT_BRANCH is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FWD_CAM_1
      port( RST : in std_logic;  DATA_IN_1, DATA_IN_2, DATA_IN_3 : in 
            std_logic_vector (5 downto 0);  MATCH_1, MATCH_2, MATCH_3 : out 
            std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal match_op_M, match_op_W, N12, N13, N14, n1, n2, n3, n4, n5, n6, n7, n8
      , n9, n10, n11, n12_port, n13_port, n14_port, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n_1391 : std_logic;

begin
   
   SEL_reg_1_inst : DLH_X1 port map( G => N12, D => N14, Q => SEL(1));
   SEL_reg_0_inst : DLH_X1 port map( G => N12, D => N13, Q => SEL(0));
   CAM : FWD_CAM_1 port map( RST => Rst, DATA_IN_1(5) => ICODE(5), DATA_IN_1(4)
                           => ICODE(4), DATA_IN_1(3) => ICODE(3), DATA_IN_1(2) 
                           => ICODE(2), DATA_IN_1(1) => ICODE(1), DATA_IN_1(0) 
                           => ICODE(0), DATA_IN_2(5) => ICODE_M(5), 
                           DATA_IN_2(4) => ICODE_M(4), DATA_IN_2(3) => 
                           ICODE_M(3), DATA_IN_2(2) => ICODE_M(2), DATA_IN_2(1)
                           => ICODE_M(1), DATA_IN_2(0) => ICODE_M(0), 
                           DATA_IN_3(5) => ICODE_W(5), DATA_IN_3(4) => 
                           ICODE_W(4), DATA_IN_3(3) => ICODE_W(3), DATA_IN_3(2)
                           => ICODE_W(2), DATA_IN_3(1) => ICODE_W(1), 
                           DATA_IN_3(0) => ICODE_W(0), MATCH_1 => n_1391, 
                           MATCH_2 => match_op_M, MATCH_3 => match_op_W);
   U3 : INV_X1 port map( A => Rst, ZN => n1);
   U4 : NOR4_X1 port map( A1 => n2, A2 => n3, A3 => n1, A4 => n4, ZN => N14);
   U5 : XOR2_X1 port map( A => Rs1(3), B => Rd_W(3), Z => n4);
   U6 : OAI221_X1 port map( B1 => match_op_W, B2 => n5, C1 => n6, C2 => n7, A 
                           => n8, ZN => n3);
   U7 : OR2_X1 port map( A1 => Rd_W(0), A2 => Rd_W(1), ZN => n7);
   U8 : OR3_X1 port map( A1 => Rd_W(3), A2 => Rd_W(4), A3 => Rd_W(2), ZN => n6)
                           ;
   U9 : NOR4_X1 port map( A1 => n9, A2 => ICODE_W(0), A3 => ICODE_W(2), A4 => 
                           ICODE_W(1), ZN => n5);
   U10 : OR3_X1 port map( A1 => ICODE_W(5), A2 => ICODE_W(4), A3 => ICODE_W(3),
                           ZN => n9);
   U11 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12_port, A4 => 
                           n13_port, ZN => n2);
   U12 : XNOR2_X1 port map( A => Rd_W(0), B => Rs1(0), ZN => n13_port);
   U13 : XNOR2_X1 port map( A => Rd_W(1), B => Rs1(1), ZN => n12_port);
   U14 : XNOR2_X1 port map( A => Rd_W(2), B => Rs1(2), ZN => n11);
   U15 : XOR2_X1 port map( A => Rd_W(4), B => n14_port, Z => n10);
   U16 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => N13);
   U17 : OR4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => n8)
                           ;
   U18 : OAI211_X1 port map( C1 => match_op_M, C2 => n19, A => n20, B => n21, 
                           ZN => n18);
   U19 : XNOR2_X1 port map( A => Rd_M(0), B => Rs1(0), ZN => n21);
   U20 : XNOR2_X1 port map( A => Rd_M(1), B => Rs1(1), ZN => n20);
   U21 : NOR4_X1 port map( A1 => n22, A2 => ICODE_M(0), A3 => ICODE_M(2), A4 =>
                           ICODE_M(1), ZN => n19);
   U22 : OR3_X1 port map( A1 => ICODE_M(5), A2 => ICODE_M(4), A3 => ICODE_M(3),
                           ZN => n22);
   U23 : MUX2_X1 port map( A => n23, B => n14_port, S => Rd_M(4), Z => n17);
   U24 : NAND2_X1 port map( A1 => n14_port, A2 => n24, ZN => n23);
   U25 : OR4_X1 port map( A1 => Rd_M(0), A2 => Rd_M(1), A3 => Rd_M(2), A4 => 
                           Rd_M(3), ZN => n24);
   U26 : INV_X1 port map( A => Rs1(4), ZN => n14_port);
   U27 : XOR2_X1 port map( A => Rs1(3), B => Rd_M(3), Z => n16);
   U28 : XOR2_X1 port map( A => Rs1(2), B => Rd_M(2), Z => n15);
   U29 : NAND2_X1 port map( A1 => Rst, A2 => n25, ZN => N12);
   U30 : NAND3_X1 port map( A1 => ICODE(2), A2 => n26, A3 => n27, ZN => n25);
   U31 : NOR3_X1 port map( A1 => ICODE(3), A2 => ICODE(5), A3 => ICODE(4), ZN 
                           => n27);
   U32 : INV_X1 port map( A => ICODE(1), ZN => n26);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity ALU_N32 is

   port( INA, INB : in std_logic_vector (31 downto 0);  OP : in 
         std_logic_vector (0 to 4);  alu_out : out std_logic_vector (31 downto 
         0));

end ALU_N32;

architecture SYN_Behavioral of ALU_N32 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux4to1_N32
      port( inadd, inlog, insh, incom : in std_logic_vector (31 downto 0);  sel
            : in std_logic_vector (0 to 4);  O : out std_logic_vector (31 
            downto 0));
   end component;
   
   component comparator_N32
      port( inA, inB : in std_logic_vector (31 downto 0);  op : in 
            std_logic_vector (0 to 4);  res : out std_logic_vector (31 downto 
            0));
   end component;
   
   component SHIFTER_GENERIC_N32
      port( A, B : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (0 to 4);  OUTPUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component logic_N32
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (0 to 4);  O : out std_logic_vector (31 downto 0)
            );
   end component;
   
   component add_wrapper_N32
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (0 to 4);  O : out std_logic_vector (31 downto 0)
            );
   end component;
   
   signal res1_31_port, res1_30_port, res1_29_port, res1_28_port, res1_27_port,
      res1_26_port, res1_25_port, res1_24_port, res1_23_port, res1_22_port, 
      res1_21_port, res1_20_port, res1_19_port, res1_18_port, res1_17_port, 
      res1_16_port, res1_15_port, res1_14_port, res1_13_port, res1_12_port, 
      res1_11_port, res1_10_port, res1_9_port, res1_8_port, res1_7_port, 
      res1_6_port, res1_5_port, res1_4_port, res1_3_port, res1_2_port, 
      res1_1_port, res1_0_port, res2_31_port, res2_30_port, res2_29_port, 
      res2_28_port, res2_27_port, res2_26_port, res2_25_port, res2_24_port, 
      res2_23_port, res2_22_port, res2_21_port, res2_20_port, res2_19_port, 
      res2_18_port, res2_17_port, res2_16_port, res2_15_port, res2_14_port, 
      res2_13_port, res2_12_port, res2_11_port, res2_10_port, res2_9_port, 
      res2_8_port, res2_7_port, res2_6_port, res2_5_port, res2_4_port, 
      res2_3_port, res2_2_port, res2_1_port, res2_0_port, res3_31_port, 
      res3_30_port, res3_29_port, res3_28_port, res3_27_port, res3_26_port, 
      res3_25_port, res3_24_port, res3_23_port, res3_22_port, res3_21_port, 
      res3_20_port, res3_19_port, res3_18_port, res3_17_port, res3_16_port, 
      res3_15_port, res3_14_port, res3_13_port, res3_12_port, res3_11_port, 
      res3_10_port, res3_9_port, res3_8_port, res3_7_port, res3_6_port, 
      res3_5_port, res3_4_port, res3_3_port, res3_2_port, res3_1_port, 
      res3_0_port, res4_31_port, res4_30_port, res4_29_port, res4_28_port, 
      res4_27_port, res4_26_port, res4_25_port, res4_24_port, res4_23_port, 
      res4_22_port, res4_21_port, res4_20_port, res4_19_port, res4_18_port, 
      res4_17_port, res4_16_port, res4_15_port, res4_14_port, res4_13_port, 
      res4_12_port, res4_11_port, res4_10_port, res4_9_port, res4_8_port, 
      res4_7_port, res4_6_port, res4_5_port, res4_4_port, res4_3_port, 
      res4_2_port, res4_1_port, res4_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422 : std_logic;

begin
   
   adder : add_wrapper_N32 port map( A(31) => INA(31), A(30) => n6, A(29) => 
                           INA(29), A(28) => n5, A(27) => INA(27), A(26) => 
                           INA(26), A(25) => n9, A(24) => INA(24), A(23) => 
                           INA(23), A(22) => INA(22), A(21) => n12, A(20) => 
                           INA(20), A(19) => INA(19), A(18) => INA(18), A(17) 
                           => INA(17), A(16) => INA(16), A(15) => INA(15), 
                           A(14) => INA(14), A(13) => n4, A(12) => n8, A(11) =>
                           n35, A(10) => n1, A(9) => INA(9), A(8) => INA(8), 
                           A(7) => INA(7), A(6) => INA(6), A(5) => n38, A(4) =>
                           n33, A(3) => n47, A(2) => n45, A(1) => n39, A(0) => 
                           n40, B(31) => INB(31), B(30) => INB(30), B(29) => 
                           INB(29), B(28) => INB(28), B(27) => INB(27), B(26) 
                           => INB(26), B(25) => INB(25), B(24) => INB(24), 
                           B(23) => INB(23), B(22) => INB(22), B(21) => INB(21)
                           , B(20) => INB(20), B(19) => INB(19), B(18) => 
                           INB(18), B(17) => INB(17), B(16) => INB(16), B(15) 
                           => INB(15), B(14) => INB(14), B(13) => INB(13), 
                           B(12) => INB(12), B(11) => INB(11), B(10) => INB(10)
                           , B(9) => INB(9), B(8) => INB(8), B(7) => INB(7), 
                           B(6) => INB(6), B(5) => INB(5), B(4) => INB(4), B(3)
                           => INB(3), B(2) => INB(2), B(1) => INB(1), B(0) => 
                           INB(0), SEL(0) => OP(0), SEL(1) => OP(1), SEL(2) => 
                           OP(2), SEL(3) => OP(3), SEL(4) => OP(4), O(31) => 
                           res1_31_port, O(30) => res1_30_port, O(29) => 
                           res1_29_port, O(28) => res1_28_port, O(27) => 
                           res1_27_port, O(26) => res1_26_port, O(25) => 
                           res1_25_port, O(24) => res1_24_port, O(23) => 
                           res1_23_port, O(22) => res1_22_port, O(21) => 
                           res1_21_port, O(20) => res1_20_port, O(19) => 
                           res1_19_port, O(18) => res1_18_port, O(17) => 
                           res1_17_port, O(16) => res1_16_port, O(15) => 
                           res1_15_port, O(14) => res1_14_port, O(13) => 
                           res1_13_port, O(12) => res1_12_port, O(11) => 
                           res1_11_port, O(10) => res1_10_port, O(9) => 
                           res1_9_port, O(8) => res1_8_port, O(7) => 
                           res1_7_port, O(6) => res1_6_port, O(5) => 
                           res1_5_port, O(4) => res1_4_port, O(3) => 
                           res1_3_port, O(2) => res1_2_port, O(1) => 
                           res1_1_port, O(0) => res1_0_port);
   log : logic_N32 port map( A(31) => INA(31), A(30) => n6, A(29) => INA(29), 
                           A(28) => n5, A(27) => INA(27), A(26) => INA(26), 
                           A(25) => n9, A(24) => INA(24), A(23) => INA(23), 
                           A(22) => INA(22), A(21) => n12, A(20) => INA(20), 
                           A(19) => INA(19), A(18) => INA(18), A(17) => INA(17)
                           , A(16) => INA(16), A(15) => INA(15), A(14) => 
                           INA(14), A(13) => n4, A(12) => n8, A(11) => n35, 
                           A(10) => n1, A(9) => INA(9), A(8) => INA(8), A(7) =>
                           INA(7), A(6) => INA(6), A(5) => n38, A(4) => n33, 
                           A(3) => n47, A(2) => n45, A(1) => n39, A(0) => n40, 
                           B(31) => INB(31), B(30) => INB(30), B(29) => INB(29)
                           , B(28) => INB(28), B(27) => INB(27), B(26) => 
                           INB(26), B(25) => INB(25), B(24) => INB(24), B(23) 
                           => INB(23), B(22) => INB(22), B(21) => n15, B(20) =>
                           n13, B(19) => n29, B(18) => n32, B(17) => n30, B(16)
                           => n10, B(15) => n21, B(14) => n18, B(13) => n2, 
                           B(12) => n23, B(11) => n28, B(10) => n25, B(9) => 
                           n20, B(8) => n41, B(7) => n27, B(6) => n42, B(5) => 
                           n22, B(4) => n26, B(3) => n31, B(2) => n44, B(1) => 
                           n19, B(0) => n43, SEL(0) => OP(0), SEL(1) => OP(1), 
                           SEL(2) => OP(2), SEL(3) => OP(3), SEL(4) => OP(4), 
                           O(31) => res2_31_port, O(30) => res2_30_port, O(29) 
                           => res2_29_port, O(28) => res2_28_port, O(27) => 
                           res2_27_port, O(26) => res2_26_port, O(25) => 
                           res2_25_port, O(24) => res2_24_port, O(23) => 
                           res2_23_port, O(22) => res2_22_port, O(21) => 
                           res2_21_port, O(20) => res2_20_port, O(19) => 
                           res2_19_port, O(18) => res2_18_port, O(17) => 
                           res2_17_port, O(16) => res2_16_port, O(15) => 
                           res2_15_port, O(14) => res2_14_port, O(13) => 
                           res2_13_port, O(12) => res2_12_port, O(11) => 
                           res2_11_port, O(10) => res2_10_port, O(9) => 
                           res2_9_port, O(8) => res2_8_port, O(7) => 
                           res2_7_port, O(6) => res2_6_port, O(5) => 
                           res2_5_port, O(4) => res2_4_port, O(3) => 
                           res2_3_port, O(2) => res2_2_port, O(1) => 
                           res2_1_port, O(0) => res2_0_port);
   shifter : SHIFTER_GENERIC_N32 port map( A(31) => INA(31), A(30) => n6, A(29)
                           => INA(29), A(28) => n5, A(27) => INA(27), A(26) => 
                           INA(26), A(25) => n9, A(24) => INA(24), A(23) => 
                           INA(23), A(22) => INA(22), A(21) => n12, A(20) => 
                           INA(20), A(19) => INA(19), A(18) => INA(18), A(17) 
                           => INA(17), A(16) => INA(16), A(15) => INA(15), 
                           A(14) => INA(14), A(13) => n4, A(12) => n8, A(11) =>
                           n35, A(10) => INA(10), A(9) => INA(9), A(8) => 
                           INA(8), A(7) => INA(7), A(6) => INA(6), A(5) => n38,
                           A(4) => n33, A(3) => n47, A(2) => n45, A(1) => n39, 
                           A(0) => n40, B(31) => INB(31), B(30) => INB(30), 
                           B(29) => INB(29), B(28) => INB(28), B(27) => INB(27)
                           , B(26) => INB(26), B(25) => INB(25), B(24) => 
                           INB(24), B(23) => INB(23), B(22) => INB(22), B(21) 
                           => n15, B(20) => n13, B(19) => n29, B(18) => n32, 
                           B(17) => n30, B(16) => n10, B(15) => n21, B(14) => 
                           n18, B(13) => n2, B(12) => n23, B(11) => n28, B(10) 
                           => n25, B(9) => n20, B(8) => INB(8), B(7) => n27, 
                           B(6) => n42, B(5) => n22, B(4) => n26, B(3) => n31, 
                           B(2) => n44, B(1) => n16, B(0) => n37, sel(0) => 
                           OP(0), sel(1) => OP(1), sel(2) => OP(2), sel(3) => 
                           OP(3), sel(4) => OP(4), OUTPUT(31) => res3_31_port, 
                           OUTPUT(30) => res3_30_port, OUTPUT(29) => 
                           res3_29_port, OUTPUT(28) => res3_28_port, OUTPUT(27)
                           => res3_27_port, OUTPUT(26) => res3_26_port, 
                           OUTPUT(25) => res3_25_port, OUTPUT(24) => 
                           res3_24_port, OUTPUT(23) => res3_23_port, OUTPUT(22)
                           => res3_22_port, OUTPUT(21) => res3_21_port, 
                           OUTPUT(20) => res3_20_port, OUTPUT(19) => 
                           res3_19_port, OUTPUT(18) => res3_18_port, OUTPUT(17)
                           => res3_17_port, OUTPUT(16) => res3_16_port, 
                           OUTPUT(15) => res3_15_port, OUTPUT(14) => 
                           res3_14_port, OUTPUT(13) => res3_13_port, OUTPUT(12)
                           => res3_12_port, OUTPUT(11) => res3_11_port, 
                           OUTPUT(10) => res3_10_port, OUTPUT(9) => res3_9_port
                           , OUTPUT(8) => res3_8_port, OUTPUT(7) => res3_7_port
                           , OUTPUT(6) => res3_6_port, OUTPUT(5) => res3_5_port
                           , OUTPUT(4) => res3_4_port, OUTPUT(3) => res3_3_port
                           , OUTPUT(2) => res3_2_port, OUTPUT(1) => res3_1_port
                           , OUTPUT(0) => res3_0_port);
   comp : comparator_N32 port map( inA(31) => INA(31), inA(30) => INA(30), 
                           inA(29) => INA(29), inA(28) => INA(28), inA(27) => 
                           INA(27), inA(26) => INA(26), inA(25) => INA(25), 
                           inA(24) => INA(24), inA(23) => INA(23), inA(22) => 
                           INA(22), inA(21) => INA(21), inA(20) => INA(20), 
                           inA(19) => INA(19), inA(18) => INA(18), inA(17) => 
                           INA(17), inA(16) => INA(16), inA(15) => INA(15), 
                           inA(14) => INA(14), inA(13) => INA(13), inA(12) => 
                           INA(12), inA(11) => INA(11), inA(10) => INA(10), 
                           inA(9) => INA(9), inA(8) => INA(8), inA(7) => INA(7)
                           , inA(6) => INA(6), inA(5) => INA(5), inA(4) => 
                           INA(4), inA(3) => INA(3), inA(2) => INA(2), inA(1) 
                           => INA(1), inA(0) => INA(0), inB(31) => INB(31), 
                           inB(30) => INB(30), inB(29) => INB(29), inB(28) => 
                           INB(28), inB(27) => INB(27), inB(26) => INB(26), 
                           inB(25) => INB(25), inB(24) => INB(24), inB(23) => 
                           INB(23), inB(22) => INB(22), inB(21) => n15, inB(20)
                           => n13, inB(19) => n29, inB(18) => n32, inB(17) => 
                           n30, inB(16) => n10, inB(15) => n21, inB(14) => n18,
                           inB(13) => n2, inB(12) => n23, inB(11) => n28, 
                           inB(10) => n25, inB(9) => n20, inB(8) => n41, inB(7)
                           => n27, inB(6) => n42, inB(5) => n22, inB(4) => n26,
                           inB(3) => n3, inB(2) => n24, inB(1) => n16, inB(0) 
                           => n17, op(0) => OP(0), op(1) => OP(1), op(2) => 
                           OP(2), op(3) => OP(3), op(4) => OP(4), res(31) => 
                           n_1392, res(30) => n_1393, res(29) => n_1394, 
                           res(28) => n_1395, res(27) => n_1396, res(26) => 
                           n_1397, res(25) => n_1398, res(24) => n_1399, 
                           res(23) => n_1400, res(22) => n_1401, res(21) => 
                           n_1402, res(20) => n_1403, res(19) => n_1404, 
                           res(18) => n_1405, res(17) => n_1406, res(16) => 
                           n_1407, res(15) => n_1408, res(14) => n_1409, 
                           res(13) => n_1410, res(12) => n_1411, res(11) => 
                           n_1412, res(10) => n_1413, res(9) => n_1414, res(8) 
                           => n_1415, res(7) => n_1416, res(6) => n_1417, 
                           res(5) => n_1418, res(4) => n_1419, res(3) => n_1420
                           , res(2) => n_1421, res(1) => n_1422, res(0) => 
                           res4_0_port);
   mux : mux4to1_N32 port map( inadd(31) => res1_31_port, inadd(30) => 
                           res1_30_port, inadd(29) => res1_29_port, inadd(28) 
                           => res1_28_port, inadd(27) => res1_27_port, 
                           inadd(26) => res1_26_port, inadd(25) => res1_25_port
                           , inadd(24) => res1_24_port, inadd(23) => 
                           res1_23_port, inadd(22) => res1_22_port, inadd(21) 
                           => res1_21_port, inadd(20) => res1_20_port, 
                           inadd(19) => res1_19_port, inadd(18) => res1_18_port
                           , inadd(17) => res1_17_port, inadd(16) => 
                           res1_16_port, inadd(15) => res1_15_port, inadd(14) 
                           => res1_14_port, inadd(13) => res1_13_port, 
                           inadd(12) => res1_12_port, inadd(11) => res1_11_port
                           , inadd(10) => res1_10_port, inadd(9) => res1_9_port
                           , inadd(8) => res1_8_port, inadd(7) => res1_7_port, 
                           inadd(6) => res1_6_port, inadd(5) => res1_5_port, 
                           inadd(4) => res1_4_port, inadd(3) => res1_3_port, 
                           inadd(2) => res1_2_port, inadd(1) => res1_1_port, 
                           inadd(0) => res1_0_port, inlog(31) => res2_31_port, 
                           inlog(30) => res2_30_port, inlog(29) => res2_29_port
                           , inlog(28) => res2_28_port, inlog(27) => 
                           res2_27_port, inlog(26) => res2_26_port, inlog(25) 
                           => res2_25_port, inlog(24) => res2_24_port, 
                           inlog(23) => res2_23_port, inlog(22) => res2_22_port
                           , inlog(21) => res2_21_port, inlog(20) => 
                           res2_20_port, inlog(19) => res2_19_port, inlog(18) 
                           => res2_18_port, inlog(17) => res2_17_port, 
                           inlog(16) => res2_16_port, inlog(15) => res2_15_port
                           , inlog(14) => res2_14_port, inlog(13) => 
                           res2_13_port, inlog(12) => res2_12_port, inlog(11) 
                           => res2_11_port, inlog(10) => res2_10_port, inlog(9)
                           => res2_9_port, inlog(8) => res2_8_port, inlog(7) =>
                           res2_7_port, inlog(6) => res2_6_port, inlog(5) => 
                           res2_5_port, inlog(4) => res2_4_port, inlog(3) => 
                           res2_3_port, inlog(2) => res2_2_port, inlog(1) => 
                           res2_1_port, inlog(0) => res2_0_port, insh(31) => 
                           res3_31_port, insh(30) => res3_30_port, insh(29) => 
                           res3_29_port, insh(28) => res3_28_port, insh(27) => 
                           res3_27_port, insh(26) => res3_26_port, insh(25) => 
                           res3_25_port, insh(24) => res3_24_port, insh(23) => 
                           res3_23_port, insh(22) => res3_22_port, insh(21) => 
                           res3_21_port, insh(20) => res3_20_port, insh(19) => 
                           res3_19_port, insh(18) => res3_18_port, insh(17) => 
                           res3_17_port, insh(16) => res3_16_port, insh(15) => 
                           res3_15_port, insh(14) => res3_14_port, insh(13) => 
                           res3_13_port, insh(12) => res3_12_port, insh(11) => 
                           res3_11_port, insh(10) => res3_10_port, insh(9) => 
                           res3_9_port, insh(8) => res3_8_port, insh(7) => 
                           res3_7_port, insh(6) => res3_6_port, insh(5) => 
                           res3_5_port, insh(4) => res3_4_port, insh(3) => 
                           res3_3_port, insh(2) => res3_2_port, insh(1) => 
                           res3_1_port, insh(0) => res3_0_port, incom(31) => 
                           res4_31_port, incom(30) => res4_30_port, incom(29) 
                           => res4_29_port, incom(28) => res4_28_port, 
                           incom(27) => res4_27_port, incom(26) => res4_26_port
                           , incom(25) => res4_25_port, incom(24) => 
                           res4_24_port, incom(23) => res4_23_port, incom(22) 
                           => res4_22_port, incom(21) => res4_21_port, 
                           incom(20) => res4_20_port, incom(19) => res4_19_port
                           , incom(18) => res4_18_port, incom(17) => 
                           res4_17_port, incom(16) => res4_16_port, incom(15) 
                           => res4_15_port, incom(14) => res4_14_port, 
                           incom(13) => res4_13_port, incom(12) => res4_12_port
                           , incom(11) => res4_11_port, incom(10) => 
                           res4_10_port, incom(9) => res4_9_port, incom(8) => 
                           res4_8_port, incom(7) => res4_7_port, incom(6) => 
                           res4_6_port, incom(5) => res4_5_port, incom(4) => 
                           res4_4_port, incom(3) => res4_3_port, incom(2) => 
                           res4_2_port, incom(1) => res4_1_port, incom(0) => 
                           res4_0_port, sel(0) => OP(0), sel(1) => OP(1), 
                           sel(2) => OP(2), sel(3) => OP(3), sel(4) => OP(4), 
                           O(31) => alu_out(31), O(30) => alu_out(30), O(29) =>
                           alu_out(29), O(28) => alu_out(28), O(27) => 
                           alu_out(27), O(26) => alu_out(26), O(25) => 
                           alu_out(25), O(24) => alu_out(24), O(23) => 
                           alu_out(23), O(22) => alu_out(22), O(21) => 
                           alu_out(21), O(20) => alu_out(20), O(19) => 
                           alu_out(19), O(18) => alu_out(18), O(17) => 
                           alu_out(17), O(16) => alu_out(16), O(15) => 
                           alu_out(15), O(14) => alu_out(14), O(13) => 
                           alu_out(13), O(12) => alu_out(12), O(11) => 
                           alu_out(11), O(10) => alu_out(10), O(9) => 
                           alu_out(9), O(8) => alu_out(8), O(7) => alu_out(7), 
                           O(6) => alu_out(6), O(5) => alu_out(5), O(4) => 
                           alu_out(4), O(3) => alu_out(3), O(2) => alu_out(2), 
                           O(1) => alu_out(1), O(0) => alu_out(0));
   U1 : BUF_X2 port map( A => INA(1), Z => n39);
   U2 : BUF_X2 port map( A => INA(5), Z => n38);
   U3 : BUF_X1 port map( A => INA(30), Z => n6);
   U4 : BUF_X1 port map( A => INA(4), Z => n33);
   U5 : BUF_X1 port map( A => INA(0), Z => n40);
   U6 : BUF_X1 port map( A => n24, Z => n44);
   U7 : CLKBUF_X2 port map( A => INB(1), Z => n16);
   U8 : CLKBUF_X1 port map( A => INB(4), Z => n26);
   U9 : CLKBUF_X1 port map( A => INA(10), Z => n1);
   U10 : CLKBUF_X1 port map( A => INB(13), Z => n2);
   U11 : CLKBUF_X1 port map( A => INB(3), Z => n3);
   U12 : INV_X2 port map( A => n14, ZN => n37);
   U13 : BUF_X2 port map( A => INA(13), Z => n4);
   U14 : BUF_X2 port map( A => INA(28), Z => n5);
   U15 : INV_X1 port map( A => INA(12), ZN => n7);
   U16 : INV_X2 port map( A => n7, ZN => n8);
   U17 : BUF_X2 port map( A => INA(25), Z => n9);
   U18 : CLKBUF_X1 port map( A => INB(16), Z => n10);
   U19 : INV_X1 port map( A => INA(21), ZN => n11);
   U20 : INV_X2 port map( A => n11, ZN => n12);
   U21 : CLKBUF_X1 port map( A => INB(2), Z => n24);
   U22 : CLKBUF_X1 port map( A => INB(20), Z => n13);
   U23 : CLKBUF_X1 port map( A => n36, Z => n14);
   U24 : CLKBUF_X1 port map( A => INB(21), Z => n15);
   U25 : CLKBUF_X1 port map( A => INB(5), Z => n22);
   U26 : INV_X1 port map( A => n36, ZN => n17);
   U27 : CLKBUF_X1 port map( A => INB(14), Z => n18);
   U28 : CLKBUF_X1 port map( A => n16, Z => n19);
   U29 : CLKBUF_X1 port map( A => INB(9), Z => n20);
   U30 : CLKBUF_X1 port map( A => INB(15), Z => n21);
   U31 : CLKBUF_X1 port map( A => INB(12), Z => n23);
   U32 : CLKBUF_X1 port map( A => INB(10), Z => n25);
   U33 : CLKBUF_X1 port map( A => INB(7), Z => n27);
   U34 : CLKBUF_X1 port map( A => INB(11), Z => n28);
   U35 : CLKBUF_X1 port map( A => INB(19), Z => n29);
   U36 : CLKBUF_X1 port map( A => INB(17), Z => n30);
   U37 : CLKBUF_X1 port map( A => n3, Z => n31);
   U38 : CLKBUF_X1 port map( A => INB(18), Z => n32);
   U39 : INV_X1 port map( A => INA(11), ZN => n34);
   U40 : INV_X2 port map( A => n34, ZN => n35);
   U41 : INV_X1 port map( A => INB(0), ZN => n36);
   U42 : CLKBUF_X1 port map( A => INB(6), Z => n42);
   U43 : CLKBUF_X1 port map( A => INB(8), Z => n41);
   U44 : CLKBUF_X1 port map( A => n37, Z => n43);
   U45 : CLKBUF_X1 port map( A => INA(2), Z => n45);
   U46 : INV_X1 port map( A => INA(3), ZN => n46);
   U47 : INV_X2 port map( A => n46, ZN => n47);
   res4_1_port <= '0';
   res4_2_port <= '0';
   res4_3_port <= '0';
   res4_4_port <= '0';
   res4_5_port <= '0';
   res4_6_port <= '0';
   res4_7_port <= '0';
   res4_8_port <= '0';
   res4_9_port <= '0';
   res4_10_port <= '0';
   res4_11_port <= '0';
   res4_12_port <= '0';
   res4_13_port <= '0';
   res4_14_port <= '0';
   res4_15_port <= '0';
   res4_16_port <= '0';
   res4_17_port <= '0';
   res4_18_port <= '0';
   res4_19_port <= '0';
   res4_20_port <= '0';
   res4_21_port <= '0';
   res4_22_port <= '0';
   res4_23_port <= '0';
   res4_24_port <= '0';
   res4_25_port <= '0';
   res4_26_port <= '0';
   res4_27_port <= '0';
   res4_28_port <= '0';
   res4_29_port <= '0';
   res4_30_port <= '0';
   res4_31_port <= '0';

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity mux_3to1_N32_0 is

   port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux_3to1_N32_0;

architecture SYN_BEHAVIORAL of mux_3to1_N32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n18, n19, n20, 
      n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67 : std_logic;

begin
   
   U1 : CLKBUF_X3 port map( A => n65, Z => n33);
   U2 : OR3_X2 port map( A1 => n28, A2 => n29, A3 => n30, ZN => Y(2));
   U3 : INV_X2 port map( A => n59, ZN => Y(24));
   U4 : NAND3_X2 port map( A1 => n14, A2 => n15, A3 => n16, ZN => Y(26));
   U5 : BUF_X2 port map( A => n65, Z => n32);
   U6 : OR3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => Y(4));
   U7 : INV_X1 port map( A => n51, ZN => Y(16));
   U8 : INV_X1 port map( A => n52, ZN => Y(17));
   U9 : INV_X1 port map( A => n53, ZN => Y(18));
   U10 : INV_X1 port map( A => n50, ZN => Y(15));
   U11 : INV_X1 port map( A => n58, ZN => Y(23));
   U12 : NAND3_X1 port map( A1 => n7, A2 => n8, A3 => n9, ZN => Y(3));
   U13 : BUF_X1 port map( A => n31, Z => n34);
   U14 : BUF_X2 port map( A => n33, Z => n22);
   U15 : OR3_X2 port map( A1 => n4, A2 => n5, A3 => n6, ZN => Y(1));
   U16 : BUF_X2 port map( A => n31, Z => n21);
   U17 : AND2_X1 port map( A1 => B(1), A2 => n66, ZN => n4);
   U18 : AND2_X1 port map( A1 => A(1), A2 => n31, ZN => n5);
   U19 : AND2_X1 port map( A1 => C(1), A2 => n32, ZN => n6);
   U20 : BUF_X2 port map( A => n66, Z => n37);
   U21 : INV_X1 port map( A => n45, ZN => Y(10));
   U22 : NAND2_X1 port map( A1 => B(3), A2 => n36, ZN => n7);
   U23 : NAND2_X1 port map( A1 => A(3), A2 => n21, ZN => n8);
   U24 : NAND2_X1 port map( A1 => C(3), A2 => n33, ZN => n9);
   U25 : INV_X2 port map( A => n44, ZN => Y(9));
   U26 : NAND3_X1 port map( A1 => n10, A2 => n11, A3 => n12, ZN => Y(5));
   U27 : NAND2_X1 port map( A1 => B(5), A2 => n37, ZN => n10);
   U28 : NAND2_X1 port map( A1 => A(5), A2 => n31, ZN => n11);
   U29 : NAND2_X1 port map( A1 => C(5), A2 => n33, ZN => n12);
   U30 : INV_X2 port map( A => n55, ZN => Y(20));
   U31 : CLKBUF_X1 port map( A => n31, Z => n35);
   U32 : INV_X1 port map( A => n48, ZN => Y(13));
   U33 : NAND2_X1 port map( A1 => B(26), A2 => n37, ZN => n14);
   U34 : NAND2_X1 port map( A1 => A(26), A2 => n21, ZN => n15);
   U35 : NAND2_X1 port map( A1 => C(26), A2 => n32, ZN => n16);
   U36 : INV_X1 port map( A => n47, ZN => Y(12));
   U37 : INV_X1 port map( A => n60, ZN => Y(25));
   U38 : INV_X1 port map( A => n56, ZN => Y(21));
   U39 : AND2_X1 port map( A1 => B(4), A2 => n66, ZN => n18);
   U40 : AND2_X1 port map( A1 => A(4), A2 => n31, ZN => n19);
   U41 : AND2_X1 port map( A1 => C(4), A2 => n32, ZN => n20);
   U42 : BUF_X2 port map( A => n66, Z => n36);
   U43 : OR2_X1 port map( A1 => SEL(1), A2 => n38, ZN => n39);
   U44 : INV_X1 port map( A => n46, ZN => Y(11));
   U45 : AND2_X2 port map( A1 => n40, A2 => n39, ZN => n31);
   U46 : INV_X2 port map( A => n49, ZN => Y(14));
   U47 : OR3_X2 port map( A1 => n26, A2 => n27, A3 => n25, ZN => Y(0));
   U48 : AND2_X1 port map( A1 => n66, A2 => B(0), ZN => n25);
   U49 : AND2_X1 port map( A1 => A(0), A2 => n31, ZN => n26);
   U50 : AND2_X1 port map( A1 => C(0), A2 => n33, ZN => n27);
   U51 : AND2_X1 port map( A1 => B(2), A2 => n66, ZN => n28);
   U52 : AND2_X1 port map( A1 => A(2), A2 => n31, ZN => n29);
   U53 : AND2_X1 port map( A1 => C(2), A2 => n33, ZN => n30);
   U54 : INV_X2 port map( A => n61, ZN => Y(27));
   U55 : INV_X2 port map( A => n42, ZN => Y(7));
   U56 : INV_X2 port map( A => n41, ZN => Y(6));
   U57 : INV_X2 port map( A => n57, ZN => Y(22));
   U58 : INV_X2 port map( A => n43, ZN => Y(8));
   U59 : INV_X1 port map( A => n39, ZN => n66);
   U60 : INV_X1 port map( A => SEL(0), ZN => n38);
   U61 : NAND2_X1 port map( A1 => n38, A2 => SEL(1), ZN => n40);
   U62 : INV_X1 port map( A => n40, ZN => n65);
   U63 : AOI222_X1 port map( A1 => B(6), A2 => n36, B1 => A(6), B2 => n31, C1 
                           => C(6), C2 => n33, ZN => n41);
   U64 : AOI222_X1 port map( A1 => B(7), A2 => n37, B1 => A(7), B2 => n35, C1 
                           => C(7), C2 => n32, ZN => n42);
   U65 : AOI222_X1 port map( A1 => B(8), A2 => n36, B1 => A(8), B2 => n31, C1 
                           => C(8), C2 => n32, ZN => n43);
   U66 : AOI222_X1 port map( A1 => B(9), A2 => n36, B1 => A(9), B2 => n21, C1 
                           => C(9), C2 => n32, ZN => n44);
   U67 : AOI222_X1 port map( A1 => B(10), A2 => n36, B1 => A(10), B2 => n21, C1
                           => C(10), C2 => n33, ZN => n45);
   U68 : AOI222_X1 port map( A1 => B(11), A2 => n36, B1 => A(11), B2 => n35, C1
                           => C(11), C2 => n22, ZN => n46);
   U69 : AOI222_X1 port map( A1 => B(12), A2 => n36, B1 => A(12), B2 => n21, C1
                           => C(12), C2 => n32, ZN => n47);
   U70 : AOI222_X1 port map( A1 => B(13), A2 => n37, B1 => A(13), B2 => n34, C1
                           => C(13), C2 => n22, ZN => n48);
   U71 : AOI222_X1 port map( A1 => B(14), A2 => n36, B1 => A(14), B2 => n21, C1
                           => C(14), C2 => n33, ZN => n49);
   U72 : AOI222_X1 port map( A1 => B(15), A2 => n37, B1 => A(15), B2 => n34, C1
                           => C(15), C2 => n22, ZN => n50);
   U73 : AOI222_X1 port map( A1 => B(16), A2 => n37, B1 => A(16), B2 => n35, C1
                           => C(16), C2 => n32, ZN => n51);
   U74 : AOI222_X1 port map( A1 => B(17), A2 => n36, B1 => A(17), B2 => n21, C1
                           => C(17), C2 => n22, ZN => n52);
   U75 : AOI222_X1 port map( A1 => B(18), A2 => n36, B1 => A(18), B2 => n34, C1
                           => C(18), C2 => n22, ZN => n53);
   U76 : AOI222_X1 port map( A1 => B(19), A2 => n36, B1 => A(19), B2 => n35, C1
                           => C(19), C2 => n33, ZN => n54);
   U77 : INV_X1 port map( A => n54, ZN => Y(19));
   U78 : AOI222_X1 port map( A1 => B(20), A2 => n37, B1 => A(20), B2 => n21, C1
                           => C(20), C2 => n22, ZN => n55);
   U79 : AOI222_X1 port map( A1 => B(21), A2 => n37, B1 => A(21), B2 => n21, C1
                           => C(21), C2 => n22, ZN => n56);
   U80 : AOI222_X1 port map( A1 => B(22), A2 => n36, B1 => A(22), B2 => n21, C1
                           => C(22), C2 => n32, ZN => n57);
   U81 : AOI222_X1 port map( A1 => B(23), A2 => n36, B1 => A(23), B2 => n34, C1
                           => C(23), C2 => n32, ZN => n58);
   U82 : AOI222_X1 port map( A1 => B(24), A2 => n36, B1 => A(24), B2 => n31, C1
                           => C(24), C2 => n22, ZN => n59);
   U83 : AOI222_X1 port map( A1 => B(25), A2 => n37, B1 => A(25), B2 => n35, C1
                           => C(25), C2 => n32, ZN => n60);
   U84 : AOI222_X1 port map( A1 => B(27), A2 => n37, B1 => A(27), B2 => n21, C1
                           => C(27), C2 => n22, ZN => n61);
   U85 : AOI222_X1 port map( A1 => B(28), A2 => n36, B1 => A(28), B2 => n21, C1
                           => C(28), C2 => n32, ZN => n62);
   U86 : INV_X1 port map( A => n62, ZN => Y(28));
   U87 : AOI222_X1 port map( A1 => B(29), A2 => n37, B1 => A(29), B2 => n21, C1
                           => C(29), C2 => n33, ZN => n63);
   U88 : INV_X1 port map( A => n63, ZN => Y(29));
   U89 : AOI222_X1 port map( A1 => B(30), A2 => n36, B1 => A(30), B2 => n34, C1
                           => C(30), C2 => n32, ZN => n64);
   U90 : INV_X1 port map( A => n64, ZN => Y(30));
   U91 : AOI222_X1 port map( A1 => B(31), A2 => n36, B1 => A(31), B2 => n34, C1
                           => C(31), C2 => n22, ZN => n67);
   U92 : INV_X1 port map( A => n67, ZN => Y(31));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity FWD_UNIT is

   port( Rst : in std_logic;  Rs1, Rs2, Rd_M, Rd_W : in std_logic_vector (4 
         downto 0);  ICODE, ICODE_M, ICODE_W : in std_logic_vector (5 downto 0)
         ;  SEL_A, SEL_B : out std_logic_vector (1 downto 0));

end FWD_UNIT;

architecture SYN_Behavioral of FWD_UNIT is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FWD_CAM_0
      port( RST : in std_logic;  DATA_IN_1, DATA_IN_2, DATA_IN_3 : in 
            std_logic_vector (5 downto 0);  MATCH_1, MATCH_2, MATCH_3 : out 
            std_logic);
   end component;
   
   signal match_op, match_op_M, match_op_W, net28103, net28106, net28110, 
      net28111, net28112, net28113, net28115, net28123, net28125, net28127, 
      net28128, net28129, net28130, net28133, net28136, net28142, net28165, 
      net28166, net28167, net28170, net29934, net35871, net37653, net35872, 
      net28154, net28152, net28150, net28148, net28137, net28135, net28117, 
      net28105, net28169, net28168, net28138, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54 : std_logic;

begin
   
   CAM : FWD_CAM_0 port map( RST => Rst, DATA_IN_1(5) => ICODE(5), DATA_IN_1(4)
                           => ICODE(4), DATA_IN_1(3) => ICODE(3), DATA_IN_1(2) 
                           => ICODE(2), DATA_IN_1(1) => ICODE(1), DATA_IN_1(0) 
                           => ICODE(0), DATA_IN_2(5) => ICODE_M(5), 
                           DATA_IN_2(4) => ICODE_M(4), DATA_IN_2(3) => 
                           ICODE_M(3), DATA_IN_2(2) => ICODE_M(2), DATA_IN_2(1)
                           => ICODE_M(1), DATA_IN_2(0) => ICODE_M(0), 
                           DATA_IN_3(5) => ICODE_W(5), DATA_IN_3(4) => 
                           ICODE_W(4), DATA_IN_3(3) => ICODE_W(3), DATA_IN_3(2)
                           => ICODE_W(2), DATA_IN_3(1) => ICODE_W(1), 
                           DATA_IN_3(0) => ICODE_W(0), MATCH_1 => match_op, 
                           MATCH_2 => match_op_M, MATCH_3 => match_op_W);
   U2 : OR2_X1 port map( A1 => n23, A2 => net35871, ZN => n1);
   U3 : AND2_X1 port map( A1 => net28166, A2 => net28165, ZN => n2);
   U4 : AND2_X1 port map( A1 => n46, A2 => n45, ZN => n3);
   U5 : OR2_X1 port map( A1 => n1, A2 => n47, ZN => n4);
   U6 : NOR2_X1 port map( A1 => n6, A2 => net28138, ZN => SEL_B(1));
   U7 : NAND4_X1 port map( A1 => n10, A2 => n11, A3 => n12, A4 => n13, ZN => 
                           net28138);
   U8 : XOR2_X1 port map( A => n14, B => Rd_W(2), Z => n13);
   U9 : INV_X1 port map( A => Rs2(2), ZN => n14);
   U10 : XOR2_X1 port map( A => n15, B => Rd_W(3), Z => n12);
   U11 : INV_X1 port map( A => Rs2(3), ZN => n15);
   U12 : XOR2_X1 port map( A => n16, B => Rd_W(1), Z => n11);
   U13 : INV_X1 port map( A => Rs2(1), ZN => n16);
   U14 : XOR2_X1 port map( A => n16, B => Rd_M(1), Z => net28166);
   U15 : XOR2_X1 port map( A => n17, B => Rd_W(4), Z => n10);
   U16 : INV_X1 port map( A => Rs2(4), ZN => n17);
   U17 : NAND3_X1 port map( A1 => n5, A2 => n8, A3 => n19, ZN => n6);
   U18 : AND2_X1 port map( A1 => net28105, A2 => n7, ZN => n19);
   U19 : XOR2_X1 port map( A => n9, B => Rd_W(0), Z => n7);
   U20 : INV_X1 port map( A => Rs2(0), ZN => n9);
   U21 : XOR2_X1 port map( A => n9, B => Rd_M(0), Z => net28165);
   U22 : NOR3_X1 port map( A1 => net35872, A2 => n18, A3 => net28106, ZN => n8)
                           ;
   U23 : INV_X1 port map( A => Rst, ZN => n18);
   U24 : NOR4_X1 port map( A1 => net28129, A2 => net28130, A3 => net35871, A4 
                           => n18, ZN => net28127);
   U25 : NOR4_X1 port map( A1 => net28168, A2 => net28169, A3 => net28170, A4 
                           => n18, ZN => net28167);
   U26 : OR2_X1 port map( A1 => match_op_W, A2 => net28142, ZN => n5);
   U27 : XOR2_X1 port map( A => Rs1(2), B => Rd_W(2), Z => net28111);
   U28 : NOR3_X1 port map( A1 => Rd_W(2), A2 => Rd_W(1), A3 => Rd_W(0), ZN => 
                           net28148);
   U29 : XOR2_X1 port map( A => net28137, B => Rd_W(2), Z => net28150);
   U30 : XOR2_X1 port map( A => Rd_M(2), B => Rs2(2), Z => net28169);
   U31 : INV_X1 port map( A => Rd_W(3), ZN => net28115);
   U32 : XOR2_X1 port map( A => Rd_W(3), B => Rd_M(3), Z => net28154);
   U33 : XOR2_X1 port map( A => Rd_M(3), B => Rs2(3), Z => net28168);
   U34 : XNOR2_X1 port map( A => Rd_W(1), B => Rs1(1), ZN => net28113);
   U35 : XOR2_X1 port map( A => Rd_W(1), B => Rd_M(1), Z => net28152);
   U36 : NAND3_X1 port map( A1 => n21, A2 => net28150, A3 => n20, ZN => 
                           net28105);
   U37 : XOR2_X1 port map( A => net28135, B => Rd_W(0), Z => n20);
   U38 : INV_X1 port map( A => Rd_M(0), ZN => net28135);
   U39 : XOR2_X1 port map( A => net28135, B => Rs1(0), Z => net28123);
   U40 : INV_X1 port map( A => Rd_M(2), ZN => net28137);
   U41 : NOR3_X1 port map( A1 => net28152, A2 => net28154, A3 => n22, ZN => n21
                           );
   U42 : XOR2_X1 port map( A => Rd_W(4), B => Rd_M(4), Z => n22);
   U43 : XOR2_X1 port map( A => Rs1(0), B => Rd_W(0), Z => net28110);
   U44 : AND3_X1 port map( A1 => net28115, A2 => net28117, A3 => net28148, ZN 
                           => net35872);
   U45 : OR2_X1 port map( A1 => net28103, A2 => net35872, ZN => net37653);
   U46 : INV_X1 port map( A => Rd_W(4), ZN => net28117);
   U47 : XOR2_X1 port map( A => net28117, B => Rs1(4), Z => net28112);
   U48 : NAND3_X1 port map( A1 => n26, A2 => net28127, A3 => n3, ZN => n44);
   U49 : INV_X1 port map( A => n23, ZN => n46);
   U50 : NOR3_X1 port map( A1 => n53, A2 => net37653, A3 => n54, ZN => SEL_A(1)
                           );
   U51 : XOR2_X1 port map( A => Rd_M(2), B => Rs1(2), Z => n23);
   U52 : OAI21_X1 port map( B1 => match_op_M, B2 => n34, A => n33, ZN => n24);
   U53 : NOR2_X1 port map( A1 => n48, A2 => n4, ZN => n54);
   U54 : CLKBUF_X1 port map( A => ICODE_W(0), Z => n25);
   U55 : OR2_X1 port map( A1 => net28128, A2 => match_op, ZN => n26);
   U56 : NAND3_X1 port map( A1 => net28128, A2 => net28167, A3 => n2, ZN => n39
                           );
   U57 : NOR4_X2 port map( A1 => n31, A2 => n30, A3 => ICODE_M(4), A4 => 
                           ICODE_M(5), ZN => n34);
   U58 : CLKBUF_X1 port map( A => ICODE_W(1), Z => n27);
   U59 : OAI21_X1 port map( B1 => match_op_M, B2 => n34, A => n33, ZN => n28);
   U60 : OAI21_X1 port map( B1 => n34, B2 => match_op_M, A => n33, ZN => n48);
   U61 : XNOR2_X1 port map( A => Rd_M(1), B => Rs1(1), ZN => net28125);
   U62 : OR3_X1 port map( A1 => ICODE_M(1), A2 => ICODE_M(2), A3 => ICODE_M(0),
                           ZN => n31);
   U63 : XNOR2_X1 port map( A => net28133, B => Rs1(4), ZN => net35871);
   U64 : OR2_X1 port map( A1 => match_op, A2 => net28128, ZN => n51);
   U65 : OR2_X1 port map( A1 => net28142, A2 => match_op_W, ZN => net29934);
   U66 : CLKBUF_X1 port map( A => ICODE_W(3), Z => n29);
   U67 : CLKBUF_X1 port map( A => ICODE_M(3), Z => n30);
   U68 : INV_X1 port map( A => Rd_M(4), ZN => net28133);
   U69 : INV_X1 port map( A => Rd_M(3), ZN => net28136);
   U70 : NOR3_X1 port map( A1 => Rd_M(2), A2 => Rd_M(0), A3 => Rd_M(1), ZN => 
                           n32);
   U71 : NAND3_X1 port map( A1 => net28133, A2 => net28136, A3 => n32, ZN => 
                           n33);
   U72 : INV_X1 port map( A => ICODE(0), ZN => n38);
   U73 : INV_X1 port map( A => ICODE(1), ZN => n37);
   U74 : INV_X1 port map( A => ICODE(2), ZN => n36);
   U75 : NOR3_X1 port map( A1 => ICODE(5), A2 => ICODE(4), A3 => ICODE(3), ZN 
                           => n35);
   U76 : NAND4_X1 port map( A1 => n38, A2 => n37, A3 => n36, A4 => n35, ZN => 
                           net28106);
   U77 : INV_X1 port map( A => net28106, ZN => net28128);
   U78 : XOR2_X1 port map( A => Rd_M(4), B => Rs2(4), Z => net28170);
   U79 : NOR2_X1 port map( A1 => n28, A2 => n39, ZN => SEL_B(0));
   U80 : INV_X1 port map( A => ICODE_W(2), ZN => n42);
   U81 : INV_X1 port map( A => n27, ZN => n41);
   U82 : INV_X1 port map( A => n25, ZN => n40);
   U83 : NAND3_X1 port map( A1 => n42, A2 => n41, A3 => n40, ZN => n43);
   U84 : NOR4_X1 port map( A1 => n43, A2 => n29, A3 => ICODE_W(4), A4 => 
                           ICODE_W(5), ZN => net28142);
   U85 : XOR2_X1 port map( A => net28136, B => Rs1(3), Z => n45);
   U86 : INV_X1 port map( A => net28123, ZN => net28129);
   U87 : INV_X1 port map( A => net28125, ZN => net28130);
   U88 : NOR2_X1 port map( A1 => n44, A2 => n24, ZN => SEL_A(0));
   U89 : NAND3_X1 port map( A1 => net28123, A2 => n45, A3 => net28125, ZN => 
                           n47);
   U90 : XOR2_X1 port map( A => net28115, B => Rs1(3), Z => n49);
   U91 : NAND4_X1 port map( A1 => Rst, A2 => net28112, A3 => net28113, A4 => 
                           n49, ZN => n50);
   U92 : NOR3_X1 port map( A1 => n50, A2 => net28110, A3 => net28111, ZN => n52
                           );
   U93 : OAI211_X1 port map( C1 => net28105, C2 => net28106, A => n51, B => n52
                           , ZN => n53);
   U94 : INV_X1 port map( A => net29934, ZN => net28103);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity ID_EX is

   port( CLK, RST : in std_logic;  NPC_IN, NPC_L_IN, A_IN, B_IN, IMM_IN : in 
         std_logic_vector (31 downto 0);  RS1_IN, RS2_IN, RD_IN : in 
         std_logic_vector (4 downto 0);  OPCODE_IN : in std_logic_vector (5 
         downto 0);  IR_IN : in std_logic_vector (15 downto 0);  PR_IN : in 
         std_logic;  NPC_OUT, NPC_L_OUT, A_OUT, B_OUT, IMM_OUT : out 
         std_logic_vector (31 downto 0);  RS1_OUT, RS2_OUT, RD_OUT : out 
         std_logic_vector (4 downto 0);  OPCODE_OUT : out std_logic_vector (5 
         downto 0);  IR_OUT : out std_logic_vector (15 downto 0);  PR_OUT : out
         std_logic);

end ID_EX;

architecture SYN_Behavioral of ID_EX is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620 : std_logic;

begin
   
   PR_OUT_reg : DFFR_X1 port map( D => PR_IN, CK => CLK, RN => n7, Q => PR_OUT,
                           QN => n_1423);
   A_OUT_reg_31_inst : DFFR_X1 port map( D => A_IN(31), CK => CLK, RN => n7, Q 
                           => A_OUT(31), QN => n_1424);
   A_OUT_reg_30_inst : DFFR_X1 port map( D => A_IN(30), CK => CLK, RN => n7, Q 
                           => A_OUT(30), QN => n_1425);
   A_OUT_reg_29_inst : DFFR_X1 port map( D => A_IN(29), CK => CLK, RN => n7, Q 
                           => A_OUT(29), QN => n_1426);
   A_OUT_reg_28_inst : DFFR_X1 port map( D => A_IN(28), CK => CLK, RN => n7, Q 
                           => A_OUT(28), QN => n_1427);
   A_OUT_reg_27_inst : DFFR_X1 port map( D => A_IN(27), CK => CLK, RN => n7, Q 
                           => A_OUT(27), QN => n_1428);
   A_OUT_reg_26_inst : DFFR_X1 port map( D => A_IN(26), CK => CLK, RN => n7, Q 
                           => A_OUT(26), QN => n_1429);
   A_OUT_reg_25_inst : DFFR_X1 port map( D => A_IN(25), CK => CLK, RN => n7, Q 
                           => A_OUT(25), QN => n_1430);
   A_OUT_reg_24_inst : DFFR_X1 port map( D => A_IN(24), CK => CLK, RN => n7, Q 
                           => A_OUT(24), QN => n_1431);
   A_OUT_reg_23_inst : DFFR_X1 port map( D => A_IN(23), CK => CLK, RN => n7, Q 
                           => A_OUT(23), QN => n_1432);
   A_OUT_reg_22_inst : DFFR_X1 port map( D => A_IN(22), CK => CLK, RN => n7, Q 
                           => A_OUT(22), QN => n_1433);
   A_OUT_reg_21_inst : DFFR_X1 port map( D => A_IN(21), CK => CLK, RN => n7, Q 
                           => A_OUT(21), QN => n_1434);
   A_OUT_reg_20_inst : DFFR_X1 port map( D => A_IN(20), CK => CLK, RN => n8, Q 
                           => A_OUT(20), QN => n_1435);
   A_OUT_reg_19_inst : DFFR_X1 port map( D => A_IN(19), CK => CLK, RN => n8, Q 
                           => A_OUT(19), QN => n_1436);
   A_OUT_reg_18_inst : DFFR_X1 port map( D => A_IN(18), CK => CLK, RN => n8, Q 
                           => A_OUT(18), QN => n_1437);
   A_OUT_reg_17_inst : DFFR_X1 port map( D => A_IN(17), CK => CLK, RN => n8, Q 
                           => A_OUT(17), QN => n_1438);
   A_OUT_reg_16_inst : DFFR_X1 port map( D => A_IN(16), CK => CLK, RN => n8, Q 
                           => A_OUT(16), QN => n_1439);
   A_OUT_reg_15_inst : DFFR_X1 port map( D => A_IN(15), CK => CLK, RN => n8, Q 
                           => A_OUT(15), QN => n_1440);
   A_OUT_reg_14_inst : DFFR_X1 port map( D => A_IN(14), CK => CLK, RN => n8, Q 
                           => A_OUT(14), QN => n_1441);
   A_OUT_reg_13_inst : DFFR_X1 port map( D => A_IN(13), CK => CLK, RN => n8, Q 
                           => A_OUT(13), QN => n_1442);
   A_OUT_reg_12_inst : DFFR_X1 port map( D => A_IN(12), CK => CLK, RN => n8, Q 
                           => A_OUT(12), QN => n_1443);
   A_OUT_reg_11_inst : DFFR_X1 port map( D => A_IN(11), CK => CLK, RN => n8, Q 
                           => A_OUT(11), QN => n_1444);
   A_OUT_reg_10_inst : DFFR_X1 port map( D => A_IN(10), CK => CLK, RN => n8, Q 
                           => A_OUT(10), QN => n_1445);
   A_OUT_reg_9_inst : DFFR_X1 port map( D => A_IN(9), CK => CLK, RN => n8, Q =>
                           A_OUT(9), QN => n_1446);
   A_OUT_reg_8_inst : DFFR_X1 port map( D => A_IN(8), CK => CLK, RN => n9, Q =>
                           A_OUT(8), QN => n_1447);
   A_OUT_reg_7_inst : DFFR_X1 port map( D => A_IN(7), CK => CLK, RN => n9, Q =>
                           A_OUT(7), QN => n_1448);
   A_OUT_reg_6_inst : DFFR_X1 port map( D => A_IN(6), CK => CLK, RN => n9, Q =>
                           A_OUT(6), QN => n_1449);
   A_OUT_reg_5_inst : DFFR_X1 port map( D => A_IN(5), CK => CLK, RN => n9, Q =>
                           A_OUT(5), QN => n_1450);
   A_OUT_reg_4_inst : DFFR_X1 port map( D => A_IN(4), CK => CLK, RN => n9, Q =>
                           A_OUT(4), QN => n_1451);
   A_OUT_reg_3_inst : DFFR_X1 port map( D => A_IN(3), CK => CLK, RN => n9, Q =>
                           A_OUT(3), QN => n_1452);
   A_OUT_reg_2_inst : DFFR_X1 port map( D => A_IN(2), CK => CLK, RN => n9, Q =>
                           A_OUT(2), QN => n_1453);
   A_OUT_reg_1_inst : DFFR_X1 port map( D => A_IN(1), CK => CLK, RN => n9, Q =>
                           A_OUT(1), QN => n_1454);
   A_OUT_reg_0_inst : DFFR_X1 port map( D => A_IN(0), CK => CLK, RN => n9, Q =>
                           A_OUT(0), QN => n_1455);
   B_OUT_reg_31_inst : DFFR_X1 port map( D => B_IN(31), CK => CLK, RN => n9, Q 
                           => B_OUT(31), QN => n_1456);
   B_OUT_reg_30_inst : DFFR_X1 port map( D => B_IN(30), CK => CLK, RN => n9, Q 
                           => B_OUT(30), QN => n_1457);
   B_OUT_reg_29_inst : DFFR_X1 port map( D => B_IN(29), CK => CLK, RN => n9, Q 
                           => B_OUT(29), QN => n_1458);
   B_OUT_reg_28_inst : DFFR_X1 port map( D => B_IN(28), CK => CLK, RN => n10, Q
                           => B_OUT(28), QN => n_1459);
   B_OUT_reg_27_inst : DFFR_X1 port map( D => B_IN(27), CK => CLK, RN => n10, Q
                           => B_OUT(27), QN => n_1460);
   B_OUT_reg_26_inst : DFFR_X1 port map( D => B_IN(26), CK => CLK, RN => n10, Q
                           => B_OUT(26), QN => n_1461);
   B_OUT_reg_25_inst : DFFR_X1 port map( D => B_IN(25), CK => CLK, RN => n10, Q
                           => B_OUT(25), QN => n_1462);
   B_OUT_reg_24_inst : DFFR_X1 port map( D => B_IN(24), CK => CLK, RN => n10, Q
                           => B_OUT(24), QN => n_1463);
   B_OUT_reg_23_inst : DFFR_X1 port map( D => B_IN(23), CK => CLK, RN => n10, Q
                           => B_OUT(23), QN => n_1464);
   B_OUT_reg_22_inst : DFFR_X1 port map( D => B_IN(22), CK => CLK, RN => n10, Q
                           => B_OUT(22), QN => n_1465);
   B_OUT_reg_21_inst : DFFR_X1 port map( D => B_IN(21), CK => CLK, RN => n10, Q
                           => B_OUT(21), QN => n_1466);
   B_OUT_reg_20_inst : DFFR_X1 port map( D => B_IN(20), CK => CLK, RN => n10, Q
                           => B_OUT(20), QN => n_1467);
   B_OUT_reg_19_inst : DFFR_X1 port map( D => B_IN(19), CK => CLK, RN => n10, Q
                           => B_OUT(19), QN => n_1468);
   B_OUT_reg_18_inst : DFFR_X1 port map( D => B_IN(18), CK => CLK, RN => n10, Q
                           => B_OUT(18), QN => n_1469);
   B_OUT_reg_17_inst : DFFR_X1 port map( D => B_IN(17), CK => CLK, RN => n10, Q
                           => B_OUT(17), QN => n_1470);
   B_OUT_reg_16_inst : DFFR_X1 port map( D => B_IN(16), CK => CLK, RN => n11, Q
                           => B_OUT(16), QN => n_1471);
   B_OUT_reg_15_inst : DFFR_X1 port map( D => B_IN(15), CK => CLK, RN => n11, Q
                           => B_OUT(15), QN => n_1472);
   B_OUT_reg_14_inst : DFFR_X1 port map( D => B_IN(14), CK => CLK, RN => n11, Q
                           => B_OUT(14), QN => n_1473);
   B_OUT_reg_13_inst : DFFR_X1 port map( D => B_IN(13), CK => CLK, RN => n11, Q
                           => B_OUT(13), QN => n_1474);
   B_OUT_reg_12_inst : DFFR_X1 port map( D => B_IN(12), CK => CLK, RN => n11, Q
                           => B_OUT(12), QN => n_1475);
   B_OUT_reg_11_inst : DFFR_X1 port map( D => B_IN(11), CK => CLK, RN => n11, Q
                           => B_OUT(11), QN => n_1476);
   B_OUT_reg_10_inst : DFFR_X1 port map( D => B_IN(10), CK => CLK, RN => n11, Q
                           => B_OUT(10), QN => n_1477);
   B_OUT_reg_9_inst : DFFR_X1 port map( D => B_IN(9), CK => CLK, RN => n11, Q 
                           => B_OUT(9), QN => n_1478);
   B_OUT_reg_8_inst : DFFR_X1 port map( D => B_IN(8), CK => CLK, RN => n11, Q 
                           => B_OUT(8), QN => n_1479);
   B_OUT_reg_7_inst : DFFR_X1 port map( D => B_IN(7), CK => CLK, RN => n11, Q 
                           => B_OUT(7), QN => n_1480);
   B_OUT_reg_6_inst : DFFR_X1 port map( D => B_IN(6), CK => CLK, RN => n11, Q 
                           => B_OUT(6), QN => n_1481);
   B_OUT_reg_5_inst : DFFR_X1 port map( D => B_IN(5), CK => CLK, RN => n11, Q 
                           => B_OUT(5), QN => n_1482);
   B_OUT_reg_4_inst : DFFR_X1 port map( D => B_IN(4), CK => CLK, RN => n12, Q 
                           => B_OUT(4), QN => n_1483);
   B_OUT_reg_3_inst : DFFR_X1 port map( D => B_IN(3), CK => CLK, RN => n12, Q 
                           => B_OUT(3), QN => n_1484);
   B_OUT_reg_2_inst : DFFR_X1 port map( D => B_IN(2), CK => CLK, RN => n12, Q 
                           => B_OUT(2), QN => n_1485);
   B_OUT_reg_1_inst : DFFR_X1 port map( D => B_IN(1), CK => CLK, RN => n12, Q 
                           => B_OUT(1), QN => n_1486);
   B_OUT_reg_0_inst : DFFR_X1 port map( D => B_IN(0), CK => CLK, RN => n12, Q 
                           => B_OUT(0), QN => n_1487);
   IMM_OUT_reg_31_inst : DFFR_X1 port map( D => IMM_IN(31), CK => CLK, RN => 
                           n12, Q => IMM_OUT(31), QN => n_1488);
   IMM_OUT_reg_30_inst : DFFR_X1 port map( D => IMM_IN(30), CK => CLK, RN => 
                           n12, Q => IMM_OUT(30), QN => n_1489);
   IMM_OUT_reg_29_inst : DFFR_X1 port map( D => IMM_IN(29), CK => CLK, RN => 
                           n12, Q => IMM_OUT(29), QN => n_1490);
   IMM_OUT_reg_28_inst : DFFR_X1 port map( D => IMM_IN(28), CK => CLK, RN => 
                           n12, Q => IMM_OUT(28), QN => n_1491);
   IMM_OUT_reg_27_inst : DFFR_X1 port map( D => IMM_IN(27), CK => CLK, RN => 
                           n12, Q => IMM_OUT(27), QN => n_1492);
   IMM_OUT_reg_26_inst : DFFR_X1 port map( D => IMM_IN(26), CK => CLK, RN => 
                           n12, Q => IMM_OUT(26), QN => n_1493);
   IMM_OUT_reg_25_inst : DFFR_X1 port map( D => IMM_IN(25), CK => CLK, RN => 
                           n12, Q => IMM_OUT(25), QN => n_1494);
   IMM_OUT_reg_24_inst : DFFR_X1 port map( D => IMM_IN(24), CK => CLK, RN => 
                           n13, Q => IMM_OUT(24), QN => n_1495);
   IMM_OUT_reg_23_inst : DFFR_X1 port map( D => IMM_IN(23), CK => CLK, RN => 
                           n13, Q => IMM_OUT(23), QN => n_1496);
   IMM_OUT_reg_22_inst : DFFR_X1 port map( D => IMM_IN(22), CK => CLK, RN => 
                           n13, Q => IMM_OUT(22), QN => n_1497);
   IMM_OUT_reg_21_inst : DFFR_X1 port map( D => IMM_IN(21), CK => CLK, RN => 
                           n13, Q => IMM_OUT(21), QN => n_1498);
   IMM_OUT_reg_20_inst : DFFR_X1 port map( D => IMM_IN(20), CK => CLK, RN => 
                           n13, Q => IMM_OUT(20), QN => n_1499);
   IMM_OUT_reg_19_inst : DFFR_X1 port map( D => IMM_IN(19), CK => CLK, RN => 
                           n13, Q => IMM_OUT(19), QN => n_1500);
   IMM_OUT_reg_18_inst : DFFR_X1 port map( D => IMM_IN(18), CK => CLK, RN => 
                           n13, Q => IMM_OUT(18), QN => n_1501);
   IMM_OUT_reg_17_inst : DFFR_X1 port map( D => IMM_IN(17), CK => CLK, RN => 
                           n13, Q => IMM_OUT(17), QN => n_1502);
   IMM_OUT_reg_16_inst : DFFR_X1 port map( D => IMM_IN(16), CK => CLK, RN => 
                           n13, Q => IMM_OUT(16), QN => n_1503);
   IMM_OUT_reg_15_inst : DFFR_X1 port map( D => IMM_IN(15), CK => CLK, RN => 
                           n13, Q => IMM_OUT(15), QN => n_1504);
   IMM_OUT_reg_14_inst : DFFR_X1 port map( D => IMM_IN(14), CK => CLK, RN => 
                           n13, Q => IMM_OUT(14), QN => n_1505);
   IMM_OUT_reg_13_inst : DFFR_X1 port map( D => IMM_IN(13), CK => CLK, RN => 
                           n13, Q => IMM_OUT(13), QN => n_1506);
   IMM_OUT_reg_12_inst : DFFR_X1 port map( D => IMM_IN(12), CK => CLK, RN => 
                           n14, Q => IMM_OUT(12), QN => n_1507);
   IMM_OUT_reg_11_inst : DFFR_X1 port map( D => IMM_IN(11), CK => CLK, RN => 
                           n14, Q => IMM_OUT(11), QN => n_1508);
   IMM_OUT_reg_10_inst : DFFR_X1 port map( D => IMM_IN(10), CK => CLK, RN => 
                           n14, Q => IMM_OUT(10), QN => n_1509);
   IMM_OUT_reg_9_inst : DFFR_X1 port map( D => IMM_IN(9), CK => CLK, RN => n14,
                           Q => IMM_OUT(9), QN => n_1510);
   IMM_OUT_reg_8_inst : DFFR_X1 port map( D => IMM_IN(8), CK => CLK, RN => n14,
                           Q => IMM_OUT(8), QN => n_1511);
   IMM_OUT_reg_7_inst : DFFR_X1 port map( D => IMM_IN(7), CK => CLK, RN => n14,
                           Q => IMM_OUT(7), QN => n_1512);
   IMM_OUT_reg_6_inst : DFFR_X1 port map( D => IMM_IN(6), CK => CLK, RN => n14,
                           Q => IMM_OUT(6), QN => n_1513);
   IMM_OUT_reg_5_inst : DFFR_X1 port map( D => IMM_IN(5), CK => CLK, RN => n14,
                           Q => IMM_OUT(5), QN => n_1514);
   IMM_OUT_reg_4_inst : DFFR_X1 port map( D => IMM_IN(4), CK => CLK, RN => n14,
                           Q => IMM_OUT(4), QN => n_1515);
   IMM_OUT_reg_3_inst : DFFR_X1 port map( D => IMM_IN(3), CK => CLK, RN => n14,
                           Q => IMM_OUT(3), QN => n_1516);
   IMM_OUT_reg_2_inst : DFFR_X1 port map( D => IMM_IN(2), CK => CLK, RN => n14,
                           Q => IMM_OUT(2), QN => n_1517);
   IMM_OUT_reg_1_inst : DFFR_X1 port map( D => IMM_IN(1), CK => CLK, RN => n14,
                           Q => IMM_OUT(1), QN => n_1518);
   IMM_OUT_reg_0_inst : DFFR_X1 port map( D => IMM_IN(0), CK => CLK, RN => n15,
                           Q => IMM_OUT(0), QN => n_1519);
   NPC_OUT_reg_31_inst : DFFR_X1 port map( D => NPC_IN(31), CK => CLK, RN => 
                           n15, Q => NPC_OUT(31), QN => n_1520);
   NPC_OUT_reg_30_inst : DFFR_X1 port map( D => NPC_IN(30), CK => CLK, RN => 
                           n15, Q => NPC_OUT(30), QN => n_1521);
   NPC_OUT_reg_29_inst : DFFR_X1 port map( D => NPC_IN(29), CK => CLK, RN => 
                           n15, Q => NPC_OUT(29), QN => n_1522);
   NPC_OUT_reg_28_inst : DFFR_X1 port map( D => NPC_IN(28), CK => CLK, RN => 
                           n15, Q => NPC_OUT(28), QN => n_1523);
   NPC_OUT_reg_27_inst : DFFR_X1 port map( D => NPC_IN(27), CK => CLK, RN => 
                           n15, Q => NPC_OUT(27), QN => n_1524);
   NPC_OUT_reg_26_inst : DFFR_X1 port map( D => NPC_IN(26), CK => CLK, RN => 
                           n15, Q => NPC_OUT(26), QN => n_1525);
   NPC_OUT_reg_25_inst : DFFR_X1 port map( D => NPC_IN(25), CK => CLK, RN => 
                           n15, Q => NPC_OUT(25), QN => n_1526);
   NPC_OUT_reg_24_inst : DFFR_X1 port map( D => NPC_IN(24), CK => CLK, RN => 
                           n15, Q => NPC_OUT(24), QN => n_1527);
   NPC_OUT_reg_23_inst : DFFR_X1 port map( D => NPC_IN(23), CK => CLK, RN => 
                           n15, Q => NPC_OUT(23), QN => n_1528);
   NPC_OUT_reg_22_inst : DFFR_X1 port map( D => NPC_IN(22), CK => CLK, RN => 
                           n15, Q => NPC_OUT(22), QN => n_1529);
   NPC_OUT_reg_21_inst : DFFR_X1 port map( D => NPC_IN(21), CK => CLK, RN => 
                           n15, Q => NPC_OUT(21), QN => n_1530);
   NPC_OUT_reg_20_inst : DFFR_X1 port map( D => NPC_IN(20), CK => CLK, RN => 
                           n16, Q => NPC_OUT(20), QN => n_1531);
   NPC_OUT_reg_19_inst : DFFR_X1 port map( D => NPC_IN(19), CK => CLK, RN => 
                           n16, Q => NPC_OUT(19), QN => n_1532);
   NPC_OUT_reg_18_inst : DFFR_X1 port map( D => NPC_IN(18), CK => CLK, RN => 
                           n16, Q => NPC_OUT(18), QN => n_1533);
   NPC_OUT_reg_17_inst : DFFR_X1 port map( D => NPC_IN(17), CK => CLK, RN => 
                           n16, Q => NPC_OUT(17), QN => n_1534);
   NPC_OUT_reg_16_inst : DFFR_X1 port map( D => NPC_IN(16), CK => CLK, RN => 
                           n16, Q => NPC_OUT(16), QN => n_1535);
   NPC_OUT_reg_15_inst : DFFR_X1 port map( D => NPC_IN(15), CK => CLK, RN => 
                           n16, Q => NPC_OUT(15), QN => n_1536);
   NPC_OUT_reg_14_inst : DFFR_X1 port map( D => NPC_IN(14), CK => CLK, RN => 
                           n16, Q => NPC_OUT(14), QN => n_1537);
   NPC_OUT_reg_13_inst : DFFR_X1 port map( D => NPC_IN(13), CK => CLK, RN => 
                           n16, Q => NPC_OUT(13), QN => n_1538);
   NPC_OUT_reg_12_inst : DFFR_X1 port map( D => NPC_IN(12), CK => CLK, RN => 
                           n16, Q => NPC_OUT(12), QN => n_1539);
   NPC_OUT_reg_11_inst : DFFR_X1 port map( D => NPC_IN(11), CK => CLK, RN => 
                           n16, Q => NPC_OUT(11), QN => n_1540);
   NPC_OUT_reg_10_inst : DFFR_X1 port map( D => NPC_IN(10), CK => CLK, RN => 
                           n16, Q => NPC_OUT(10), QN => n_1541);
   NPC_OUT_reg_9_inst : DFFR_X1 port map( D => NPC_IN(9), CK => CLK, RN => n16,
                           Q => NPC_OUT(9), QN => n_1542);
   NPC_OUT_reg_8_inst : DFFR_X1 port map( D => NPC_IN(8), CK => CLK, RN => n17,
                           Q => NPC_OUT(8), QN => n_1543);
   NPC_OUT_reg_7_inst : DFFR_X1 port map( D => NPC_IN(7), CK => CLK, RN => n17,
                           Q => NPC_OUT(7), QN => n_1544);
   NPC_OUT_reg_6_inst : DFFR_X1 port map( D => NPC_IN(6), CK => CLK, RN => n17,
                           Q => NPC_OUT(6), QN => n_1545);
   NPC_OUT_reg_5_inst : DFFR_X1 port map( D => NPC_IN(5), CK => CLK, RN => n17,
                           Q => NPC_OUT(5), QN => n_1546);
   NPC_OUT_reg_4_inst : DFFR_X1 port map( D => NPC_IN(4), CK => CLK, RN => n17,
                           Q => NPC_OUT(4), QN => n_1547);
   NPC_OUT_reg_3_inst : DFFR_X1 port map( D => NPC_IN(3), CK => CLK, RN => n17,
                           Q => NPC_OUT(3), QN => n_1548);
   NPC_OUT_reg_2_inst : DFFR_X1 port map( D => NPC_IN(2), CK => CLK, RN => n17,
                           Q => NPC_OUT(2), QN => n_1549);
   NPC_OUT_reg_1_inst : DFFR_X1 port map( D => NPC_IN(1), CK => CLK, RN => n17,
                           Q => NPC_OUT(1), QN => n_1550);
   NPC_OUT_reg_0_inst : DFFR_X1 port map( D => NPC_IN(0), CK => CLK, RN => n17,
                           Q => NPC_OUT(0), QN => n_1551);
   NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => NPC_L_IN(31), CK => CLK, RN 
                           => n17, Q => NPC_L_OUT(31), QN => n_1552);
   NPC_L_OUT_reg_30_inst : DFFR_X1 port map( D => NPC_L_IN(30), CK => CLK, RN 
                           => n17, Q => NPC_L_OUT(30), QN => n_1553);
   NPC_L_OUT_reg_29_inst : DFFR_X1 port map( D => NPC_L_IN(29), CK => CLK, RN 
                           => n17, Q => NPC_L_OUT(29), QN => n_1554);
   NPC_L_OUT_reg_28_inst : DFFR_X1 port map( D => NPC_L_IN(28), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(28), QN => n_1555);
   NPC_L_OUT_reg_27_inst : DFFR_X1 port map( D => NPC_L_IN(27), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(27), QN => n_1556);
   NPC_L_OUT_reg_26_inst : DFFR_X1 port map( D => NPC_L_IN(26), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(26), QN => n_1557);
   NPC_L_OUT_reg_25_inst : DFFR_X1 port map( D => NPC_L_IN(25), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(25), QN => n_1558);
   NPC_L_OUT_reg_24_inst : DFFR_X1 port map( D => NPC_L_IN(24), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(24), QN => n_1559);
   NPC_L_OUT_reg_23_inst : DFFR_X1 port map( D => NPC_L_IN(23), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(23), QN => n_1560);
   NPC_L_OUT_reg_22_inst : DFFR_X1 port map( D => NPC_L_IN(22), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(22), QN => n_1561);
   NPC_L_OUT_reg_21_inst : DFFR_X1 port map( D => NPC_L_IN(21), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(21), QN => n_1562);
   NPC_L_OUT_reg_20_inst : DFFR_X1 port map( D => NPC_L_IN(20), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(20), QN => n_1563);
   NPC_L_OUT_reg_19_inst : DFFR_X1 port map( D => NPC_L_IN(19), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(19), QN => n_1564);
   NPC_L_OUT_reg_18_inst : DFFR_X1 port map( D => NPC_L_IN(18), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(18), QN => n_1565);
   NPC_L_OUT_reg_17_inst : DFFR_X1 port map( D => NPC_L_IN(17), CK => CLK, RN 
                           => n18, Q => NPC_L_OUT(17), QN => n_1566);
   NPC_L_OUT_reg_16_inst : DFFR_X1 port map( D => NPC_L_IN(16), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(16), QN => n_1567);
   NPC_L_OUT_reg_15_inst : DFFR_X1 port map( D => NPC_L_IN(15), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(15), QN => n_1568);
   NPC_L_OUT_reg_14_inst : DFFR_X1 port map( D => NPC_L_IN(14), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(14), QN => n_1569);
   NPC_L_OUT_reg_13_inst : DFFR_X1 port map( D => NPC_L_IN(13), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(13), QN => n_1570);
   NPC_L_OUT_reg_12_inst : DFFR_X1 port map( D => NPC_L_IN(12), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(12), QN => n_1571);
   NPC_L_OUT_reg_11_inst : DFFR_X1 port map( D => NPC_L_IN(11), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(11), QN => n_1572);
   NPC_L_OUT_reg_10_inst : DFFR_X1 port map( D => NPC_L_IN(10), CK => CLK, RN 
                           => n19, Q => NPC_L_OUT(10), QN => n_1573);
   NPC_L_OUT_reg_9_inst : DFFR_X1 port map( D => NPC_L_IN(9), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(9), QN => n_1574);
   NPC_L_OUT_reg_8_inst : DFFR_X1 port map( D => NPC_L_IN(8), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(8), QN => n_1575);
   NPC_L_OUT_reg_7_inst : DFFR_X1 port map( D => NPC_L_IN(7), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(7), QN => n_1576);
   NPC_L_OUT_reg_6_inst : DFFR_X1 port map( D => NPC_L_IN(6), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(6), QN => n_1577);
   NPC_L_OUT_reg_5_inst : DFFR_X1 port map( D => NPC_L_IN(5), CK => CLK, RN => 
                           n19, Q => NPC_L_OUT(5), QN => n_1578);
   NPC_L_OUT_reg_4_inst : DFFR_X1 port map( D => NPC_L_IN(4), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(4), QN => n_1579);
   NPC_L_OUT_reg_3_inst : DFFR_X1 port map( D => NPC_L_IN(3), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(3), QN => n_1580);
   NPC_L_OUT_reg_2_inst : DFFR_X1 port map( D => NPC_L_IN(2), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(2), QN => n_1581);
   NPC_L_OUT_reg_1_inst : DFFR_X1 port map( D => NPC_L_IN(1), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(1), QN => n_1582);
   NPC_L_OUT_reg_0_inst : DFFR_X1 port map( D => NPC_L_IN(0), CK => CLK, RN => 
                           n20, Q => NPC_L_OUT(0), QN => n_1583);
   RS1_OUT_reg_4_inst : DFFR_X1 port map( D => RS1_IN(4), CK => CLK, RN => n20,
                           Q => RS1_OUT(4), QN => n_1584);
   RS1_OUT_reg_3_inst : DFFR_X1 port map( D => RS1_IN(3), CK => CLK, RN => n20,
                           Q => RS1_OUT(3), QN => n_1585);
   RS1_OUT_reg_2_inst : DFFR_X1 port map( D => RS1_IN(2), CK => CLK, RN => n20,
                           Q => RS1_OUT(2), QN => n_1586);
   RS1_OUT_reg_1_inst : DFFR_X1 port map( D => RS1_IN(1), CK => CLK, RN => n20,
                           Q => RS1_OUT(1), QN => n_1587);
   RS1_OUT_reg_0_inst : DFFR_X1 port map( D => RS1_IN(0), CK => CLK, RN => n20,
                           Q => RS1_OUT(0), QN => n_1588);
   RS2_OUT_reg_4_inst : DFFR_X1 port map( D => RS2_IN(4), CK => CLK, RN => n20,
                           Q => RS2_OUT(4), QN => n_1589);
   RS2_OUT_reg_3_inst : DFFR_X1 port map( D => RS2_IN(3), CK => CLK, RN => n20,
                           Q => RS2_OUT(3), QN => n_1590);
   RS2_OUT_reg_2_inst : DFFR_X1 port map( D => RS2_IN(2), CK => CLK, RN => n21,
                           Q => RS2_OUT(2), QN => n_1591);
   RS2_OUT_reg_1_inst : DFFR_X1 port map( D => RS2_IN(1), CK => CLK, RN => n21,
                           Q => RS2_OUT(1), QN => n_1592);
   RS2_OUT_reg_0_inst : DFFR_X1 port map( D => RS2_IN(0), CK => CLK, RN => n21,
                           Q => RS2_OUT(0), QN => n_1593);
   RD_OUT_reg_4_inst : DFFR_X1 port map( D => RD_IN(4), CK => CLK, RN => n21, Q
                           => RD_OUT(4), QN => n_1594);
   RD_OUT_reg_3_inst : DFFR_X1 port map( D => RD_IN(3), CK => CLK, RN => n21, Q
                           => RD_OUT(3), QN => n_1595);
   RD_OUT_reg_2_inst : DFFR_X1 port map( D => RD_IN(2), CK => CLK, RN => n21, Q
                           => RD_OUT(2), QN => n_1596);
   RD_OUT_reg_1_inst : DFFR_X1 port map( D => RD_IN(1), CK => CLK, RN => n21, Q
                           => RD_OUT(1), QN => n_1597);
   RD_OUT_reg_0_inst : DFFR_X1 port map( D => RD_IN(0), CK => CLK, RN => n21, Q
                           => RD_OUT(0), QN => n_1598);
   OPCODE_OUT_reg_5_inst : DFFR_X1 port map( D => OPCODE_IN(5), CK => CLK, RN 
                           => n21, Q => OPCODE_OUT(5), QN => n_1599);
   OPCODE_OUT_reg_4_inst : DFFR_X1 port map( D => OPCODE_IN(4), CK => CLK, RN 
                           => n21, Q => OPCODE_OUT(4), QN => n_1600);
   OPCODE_OUT_reg_3_inst : DFFR_X1 port map( D => OPCODE_IN(3), CK => CLK, RN 
                           => n21, Q => OPCODE_OUT(3), QN => n_1601);
   OPCODE_OUT_reg_2_inst : DFFR_X1 port map( D => OPCODE_IN(2), CK => CLK, RN 
                           => n21, Q => n_1602, QN => n2);
   OPCODE_OUT_reg_1_inst : DFFR_X1 port map( D => OPCODE_IN(1), CK => CLK, RN 
                           => n22, Q => OPCODE_OUT(1), QN => n_1603);
   OPCODE_OUT_reg_0_inst : DFFR_X1 port map( D => OPCODE_IN(0), CK => CLK, RN 
                           => n22, Q => OPCODE_OUT(0), QN => n_1604);
   IR_OUT_reg_15_inst : DFFR_X1 port map( D => IR_IN(15), CK => CLK, RN => n22,
                           Q => IR_OUT(15), QN => n_1605);
   IR_OUT_reg_14_inst : DFFR_X1 port map( D => IR_IN(14), CK => CLK, RN => n22,
                           Q => IR_OUT(14), QN => n_1606);
   IR_OUT_reg_13_inst : DFFR_X1 port map( D => IR_IN(13), CK => CLK, RN => n22,
                           Q => IR_OUT(13), QN => n_1607);
   IR_OUT_reg_12_inst : DFFR_X1 port map( D => IR_IN(12), CK => CLK, RN => n22,
                           Q => IR_OUT(12), QN => n_1608);
   IR_OUT_reg_11_inst : DFFR_X1 port map( D => IR_IN(11), CK => CLK, RN => n22,
                           Q => IR_OUT(11), QN => n_1609);
   IR_OUT_reg_10_inst : DFFR_X1 port map( D => IR_IN(10), CK => CLK, RN => n22,
                           Q => IR_OUT(10), QN => n_1610);
   IR_OUT_reg_9_inst : DFFR_X1 port map( D => IR_IN(9), CK => CLK, RN => n22, Q
                           => IR_OUT(9), QN => n_1611);
   IR_OUT_reg_8_inst : DFFR_X1 port map( D => IR_IN(8), CK => CLK, RN => n22, Q
                           => IR_OUT(8), QN => n_1612);
   IR_OUT_reg_7_inst : DFFR_X1 port map( D => IR_IN(7), CK => CLK, RN => n22, Q
                           => IR_OUT(7), QN => n_1613);
   IR_OUT_reg_6_inst : DFFR_X1 port map( D => IR_IN(6), CK => CLK, RN => n22, Q
                           => IR_OUT(6), QN => n_1614);
   IR_OUT_reg_5_inst : DFFR_X1 port map( D => IR_IN(5), CK => CLK, RN => n23, Q
                           => IR_OUT(5), QN => n_1615);
   IR_OUT_reg_4_inst : DFFR_X1 port map( D => IR_IN(4), CK => CLK, RN => n23, Q
                           => IR_OUT(4), QN => n_1616);
   IR_OUT_reg_3_inst : DFFR_X1 port map( D => IR_IN(3), CK => CLK, RN => n23, Q
                           => IR_OUT(3), QN => n_1617);
   IR_OUT_reg_2_inst : DFFR_X1 port map( D => IR_IN(2), CK => CLK, RN => n23, Q
                           => IR_OUT(2), QN => n_1618);
   IR_OUT_reg_1_inst : DFFR_X1 port map( D => IR_IN(1), CK => CLK, RN => n23, Q
                           => IR_OUT(1), QN => n_1619);
   IR_OUT_reg_0_inst : DFFR_X1 port map( D => IR_IN(0), CK => CLK, RN => n23, Q
                           => IR_OUT(0), QN => n_1620);
   U3 : INV_X1 port map( A => n2, ZN => OPCODE_OUT(2));
   U4 : BUF_X1 port map( A => RST, Z => n5);
   U5 : BUF_X1 port map( A => RST, Z => n4);
   U6 : BUF_X1 port map( A => RST, Z => n6);
   U7 : CLKBUF_X1 port map( A => n4, Z => n7);
   U8 : CLKBUF_X1 port map( A => n4, Z => n8);
   U9 : CLKBUF_X1 port map( A => n4, Z => n9);
   U10 : CLKBUF_X1 port map( A => n4, Z => n10);
   U11 : CLKBUF_X1 port map( A => n4, Z => n11);
   U12 : CLKBUF_X1 port map( A => n4, Z => n12);
   U13 : CLKBUF_X1 port map( A => n5, Z => n13);
   U14 : CLKBUF_X1 port map( A => n5, Z => n14);
   U15 : CLKBUF_X1 port map( A => n5, Z => n15);
   U16 : CLKBUF_X1 port map( A => n5, Z => n16);
   U17 : CLKBUF_X1 port map( A => n5, Z => n17);
   U18 : CLKBUF_X1 port map( A => n5, Z => n18);
   U19 : CLKBUF_X1 port map( A => n6, Z => n19);
   U20 : CLKBUF_X1 port map( A => n6, Z => n20);
   U21 : CLKBUF_X1 port map( A => n6, Z => n21);
   U22 : CLKBUF_X1 port map( A => n6, Z => n22);
   U23 : CLKBUF_X1 port map( A => n6, Z => n23);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity sign_extender is

   port( d_in : in std_logic_vector (31 downto 0);  rst : in std_logic;  d_ext 
         : out std_logic_vector (31 downto 0));

end sign_extender;

architecture SYN_Behavioral of sign_extender is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal d_ext_31_port, d_ext_24_port, d_ext_23_port, d_ext_22_port, 
      d_ext_21_port, d_ext_20_port, d_ext_19_port, d_ext_18_port, d_ext_17_port
      , d_ext_16_port, d_ext_15_port, d_ext_14_port, d_ext_13_port, 
      d_ext_12_port, d_ext_11_port, d_ext_10_port, d_ext_9_port, d_ext_8_port, 
      d_ext_7_port, d_ext_6_port, d_ext_5_port, d_ext_4_port, d_ext_3_port, 
      d_ext_2_port, d_ext_1_port, d_ext_0_port, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n1, n2, n3, n4, n5, n6, n7, n30 : std_logic;

begin
   d_ext <= ( d_ext_31_port, d_ext_31_port, d_ext_31_port, d_ext_31_port, 
      d_ext_31_port, d_ext_31_port, d_ext_31_port, d_ext_24_port, d_ext_23_port
      , d_ext_22_port, d_ext_21_port, d_ext_20_port, d_ext_19_port, 
      d_ext_18_port, d_ext_17_port, d_ext_16_port, d_ext_15_port, d_ext_14_port
      , d_ext_13_port, d_ext_12_port, d_ext_11_port, d_ext_10_port, 
      d_ext_9_port, d_ext_8_port, d_ext_7_port, d_ext_6_port, d_ext_5_port, 
      d_ext_4_port, d_ext_3_port, d_ext_2_port, d_ext_1_port, d_ext_0_port );
   
   U56 : OAI33_X1 port map( A1 => n5, A2 => d_in(28), A3 => d_in(27), B1 => n7,
                           B2 => n27, B3 => n30, ZN => n26);
   U2 : NAND3_X1 port map( A1 => n1, A2 => n10, A3 => n9, ZN => n11);
   U3 : NOR2_X1 port map( A1 => n10, A2 => n2, ZN => n13);
   U4 : INV_X1 port map( A => rst, ZN => n2);
   U5 : AOI21_X1 port map( B1 => d_in(29), B2 => d_in(26), A => d_in(31), ZN =>
                           n27);
   U6 : OAI22_X1 port map( A1 => n6, A2 => n5, B1 => d_in(28), B2 => d_in(26), 
                           ZN => n25);
   U7 : INV_X1 port map( A => d_in(28), ZN => n7);
   U8 : NOR2_X1 port map( A1 => n8, A2 => n2, ZN => d_ext_31_port);
   U9 : AOI22_X1 port map( A1 => n9, A2 => n10, B1 => d_in(25), B2 => n4, ZN =>
                           n8);
   U10 : INV_X1 port map( A => n10, ZN => n4);
   U11 : AOI21_X1 port map( B1 => n30, B2 => d_in(26), A => d_in(31), ZN => n28
                           );
   U12 : INV_X1 port map( A => d_in(30), ZN => n5);
   U13 : INV_X1 port map( A => d_in(27), ZN => n30);
   U14 : AND2_X1 port map( A1 => d_in(15), A2 => n22, ZN => n9);
   U15 : OAI221_X1 port map( B1 => d_in(29), B2 => n23, C1 => d_in(30), C2 => 
                           n3, A => n24, ZN => n22);
   U16 : AND3_X1 port map( A1 => n28, A2 => d_in(28), A3 => d_in(30), ZN => n23
                           );
   U17 : AOI21_X1 port map( B1 => n25, B2 => n3, A => n26, ZN => n24);
   U18 : NAND2_X1 port map( A1 => n11, A2 => n21, ZN => d_ext_16_port);
   U19 : NAND2_X1 port map( A1 => d_in(16), A2 => n13, ZN => n21);
   U20 : NAND2_X1 port map( A1 => n11, A2 => n20, ZN => d_ext_17_port);
   U21 : NAND2_X1 port map( A1 => d_in(17), A2 => n13, ZN => n20);
   U22 : NAND2_X1 port map( A1 => n11, A2 => n19, ZN => d_ext_18_port);
   U23 : NAND2_X1 port map( A1 => d_in(18), A2 => n13, ZN => n19);
   U24 : NAND2_X1 port map( A1 => n11, A2 => n18, ZN => d_ext_19_port);
   U25 : NAND2_X1 port map( A1 => d_in(19), A2 => n13, ZN => n18);
   U26 : NAND2_X1 port map( A1 => n11, A2 => n17, ZN => d_ext_20_port);
   U27 : NAND2_X1 port map( A1 => d_in(20), A2 => n13, ZN => n17);
   U28 : NAND2_X1 port map( A1 => n11, A2 => n16, ZN => d_ext_21_port);
   U29 : NAND2_X1 port map( A1 => d_in(21), A2 => n13, ZN => n16);
   U30 : NAND2_X1 port map( A1 => n11, A2 => n15, ZN => d_ext_22_port);
   U31 : NAND2_X1 port map( A1 => d_in(22), A2 => n13, ZN => n15);
   U32 : NAND2_X1 port map( A1 => n11, A2 => n14, ZN => d_ext_23_port);
   U33 : NAND2_X1 port map( A1 => d_in(23), A2 => n13, ZN => n14);
   U34 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => d_ext_24_port);
   U35 : NAND2_X1 port map( A1 => d_in(24), A2 => n13, ZN => n12);
   U36 : NAND4_X1 port map( A1 => d_in(27), A2 => n7, A3 => n29, A4 => n6, ZN 
                           => n10);
   U37 : NOR2_X1 port map( A1 => d_in(31), A2 => d_in(30), ZN => n29);
   U38 : INV_X1 port map( A => d_in(29), ZN => n6);
   U39 : INV_X1 port map( A => d_in(31), ZN => n3);
   U40 : AND2_X1 port map( A1 => d_in(5), A2 => n1, ZN => d_ext_5_port);
   U41 : AND2_X1 port map( A1 => d_in(0), A2 => n1, ZN => d_ext_0_port);
   U42 : AND2_X1 port map( A1 => d_in(1), A2 => n1, ZN => d_ext_1_port);
   U43 : AND2_X1 port map( A1 => d_in(2), A2 => n1, ZN => d_ext_2_port);
   U44 : AND2_X1 port map( A1 => d_in(3), A2 => n1, ZN => d_ext_3_port);
   U45 : AND2_X1 port map( A1 => d_in(4), A2 => n1, ZN => d_ext_4_port);
   U46 : AND2_X1 port map( A1 => d_in(6), A2 => n1, ZN => d_ext_6_port);
   U47 : AND2_X1 port map( A1 => d_in(7), A2 => n1, ZN => d_ext_7_port);
   U48 : AND2_X1 port map( A1 => d_in(8), A2 => n1, ZN => d_ext_8_port);
   U49 : AND2_X1 port map( A1 => d_in(10), A2 => n1, ZN => d_ext_10_port);
   U50 : AND2_X1 port map( A1 => d_in(13), A2 => n1, ZN => d_ext_13_port);
   U51 : AND2_X1 port map( A1 => d_in(14), A2 => n1, ZN => d_ext_14_port);
   U52 : AND2_X1 port map( A1 => n1, A2 => d_in(9), ZN => d_ext_9_port);
   U53 : AND2_X1 port map( A1 => n1, A2 => d_in(15), ZN => d_ext_15_port);
   U54 : AND2_X1 port map( A1 => d_in(11), A2 => n1, ZN => d_ext_11_port);
   U55 : AND2_X1 port map( A1 => d_in(12), A2 => n1, ZN => d_ext_12_port);
   U57 : INV_X1 port map( A => n2, ZN => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity register_file_N32_addBit5 is

   port( RESET, RE, WE : in std_logic;  ADD_WR, ADD_RDA, ADD_RDB : in 
         std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUTA, OUTB : out std_logic_vector (31 downto 0));

end register_file_N32_addBit5;

architecture SYN_A of register_file_N32_addBit5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N243, N244, N245, N246, N247, 
      N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, 
      N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N307, N308, 
      N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, 
      N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, 
      N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, 
      N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, 
      N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, 
      N369, N370, N371, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, 
      n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
      n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
      n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
      n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, 
      n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, 
      n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
      n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
      n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, 
      n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
      n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
      n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, 
      n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
      n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
      n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, 
      n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, 
      n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
      n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
      n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
      n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, 
      n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
      n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
      n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, 
      n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, 
      n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
      n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, 
      n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
      n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, 
      n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
      n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, 
      n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, 
      n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
      n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, 
      n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
      n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
      n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
      n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
      n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
      n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, 
      n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
      n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
      n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
      n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
      n1785, n1786, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243_port, 
      n244_port, n245_port, n246_port, n247_port, n248_port, n249_port, 
      n250_port, n251_port, n252_port, n253_port, n254_port, n255_port, 
      n256_port, n257_port, n258_port, n259_port, n260_port, n261_port, 
      n262_port, n263_port, n264_port, n265_port, n266_port, n267_port, 
      n268_port, n269_port, n270_port, n271_port, n272_port, n273_port, 
      n274_port, n275_port, n276_port, n277_port, n278_port, n279_port, 
      n280_port, n281_port, n282_port, n283_port, n284_port, n285_port, 
      n286_port, n287_port, n288_port, n289_port, n290_port, n291_port, 
      n292_port, n293_port, n294_port, n295_port, n296_port, n297_port, 
      n298_port, n299_port, n300_port, n301_port, n302_port, n303_port, 
      n304_port, n305_port, n306, n307_port, n308_port, n309_port, n310_port, 
      n311_port, n312_port, n313_port, n314_port, n315_port, n316_port, 
      n317_port, n318_port, n319_port, n320_port, n321_port, n322_port, 
      n323_port, n324_port, n325_port, n326_port, n327_port, n328_port, 
      n329_port, n330_port, n331_port, n332_port, n333_port, n334_port, 
      n335_port, n336_port, n337_port, n338_port, n339_port, n340_port, 
      n341_port, n342_port, n343_port, n344_port, n345_port, n346_port, 
      n347_port, n348_port, n349_port, n350_port, n351_port, n352_port, 
      n353_port, n354_port, n355_port, n356_port, n357_port, n358_port, 
      n359_port, n360_port, n361_port, n362_port, n363_port, n364_port, 
      n365_port, n366_port, n367_port, n368_port, n369_port, n370_port, 
      n371_port, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n558, n1182, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794
      , n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, 
      n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, 
      n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, 
      n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
      n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
      n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
      n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
      n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
      n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
      n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
      n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
      n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, 
      n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, 
      n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, 
      n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
      n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, 
      n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
      n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
      n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157 : std_logic;

begin
   
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => n195, D => n283_port, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => n195, D => n286_port, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => n195, D => n289_port, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => n195, D => n292_port, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => n195, D => n295_port, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => n195, D => n298_port, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => n195, D => n301_port, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => n195, D => n304_port, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => n195, D => n307_port, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => n195, D => n310_port, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => n194, D => n313_port, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => n194, D => n316_port, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => n194, D => n319_port, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => n194, D => n322_port, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => n194, D => n325_port, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => n194, D => n328_port, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => n194, D => n331_port, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => n194, D => n334_port, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => n194, D => n337_port, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => n194, D => n340_port, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => n194, D => n343_port, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => n193, D => n346_port, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => n193, D => n349_port, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => n193, D => n352_port, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => n193, D => n355_port, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => n193, D => n358_port, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => n193, D => n361_port, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => n193, D => n364_port, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => n193, D => n367_port, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => n193, D => n370_port, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => n193, D => n373, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => n193, D => n376, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => n198, D => n283_port, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => n198, D => n286_port, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => n198, D => n289_port, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => n198, D => n292_port, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => n198, D => n295_port, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => n198, D => n298_port, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => n198, D => n301_port, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => n198, D => n304_port, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => n198, D => n307_port, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => n198, D => n310_port, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => n197, D => n313_port, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => n197, D => n316_port, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => n197, D => n319_port, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => n197, D => n322_port, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => n197, D => n325_port, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => n197, D => n328_port, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => n197, D => n331_port, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => n197, D => n334_port, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => n197, D => n337_port, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => n197, D => n340_port, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => n197, D => n343_port, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => n196, D => n346_port, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => n196, D => n349_port, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => n196, D => n352_port, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => n196, D => n355_port, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => n196, D => n358_port, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => n196, D => n361_port, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => n196, D => n364_port, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => n196, D => n367_port, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => n196, D => n370_port, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => n196, D => n373, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => n196, D => n376, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => n201, D => n283_port, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => n201, D => n286_port, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => n201, D => n289_port, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => n201, D => n292_port, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => n201, D => n295_port, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => n201, D => n298_port, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => n201, D => n301_port, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => n201, D => n304_port, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => n201, D => n307_port, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => n201, D => n310_port, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => n200, D => n313_port, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => n200, D => n316_port, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => n200, D => n319_port, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => n200, D => n322_port, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => n200, D => n325_port, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => n200, D => n328_port, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => n200, D => n331_port, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => n200, D => n334_port, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => n200, D => n337_port, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => n200, D => n340_port, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => n200, D => n343_port, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => n199, D => n346_port, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => n199, D => n349_port, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => n199, D => n352_port, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => n199, D => n355_port, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => n199, D => n358_port, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => n199, D => n361_port, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => n199, D => n364_port, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => n199, D => n367_port, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => n199, D => n370_port, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => n199, D => n373, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => n199, D => n376, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => n204, D => n283_port, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => n204, D => n286_port, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => n204, D => n289_port, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => n204, D => n292_port, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => n204, D => n295_port, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => n204, D => n298_port, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => n204, D => n301_port, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => n204, D => n304_port, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => n204, D => n307_port, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => n204, D => n310_port, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => n203, D => n313_port, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => n203, D => n316_port, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => n203, D => n319_port, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => n203, D => n322_port, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => n203, D => n325_port, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => n203, D => n328_port, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => n203, D => n331_port, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => n203, D => n334_port, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => n203, D => n337_port, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => n203, D => n340_port, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => n203, D => n343_port, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => n202, D => n346_port, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => n202, D => n349_port, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => n202, D => n352_port, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => n202, D => n355_port, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => n202, D => n358_port, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => n202, D => n361_port, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => n202, D => n364_port, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => n202, D => n367_port, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => n202, D => n370_port, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => n202, D => n373, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => n202, D => n376, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => n207, D => n283_port, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => n207, D => n286_port, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => n207, D => n289_port, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => n207, D => n292_port, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => n207, D => n295_port, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => n207, D => n298_port, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => n207, D => n301_port, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => n207, D => n304_port, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => n207, D => n307_port, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => n207, D => n310_port, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => n206, D => n313_port, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => n206, D => n316_port, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => n206, D => n319_port, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => n206, D => n322_port, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => n206, D => n325_port, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => n206, D => n328_port, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => n206, D => n331_port, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => n206, D => n334_port, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => n206, D => n337_port, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => n206, D => n340_port, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => n206, D => n343_port, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => n205, D => n346_port, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => n205, D => n349_port, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => n205, D => n352_port, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => n205, D => n355_port, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => n205, D => n358_port, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => n205, D => n361_port, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => n205, D => n364_port, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => n205, D => n367_port, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => n205, D => n370_port, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => n205, D => n373, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => n205, D => n376, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => n210, D => n283_port, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => n210, D => n286_port, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => n210, D => n289_port, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => n210, D => n292_port, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => n210, D => n295_port, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => n210, D => n298_port, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => n210, D => n301_port, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => n210, D => n304_port, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => n210, D => n307_port, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => n210, D => n310_port, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => n209, D => n313_port, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => n209, D => n316_port, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => n209, D => n319_port, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => n209, D => n322_port, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => n209, D => n325_port, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => n209, D => n328_port, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => n209, D => n331_port, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => n209, D => n334_port, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => n209, D => n337_port, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => n209, D => n340_port, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => n209, D => n343_port, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => n208, D => n346_port, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => n208, D => n349_port, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => n208, D => n352_port, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => n208, D => n355_port, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => n208, D => n358_port, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => n208, D => n361_port, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => n208, D => n364_port, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => n208, D => n367_port, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => n208, D => n370_port, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => n208, D => n373, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => n208, D => n376, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => n213, D => n283_port, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => n213, D => n286_port, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => n213, D => n289_port, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => n213, D => n292_port, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => n213, D => n295_port, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => n213, D => n298_port, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => n213, D => n301_port, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => n213, D => n304_port, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => n213, D => n307_port, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => n213, D => n310_port, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => n212, D => n313_port, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => n212, D => n316_port, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => n212, D => n319_port, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => n212, D => n322_port, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => n212, D => n325_port, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => n212, D => n328_port, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => n212, D => n331_port, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => n212, D => n334_port, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => n212, D => n337_port, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => n212, D => n340_port, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => n212, D => n343_port, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => n211, D => n346_port, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => n211, D => n349_port, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => n211, D => n352_port, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => n211, D => n355_port, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => n211, D => n358_port, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => n211, D => n361_port, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => n211, D => n364_port, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => n211, D => n367_port, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => n211, D => n370_port, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => n211, D => n373, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => n211, D => n376, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => n216, D => n283_port, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => n216, D => n286_port, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => n216, D => n289_port, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => n216, D => n292_port, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => n216, D => n295_port, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => n216, D => n298_port, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => n216, D => n301_port, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => n216, D => n304_port, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => n216, D => n307_port, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => n216, D => n310_port, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => n215, D => n313_port, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => n215, D => n316_port, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => n215, D => n319_port, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => n215, D => n322_port, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => n215, D => n325_port, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => n215, D => n328_port, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => n215, D => n331_port, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => n215, D => n334_port, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => n215, D => n337_port, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => n215, D => n340_port, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => n215, D => n343_port, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => n214, D => n346_port, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => n214, D => n349_port, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => n214, D => n352_port, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => n214, D => n355_port, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => n214, D => n358_port, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => n214, D => n361_port, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => n214, D => n364_port, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => n214, D => n367_port, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => n214, D => n370_port, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => n214, D => n373, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => n214, D => n376, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => n219, D => n283_port, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => n219, D => n286_port, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => n219, D => n289_port, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => n219, D => n292_port, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => n219, D => n295_port, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => n219, D => n298_port, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => n219, D => n301_port, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => n219, D => n304_port, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => n219, D => n307_port, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => n219, D => n310_port, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => n218, D => n313_port, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => n218, D => n316_port, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => n218, D => n319_port, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => n218, D => n322_port, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => n218, D => n325_port, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => n218, D => n328_port, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => n218, D => n331_port, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => n218, D => n334_port, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => n218, D => n337_port, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => n218, D => n340_port, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => n218, D => n343_port, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => n217, D => n346_port, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => n217, D => n349_port, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => n217, D => n352_port, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => n217, D => n355_port, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => n217, D => n358_port, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => n217, D => n361_port, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => n217, D => n364_port, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => n217, D => n367_port, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => n217, D => n370_port, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => n217, D => n373, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => n217, D => n376, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => n222, D => n283_port, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => n222, D => n286_port, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => n222, D => n289_port, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => n222, D => n292_port, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => n222, D => n295_port, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => n222, D => n298_port, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => n222, D => n301_port, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => n222, D => n304_port, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => n222, D => n307_port, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => n222, D => n310_port, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => n221, D => n313_port, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => n221, D => n316_port, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => n221, D => n319_port, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => n221, D => n322_port, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => n221, D => n325_port, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => n221, D => n328_port, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => n221, D => n331_port, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => n221, D => n334_port, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => n221, D => n337_port, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => n221, D => n340_port, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => n221, D => n343_port, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => n220, D => n346_port, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => n220, D => n349_port, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => n220, D => n352_port, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => n220, D => n355_port, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => n220, D => n358_port, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => n220, D => n361_port, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => n220, D => n364_port, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => n220, D => n367_port, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => n220, D => n370_port, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => n220, D => n373, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => n220, D => n376, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => n225, D => n283_port, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => n225, D => n286_port, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => n225, D => n289_port, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => n225, D => n292_port, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => n225, D => n295_port, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => n225, D => n298_port, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => n225, D => n301_port, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => n225, D => n304_port, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => n225, D => n307_port, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => n225, D => n310_port, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => n224, D => n313_port, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => n224, D => n316_port, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => n224, D => n319_port, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => n224, D => n322_port, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => n224, D => n325_port, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => n224, D => n328_port, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => n224, D => n331_port, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => n224, D => n334_port, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => n224, D => n337_port, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => n224, D => n340_port, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => n224, D => n343_port, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => n223, D => n346_port, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => n223, D => n349_port, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => n223, D => n352_port, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => n223, D => n355_port, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => n223, D => n358_port, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => n223, D => n361_port, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => n223, D => n364_port, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => n223, D => n367_port, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => n223, D => n370_port, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => n223, D => n373, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => n223, D => n376, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => n228, D => n284_port, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => n228, D => n287_port, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => n228, D => n290_port, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => n228, D => n293_port, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => n228, D => n296_port, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => n228, D => n299_port, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => n228, D => n302_port, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => n228, D => n305_port, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => n228, D => n308_port, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => n228, D => n311_port, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => n227, D => n314_port, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => n227, D => n317_port, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => n227, D => n320_port, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => n227, D => n323_port, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => n227, D => n326_port, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => n227, D => n329_port, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => n227, D => n332_port, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => n227, D => n335_port, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => n227, D => n338_port, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => n227, D => n341_port, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => n227, D => n344_port, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => n226, D => n347_port, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => n226, D => n350_port, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => n226, D => n353_port, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => n226, D => n356_port, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => n226, D => n359_port, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => n226, D => n362_port, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => n226, D => n365_port, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => n226, D => n368_port, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => n226, D => n371_port, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => n226, D => n374, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => n226, D => n377, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => n231, D => n284_port, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => n231, D => n287_port, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => n231, D => n290_port, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => n231, D => n293_port, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => n231, D => n296_port, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => n231, D => n299_port, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => n231, D => n302_port, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => n231, D => n305_port, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => n231, D => n308_port, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => n231, D => n311_port, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => n230, D => n314_port, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => n230, D => n317_port, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => n230, D => n320_port, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => n230, D => n323_port, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => n230, D => n326_port, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => n230, D => n329_port, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => n230, D => n332_port, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => n230, D => n335_port, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => n230, D => n338_port, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => n230, D => n341_port, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => n230, D => n344_port, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => n229, D => n347_port, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => n229, D => n350_port, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => n229, D => n353_port, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => n229, D => n356_port, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => n229, D => n359_port, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => n229, D => n362_port, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => n229, D => n365_port, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => n229, D => n368_port, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => n229, D => n371_port, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => n229, D => n374, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => n229, D => n377, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => n234, D => n284_port, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => n234, D => n287_port, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => n234, D => n290_port, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => n234, D => n293_port, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => n234, D => n296_port, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => n234, D => n299_port, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => n234, D => n302_port, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => n234, D => n305_port, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => n234, D => n308_port, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => n234, D => n311_port, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => n233, D => n314_port, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => n233, D => n317_port, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => n233, D => n320_port, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => n233, D => n323_port, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => n233, D => n326_port, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => n233, D => n329_port, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => n233, D => n332_port, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => n233, D => n335_port, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => n233, D => n338_port, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => n233, D => n341_port, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => n233, D => n344_port, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => n232, D => n347_port, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => n232, D => n350_port, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => n232, D => n353_port, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => n232, D => n356_port, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => n232, D => n359_port, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => n232, D => n362_port, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => n232, D => n365_port, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => n232, D => n368_port, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => n232, D => n371_port, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => n232, D => n374, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => n232, D => n377, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => n237, D => n284_port, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => n237, D => n287_port, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => n237, D => n290_port, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => n237, D => n293_port, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => n237, D => n296_port, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => n237, D => n299_port, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => n237, D => n302_port, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => n237, D => n305_port, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => n237, D => n308_port, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => n237, D => n311_port, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => n236, D => n314_port, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => n236, D => n317_port, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => n236, D => n320_port, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => n236, D => n323_port, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => n236, D => n326_port, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => n236, D => n329_port, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => n236, D => n332_port, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => n236, D => n335_port, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => n236, D => n338_port, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => n236, D => n341_port, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => n236, D => n344_port, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => n235, D => n347_port, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => n235, D => n350_port, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => n235, D => n353_port, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => n235, D => n356_port, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => n235, D => n359_port, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => n235, D => n362_port, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => n235, D => n365_port, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => n235, D => n368_port, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => n235, D => n371_port, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => n235, D => n374, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => n235, D => n377, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => n240, D => n284_port, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => n240, D => n287_port, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => n240, D => n290_port, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => n240, D => n293_port, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => n240, D => n296_port, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => n240, D => n299_port, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => n240, D => n302_port, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => n240, D => n305_port, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => n240, D => n308_port, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => n240, D => n311_port, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => n239, D => n314_port, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => n239, D => n317_port, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => n239, D => n320_port, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => n239, D => n323_port, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => n239, D => n326_port, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => n239, D => n329_port, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => n239, D => n332_port, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => n239, D => n335_port, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => n239, D => n338_port, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => n239, D => n341_port, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => n239, D => n344_port, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => n238, D => n347_port, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => n238, D => n350_port, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => n238, D => n353_port, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => n238, D => n356_port, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => n238, D => n359_port, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => n238, D => n362_port, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => n238, D => n365_port, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => n238, D => n368_port, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => n238, D => n371_port, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => n238, D => n374, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => n238, D => n377, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => n243_port, D => n284_port, 
                           Q => REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => n243_port, D => n287_port, 
                           Q => REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => n243_port, D => n290_port, 
                           Q => REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => n243_port, D => n293_port, 
                           Q => REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => n243_port, D => n296_port, 
                           Q => REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => n243_port, D => n299_port, 
                           Q => REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => n243_port, D => n302_port, 
                           Q => REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => n243_port, D => n305_port, 
                           Q => REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => n243_port, D => n308_port, 
                           Q => REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => n243_port, D => n311_port, 
                           Q => REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => n242, D => n314_port, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => n242, D => n317_port, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => n242, D => n320_port, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => n242, D => n323_port, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => n242, D => n326_port, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => n242, D => n329_port, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => n242, D => n332_port, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => n242, D => n335_port, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => n242, D => n338_port, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => n242, D => n341_port, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => n242, D => n344_port, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => n241, D => n347_port, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => n241, D => n350_port, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => n241, D => n353_port, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => n241, D => n356_port, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => n241, D => n359_port, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => n241, D => n362_port, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => n241, D => n365_port, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => n241, D => n368_port, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => n241, D => n371_port, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => n241, D => n374, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => n241, D => n377, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => n246_port, D => n284_port, 
                           Q => REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => n246_port, D => n287_port, 
                           Q => REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => n246_port, D => n290_port, 
                           Q => REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => n246_port, D => n293_port, 
                           Q => REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => n246_port, D => n296_port, 
                           Q => REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => n246_port, D => n299_port, 
                           Q => REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => n246_port, D => n302_port, 
                           Q => REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => n246_port, D => n305_port, 
                           Q => REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => n246_port, D => n308_port, 
                           Q => REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => n246_port, D => n311_port, 
                           Q => REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => n245_port, D => n314_port, 
                           Q => REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => n245_port, D => n317_port, 
                           Q => REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => n245_port, D => n320_port, 
                           Q => REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => n245_port, D => n323_port, 
                           Q => REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => n245_port, D => n326_port, 
                           Q => REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => n245_port, D => n329_port, 
                           Q => REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => n245_port, D => n332_port, 
                           Q => REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => n245_port, D => n335_port, 
                           Q => REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => n245_port, D => n338_port, 
                           Q => REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => n245_port, D => n341_port, 
                           Q => REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => n245_port, D => n344_port, 
                           Q => REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => n244_port, D => n347_port, 
                           Q => REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => n244_port, D => n350_port, Q
                           => REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => n244_port, D => n353_port, Q
                           => REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => n244_port, D => n356_port, Q
                           => REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => n244_port, D => n359_port, Q
                           => REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => n244_port, D => n362_port, Q
                           => REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => n244_port, D => n365_port, Q
                           => REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => n244_port, D => n368_port, Q
                           => REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => n244_port, D => n371_port, Q
                           => REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => n244_port, D => n374, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => n244_port, D => n377, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => n249_port, D => n284_port, 
                           Q => REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => n249_port, D => n287_port, 
                           Q => REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => n249_port, D => n290_port, 
                           Q => REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => n249_port, D => n293_port, 
                           Q => REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => n249_port, D => n296_port, 
                           Q => REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => n249_port, D => n299_port, 
                           Q => REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => n249_port, D => n302_port, 
                           Q => REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => n249_port, D => n305_port, 
                           Q => REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => n249_port, D => n308_port, 
                           Q => REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => n249_port, D => n311_port, 
                           Q => REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => n248_port, D => n314_port, 
                           Q => REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => n248_port, D => n317_port, 
                           Q => REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => n248_port, D => n320_port, 
                           Q => REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => n248_port, D => n323_port, 
                           Q => REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => n248_port, D => n326_port, 
                           Q => REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => n248_port, D => n329_port, 
                           Q => REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => n248_port, D => n332_port, 
                           Q => REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => n248_port, D => n335_port, 
                           Q => REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => n248_port, D => n338_port, 
                           Q => REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => n248_port, D => n341_port, 
                           Q => REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => n248_port, D => n344_port, 
                           Q => REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => n247_port, D => n347_port, 
                           Q => REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => n247_port, D => n350_port, Q
                           => REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => n247_port, D => n353_port, Q
                           => REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => n247_port, D => n356_port, Q
                           => REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => n247_port, D => n359_port, Q
                           => REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => n247_port, D => n362_port, Q
                           => REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => n247_port, D => n365_port, Q
                           => REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => n247_port, D => n368_port, Q
                           => REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => n247_port, D => n371_port, Q
                           => REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => n247_port, D => n374, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => n247_port, D => n377, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => n252_port, D => n284_port, 
                           Q => REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => n252_port, D => n287_port, 
                           Q => REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => n252_port, D => n290_port, 
                           Q => REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => n252_port, D => n293_port, 
                           Q => REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => n252_port, D => n296_port, 
                           Q => REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => n252_port, D => n299_port, 
                           Q => REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => n252_port, D => n302_port, 
                           Q => REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => n252_port, D => n305_port, 
                           Q => REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => n252_port, D => n308_port, 
                           Q => REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => n252_port, D => n311_port, 
                           Q => REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => n251_port, D => n314_port, 
                           Q => REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => n251_port, D => n317_port, 
                           Q => REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => n251_port, D => n320_port, 
                           Q => REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => n251_port, D => n323_port, 
                           Q => REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => n251_port, D => n326_port, 
                           Q => REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => n251_port, D => n329_port, 
                           Q => REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => n251_port, D => n332_port, 
                           Q => REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => n251_port, D => n335_port, 
                           Q => REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => n251_port, D => n338_port, 
                           Q => REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => n251_port, D => n341_port, 
                           Q => REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => n251_port, D => n344_port, 
                           Q => REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => n250_port, D => n347_port, 
                           Q => REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => n250_port, D => n350_port, Q
                           => REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => n250_port, D => n353_port, Q
                           => REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => n250_port, D => n356_port, Q
                           => REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => n250_port, D => n359_port, Q
                           => REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => n250_port, D => n362_port, Q
                           => REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => n250_port, D => n365_port, Q
                           => REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => n250_port, D => n368_port, Q
                           => REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => n250_port, D => n371_port, Q
                           => REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => n250_port, D => n374, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => n250_port, D => n377, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => n255_port, D => n284_port, 
                           Q => REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => n255_port, D => n287_port, 
                           Q => REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => n255_port, D => n290_port, 
                           Q => REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => n255_port, D => n293_port, 
                           Q => REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => n255_port, D => n296_port, 
                           Q => REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => n255_port, D => n299_port, 
                           Q => REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => n255_port, D => n302_port, 
                           Q => REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => n255_port, D => n305_port, 
                           Q => REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => n255_port, D => n308_port, 
                           Q => REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => n255_port, D => n311_port, 
                           Q => REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => n254_port, D => n314_port, 
                           Q => REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => n254_port, D => n317_port, 
                           Q => REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => n254_port, D => n320_port, 
                           Q => REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => n254_port, D => n323_port, 
                           Q => REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => n254_port, D => n326_port, 
                           Q => REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => n254_port, D => n329_port, 
                           Q => REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => n254_port, D => n332_port, 
                           Q => REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => n254_port, D => n335_port, 
                           Q => REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => n254_port, D => n338_port, 
                           Q => REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => n254_port, D => n341_port, 
                           Q => REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => n254_port, D => n344_port, 
                           Q => REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => n253_port, D => n347_port, 
                           Q => REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => n253_port, D => n350_port, Q
                           => REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => n253_port, D => n353_port, Q
                           => REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => n253_port, D => n356_port, Q
                           => REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => n253_port, D => n359_port, Q
                           => REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => n253_port, D => n362_port, Q
                           => REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => n253_port, D => n365_port, Q
                           => REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => n253_port, D => n368_port, Q
                           => REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => n253_port, D => n371_port, Q
                           => REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => n253_port, D => n374, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => n253_port, D => n377, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => n258_port, D => n284_port, 
                           Q => REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => n258_port, D => n287_port, 
                           Q => REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => n258_port, D => n290_port, 
                           Q => REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => n258_port, D => n293_port, 
                           Q => REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => n258_port, D => n296_port, 
                           Q => REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => n258_port, D => n299_port, 
                           Q => REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => n258_port, D => n302_port, 
                           Q => REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => n258_port, D => n305_port, 
                           Q => REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => n258_port, D => n308_port, 
                           Q => REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => n258_port, D => n311_port, 
                           Q => REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => n257_port, D => n314_port, 
                           Q => REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => n257_port, D => n317_port, 
                           Q => REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => n257_port, D => n320_port, 
                           Q => REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => n257_port, D => n323_port, 
                           Q => REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => n257_port, D => n326_port, 
                           Q => REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => n257_port, D => n329_port, 
                           Q => REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => n257_port, D => n332_port, 
                           Q => REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => n257_port, D => n335_port, 
                           Q => REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => n257_port, D => n338_port, 
                           Q => REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => n257_port, D => n341_port, 
                           Q => REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => n257_port, D => n344_port, 
                           Q => REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => n256_port, D => n347_port, 
                           Q => REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => n256_port, D => n350_port, Q
                           => REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => n256_port, D => n353_port, Q
                           => REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => n256_port, D => n356_port, Q
                           => REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => n256_port, D => n359_port, Q
                           => REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => n256_port, D => n362_port, Q
                           => REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => n256_port, D => n365_port, Q
                           => REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => n256_port, D => n368_port, Q
                           => REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => n256_port, D => n371_port, Q
                           => REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => n256_port, D => n374, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => n256_port, D => n377, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => n261_port, D => n285_port, 
                           Q => REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => n261_port, D => n288_port, 
                           Q => REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => n261_port, D => n291_port, 
                           Q => REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => n261_port, D => n294_port, 
                           Q => REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => n261_port, D => n297_port, 
                           Q => REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => n261_port, D => n300_port, 
                           Q => REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => n261_port, D => n303_port, 
                           Q => REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => n261_port, D => n306, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => n261_port, D => n309_port, 
                           Q => REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => n261_port, D => n312_port, 
                           Q => REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => n260_port, D => n315_port, 
                           Q => REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => n260_port, D => n318_port, 
                           Q => REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => n260_port, D => n321_port, 
                           Q => REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => n260_port, D => n324_port, 
                           Q => REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => n260_port, D => n327_port, 
                           Q => REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => n260_port, D => n330_port, 
                           Q => REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => n260_port, D => n333_port, 
                           Q => REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => n260_port, D => n336_port, 
                           Q => REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => n260_port, D => n339_port, 
                           Q => REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => n260_port, D => n342_port, 
                           Q => REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => n260_port, D => n345_port, 
                           Q => REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => n259_port, D => n348_port, 
                           Q => REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => n259_port, D => n351_port, Q
                           => REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => n259_port, D => n354_port, Q
                           => REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => n259_port, D => n357_port, Q
                           => REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => n259_port, D => n360_port, Q
                           => REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => n259_port, D => n363_port, Q
                           => REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => n259_port, D => n366_port, Q
                           => REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => n259_port, D => n369_port, Q
                           => REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => n259_port, D => n372, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => n259_port, D => n375, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => n259_port, D => n378, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => n264_port, D => n285_port, 
                           Q => REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => n264_port, D => n288_port, 
                           Q => REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => n264_port, D => n291_port, 
                           Q => REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => n264_port, D => n294_port, 
                           Q => REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => n264_port, D => n297_port, 
                           Q => REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => n264_port, D => n300_port, 
                           Q => REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => n264_port, D => n303_port, 
                           Q => REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => n264_port, D => n306, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => n264_port, D => n309_port, 
                           Q => REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => n264_port, D => n312_port, 
                           Q => REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => n263_port, D => n315_port, 
                           Q => REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => n263_port, D => n318_port, 
                           Q => REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => n263_port, D => n321_port, 
                           Q => REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => n263_port, D => n324_port, 
                           Q => REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => n263_port, D => n327_port, 
                           Q => REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => n263_port, D => n330_port, 
                           Q => REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => n263_port, D => n333_port, 
                           Q => REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => n263_port, D => n336_port, 
                           Q => REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => n263_port, D => n339_port, 
                           Q => REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => n263_port, D => n342_port, 
                           Q => REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => n263_port, D => n345_port, 
                           Q => REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => n262_port, D => n348_port, 
                           Q => REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => n262_port, D => n351_port, Q
                           => REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => n262_port, D => n354_port, Q
                           => REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => n262_port, D => n357_port, Q
                           => REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => n262_port, D => n360_port, Q
                           => REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => n262_port, D => n363_port, Q
                           => REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => n262_port, D => n366_port, Q
                           => REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => n262_port, D => n369_port, Q
                           => REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => n262_port, D => n372, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => n262_port, D => n375, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => n262_port, D => n378, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => n267_port, D => n285_port, 
                           Q => REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => n267_port, D => n288_port, 
                           Q => REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => n267_port, D => n291_port, 
                           Q => REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => n267_port, D => n294_port, 
                           Q => REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => n267_port, D => n297_port, 
                           Q => REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => n267_port, D => n300_port, 
                           Q => REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => n267_port, D => n303_port, 
                           Q => REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => n267_port, D => n306, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => n267_port, D => n309_port, 
                           Q => REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => n267_port, D => n312_port, 
                           Q => REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => n266_port, D => n315_port, 
                           Q => REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => n266_port, D => n318_port, 
                           Q => REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => n266_port, D => n321_port, 
                           Q => REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => n266_port, D => n324_port, 
                           Q => REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => n266_port, D => n327_port, 
                           Q => REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => n266_port, D => n330_port, 
                           Q => REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => n266_port, D => n333_port, 
                           Q => REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => n266_port, D => n336_port, 
                           Q => REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => n266_port, D => n339_port, 
                           Q => REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => n266_port, D => n342_port, 
                           Q => REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => n266_port, D => n345_port, 
                           Q => REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => n265_port, D => n348_port, 
                           Q => REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => n265_port, D => n351_port, Q
                           => REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => n265_port, D => n354_port, Q
                           => REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => n265_port, D => n357_port, Q
                           => REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => n265_port, D => n360_port, Q
                           => REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => n265_port, D => n363_port, Q
                           => REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => n265_port, D => n366_port, Q
                           => REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => n265_port, D => n369_port, Q
                           => REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => n265_port, D => n372, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => n265_port, D => n375, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => n265_port, D => n378, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => n270_port, D => n285_port, 
                           Q => REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => n270_port, D => n288_port, 
                           Q => REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => n270_port, D => n291_port, 
                           Q => REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => n270_port, D => n294_port, 
                           Q => REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => n270_port, D => n297_port, 
                           Q => REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => n270_port, D => n300_port, 
                           Q => REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => n270_port, D => n303_port, 
                           Q => REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => n270_port, D => n306, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => n270_port, D => n309_port, 
                           Q => REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => n270_port, D => n312_port, 
                           Q => REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => n269_port, D => n315_port, 
                           Q => REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => n269_port, D => n318_port, 
                           Q => REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => n269_port, D => n321_port, 
                           Q => REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => n269_port, D => n324_port, 
                           Q => REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => n269_port, D => n327_port, 
                           Q => REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => n269_port, D => n330_port, 
                           Q => REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => n269_port, D => n333_port, 
                           Q => REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => n269_port, D => n336_port, 
                           Q => REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => n269_port, D => n339_port, 
                           Q => REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => n269_port, D => n342_port, 
                           Q => REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => n269_port, D => n345_port, 
                           Q => REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => n268_port, D => n348_port, 
                           Q => REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => n268_port, D => n351_port, Q
                           => REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => n268_port, D => n354_port, Q
                           => REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => n268_port, D => n357_port, Q
                           => REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => n268_port, D => n360_port, Q
                           => REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => n268_port, D => n363_port, Q
                           => REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => n268_port, D => n366_port, Q
                           => REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => n268_port, D => n369_port, Q
                           => REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => n268_port, D => n372, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => n268_port, D => n375, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => n268_port, D => n378, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => n273_port, D => n285_port, 
                           Q => REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => n273_port, D => n288_port, 
                           Q => REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => n273_port, D => n291_port, 
                           Q => REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => n273_port, D => n294_port, 
                           Q => REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => n273_port, D => n297_port, 
                           Q => REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => n273_port, D => n300_port, 
                           Q => REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => n273_port, D => n303_port, 
                           Q => REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => n273_port, D => n306, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => n273_port, D => n309_port, 
                           Q => REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => n273_port, D => n312_port, 
                           Q => REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => n272_port, D => n315_port, 
                           Q => REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => n272_port, D => n318_port, 
                           Q => REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => n272_port, D => n321_port, 
                           Q => REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => n272_port, D => n324_port, 
                           Q => REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => n272_port, D => n327_port, 
                           Q => REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => n272_port, D => n330_port, 
                           Q => REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => n272_port, D => n333_port, 
                           Q => REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => n272_port, D => n336_port, 
                           Q => REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => n272_port, D => n339_port, 
                           Q => REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => n272_port, D => n342_port, 
                           Q => REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => n272_port, D => n345_port, 
                           Q => REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => n271_port, D => n348_port, 
                           Q => REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => n271_port, D => n351_port, Q
                           => REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => n271_port, D => n354_port, Q
                           => REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => n271_port, D => n357_port, Q
                           => REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => n271_port, D => n360_port, Q
                           => REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => n271_port, D => n363_port, Q
                           => REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => n271_port, D => n366_port, Q
                           => REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => n271_port, D => n369_port, Q
                           => REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => n271_port, D => n372, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => n271_port, D => n375, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => n271_port, D => n378, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => n276_port, D => n285_port, 
                           Q => REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => n276_port, D => n288_port, 
                           Q => REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => n276_port, D => n291_port, 
                           Q => REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => n276_port, D => n294_port, 
                           Q => REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => n276_port, D => n297_port, 
                           Q => REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => n276_port, D => n300_port, 
                           Q => REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => n276_port, D => n303_port, 
                           Q => REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => n276_port, D => n306, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => n276_port, D => n309_port, 
                           Q => REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => n276_port, D => n312_port, 
                           Q => REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => n275_port, D => n315_port, 
                           Q => REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => n275_port, D => n318_port, 
                           Q => REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => n275_port, D => n321_port, 
                           Q => REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => n275_port, D => n324_port, 
                           Q => REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => n275_port, D => n327_port, 
                           Q => REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => n275_port, D => n330_port, 
                           Q => REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => n275_port, D => n333_port, 
                           Q => REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => n275_port, D => n336_port, 
                           Q => REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => n275_port, D => n339_port, 
                           Q => REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => n275_port, D => n342_port, 
                           Q => REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => n275_port, D => n345_port, 
                           Q => REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => n274_port, D => n348_port, 
                           Q => REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => n274_port, D => n351_port, Q
                           => REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => n274_port, D => n354_port, Q
                           => REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => n274_port, D => n357_port, Q
                           => REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => n274_port, D => n360_port, Q
                           => REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => n274_port, D => n363_port, Q
                           => REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => n274_port, D => n366_port, Q
                           => REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => n274_port, D => n369_port, Q
                           => REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => n274_port, D => n372, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => n274_port, D => n375, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => n274_port, D => n378, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => n279_port, D => n285_port, 
                           Q => REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => n279_port, D => n288_port, 
                           Q => REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => n279_port, D => n291_port, 
                           Q => REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => n279_port, D => n294_port, 
                           Q => REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => n279_port, D => n297_port, 
                           Q => REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => n279_port, D => n300_port, 
                           Q => REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => n279_port, D => n303_port, 
                           Q => REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => n279_port, D => n306, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => n279_port, D => n309_port, 
                           Q => REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => n279_port, D => n312_port, 
                           Q => REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => n278_port, D => n315_port, 
                           Q => REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => n278_port, D => n318_port, 
                           Q => REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => n278_port, D => n321_port, 
                           Q => REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => n278_port, D => n324_port, 
                           Q => REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => n278_port, D => n327_port, 
                           Q => REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => n278_port, D => n330_port, 
                           Q => REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => n278_port, D => n333_port, 
                           Q => REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => n278_port, D => n336_port, 
                           Q => REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => n278_port, D => n339_port, 
                           Q => REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => n278_port, D => n342_port, 
                           Q => REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => n278_port, D => n345_port, 
                           Q => REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => n277_port, D => n348_port, 
                           Q => REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => n277_port, D => n351_port, Q
                           => REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => n277_port, D => n354_port, Q
                           => REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => n277_port, D => n357_port, Q
                           => REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => n277_port, D => n360_port, Q
                           => REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => n277_port, D => n363_port, Q
                           => REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => n277_port, D => n366_port, Q
                           => REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => n277_port, D => n369_port, Q
                           => REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => n277_port, D => n372, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => n277_port, D => n375, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => n277_port, D => n378, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => n282_port, D => n285_port, 
                           Q => REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => n282_port, D => n288_port, 
                           Q => REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => n282_port, D => n291_port, 
                           Q => REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => n282_port, D => n294_port, 
                           Q => REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => n282_port, D => n297_port, 
                           Q => REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => n282_port, D => n300_port, 
                           Q => REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => n282_port, D => n303_port, 
                           Q => REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => n282_port, D => n306, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => n282_port, D => n309_port, 
                           Q => REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => n282_port, D => n312_port, 
                           Q => REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => n281_port, D => n315_port, 
                           Q => REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => n281_port, D => n318_port, 
                           Q => REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => n281_port, D => n321_port, 
                           Q => REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => n281_port, D => n324_port, 
                           Q => REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => n281_port, D => n327_port, 
                           Q => REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => n281_port, D => n330_port, 
                           Q => REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => n281_port, D => n333_port, 
                           Q => REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => n281_port, D => n336_port, 
                           Q => REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => n281_port, D => n339_port, 
                           Q => REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => n281_port, D => n342_port, 
                           Q => REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => n281_port, D => n345_port, 
                           Q => REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => n280_port, D => n348_port, 
                           Q => REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => n280_port, D => n351_port, Q
                           => REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => n280_port, D => n354_port, Q
                           => REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => n280_port, D => n357_port, Q
                           => REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => n280_port, D => n360_port, Q
                           => REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => n280_port, D => n363_port, Q
                           => REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => n280_port, D => n366_port, Q
                           => REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => n280_port, D => n369_port, Q
                           => REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => n280_port, D => n372, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => n280_port, D => n375, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => n280_port, D => n378, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => n381, D => n285_port, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => n381, D => n288_port, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => n381, D => n291_port, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => n381, D => n294_port, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => n381, D => n297_port, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => n381, D => n300_port, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => n381, D => n303_port, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => n381, D => n306, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => n381, D => n309_port, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => n381, D => n312_port, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => n380, D => n315_port, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => n380, D => n318_port, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => n380, D => n321_port, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => n380, D => n324_port, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => n380, D => n327_port, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => n380, D => n330_port, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => n380, D => n333_port, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => n380, D => n336_port, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => n380, D => n339_port, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => n380, D => n342_port, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => n380, D => n345_port, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => n379, D => n348_port, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => n379, D => n351_port, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => n379, D => n354_port, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => n379, D => n357_port, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => n379, D => n360_port, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => n379, D => n363_port, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => n379, D => n366_port, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => n379, D => n369_port, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => n379, D => n372, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => n379, D => n375, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => n379, D => n378, Q => 
                           REGISTERS_31_0_port);
   OUTA_reg_31_inst : DLH_X1 port map( G => n187, D => N339, Q => OUTA(31));
   OUTA_reg_30_inst : DLH_X1 port map( G => n187, D => N338, Q => OUTA(30));
   OUTA_reg_29_inst : DLH_X1 port map( G => n187, D => N337, Q => OUTA(29));
   OUTA_reg_28_inst : DLH_X1 port map( G => n187, D => N336, Q => OUTA(28));
   OUTA_reg_27_inst : DLH_X1 port map( G => n187, D => N335, Q => OUTA(27));
   OUTA_reg_26_inst : DLH_X1 port map( G => n187, D => N334, Q => OUTA(26));
   OUTA_reg_25_inst : DLH_X1 port map( G => n187, D => N333, Q => OUTA(25));
   OUTA_reg_24_inst : DLH_X1 port map( G => n187, D => N332, Q => OUTA(24));
   OUTA_reg_23_inst : DLH_X1 port map( G => n187, D => N331, Q => OUTA(23));
   OUTA_reg_22_inst : DLH_X1 port map( G => n187, D => N330, Q => OUTA(22));
   OUTA_reg_21_inst : DLH_X1 port map( G => n187, D => N329, Q => OUTA(21));
   OUTA_reg_20_inst : DLH_X1 port map( G => n188, D => N328, Q => OUTA(20));
   OUTA_reg_19_inst : DLH_X1 port map( G => n188, D => N327, Q => OUTA(19));
   OUTA_reg_18_inst : DLH_X1 port map( G => n188, D => N326, Q => OUTA(18));
   OUTA_reg_17_inst : DLH_X1 port map( G => n188, D => N325, Q => OUTA(17));
   OUTA_reg_16_inst : DLH_X1 port map( G => n188, D => N324, Q => OUTA(16));
   OUTA_reg_15_inst : DLH_X1 port map( G => n188, D => N323, Q => OUTA(15));
   OUTA_reg_14_inst : DLH_X1 port map( G => n188, D => N322, Q => OUTA(14));
   OUTA_reg_13_inst : DLH_X1 port map( G => n188, D => N321, Q => OUTA(13));
   OUTA_reg_12_inst : DLH_X1 port map( G => n188, D => N320, Q => OUTA(12));
   OUTA_reg_11_inst : DLH_X1 port map( G => n188, D => N319, Q => OUTA(11));
   OUTA_reg_10_inst : DLH_X1 port map( G => n188, D => N318, Q => OUTA(10));
   OUTA_reg_9_inst : DLH_X1 port map( G => n189, D => N317, Q => OUTA(9));
   OUTA_reg_8_inst : DLH_X1 port map( G => n189, D => N316, Q => OUTA(8));
   OUTA_reg_7_inst : DLH_X1 port map( G => n189, D => N315, Q => OUTA(7));
   OUTA_reg_6_inst : DLH_X1 port map( G => n189, D => N314, Q => OUTA(6));
   OUTA_reg_5_inst : DLH_X1 port map( G => n189, D => N313, Q => OUTA(5));
   OUTA_reg_4_inst : DLH_X1 port map( G => n189, D => N312, Q => OUTA(4));
   OUTA_reg_3_inst : DLH_X1 port map( G => n189, D => N311, Q => OUTA(3));
   OUTA_reg_2_inst : DLH_X1 port map( G => n189, D => N310, Q => OUTA(2));
   OUTA_reg_1_inst : DLH_X1 port map( G => n189, D => N309, Q => OUTA(1));
   OUTA_reg_0_inst : DLH_X1 port map( G => n189, D => N308, Q => OUTA(0));
   OUTB_reg_31_inst : DLH_X1 port map( G => n189, D => N371, Q => OUTB(31));
   OUTB_reg_30_inst : DLH_X1 port map( G => n190, D => N370, Q => OUTB(30));
   OUTB_reg_29_inst : DLH_X1 port map( G => n190, D => N369, Q => OUTB(29));
   OUTB_reg_28_inst : DLH_X1 port map( G => n190, D => N368, Q => OUTB(28));
   OUTB_reg_27_inst : DLH_X1 port map( G => n190, D => N367, Q => OUTB(27));
   OUTB_reg_26_inst : DLH_X1 port map( G => n190, D => N366, Q => OUTB(26));
   OUTB_reg_25_inst : DLH_X1 port map( G => n190, D => N365, Q => OUTB(25));
   OUTB_reg_24_inst : DLH_X1 port map( G => n190, D => N364, Q => OUTB(24));
   OUTB_reg_23_inst : DLH_X1 port map( G => n190, D => N363, Q => OUTB(23));
   OUTB_reg_22_inst : DLH_X1 port map( G => n190, D => N362, Q => OUTB(22));
   OUTB_reg_21_inst : DLH_X1 port map( G => n190, D => N361, Q => OUTB(21));
   OUTB_reg_20_inst : DLH_X1 port map( G => n190, D => N360, Q => OUTB(20));
   OUTB_reg_19_inst : DLH_X1 port map( G => n191, D => N359, Q => OUTB(19));
   OUTB_reg_18_inst : DLH_X1 port map( G => n191, D => N358, Q => OUTB(18));
   OUTB_reg_17_inst : DLH_X1 port map( G => n191, D => N357, Q => OUTB(17));
   OUTB_reg_16_inst : DLH_X1 port map( G => n191, D => N356, Q => OUTB(16));
   OUTB_reg_15_inst : DLH_X1 port map( G => n191, D => N355, Q => OUTB(15));
   OUTB_reg_14_inst : DLH_X1 port map( G => n191, D => N354, Q => OUTB(14));
   OUTB_reg_13_inst : DLH_X1 port map( G => n191, D => N353, Q => OUTB(13));
   OUTB_reg_12_inst : DLH_X1 port map( G => n191, D => N352, Q => OUTB(12));
   OUTB_reg_11_inst : DLH_X1 port map( G => n191, D => N351, Q => OUTB(11));
   OUTB_reg_10_inst : DLH_X1 port map( G => n191, D => N350, Q => OUTB(10));
   OUTB_reg_9_inst : DLH_X1 port map( G => n191, D => N349, Q => OUTB(9));
   OUTB_reg_8_inst : DLH_X1 port map( G => n192, D => N348, Q => OUTB(8));
   OUTB_reg_7_inst : DLH_X1 port map( G => n192, D => N347, Q => OUTB(7));
   OUTB_reg_6_inst : DLH_X1 port map( G => n192, D => N346, Q => OUTB(6));
   OUTB_reg_5_inst : DLH_X1 port map( G => n192, D => N345, Q => OUTB(5));
   OUTB_reg_4_inst : DLH_X1 port map( G => n192, D => N344, Q => OUTB(4));
   OUTB_reg_3_inst : DLH_X1 port map( G => n192, D => N343, Q => OUTB(3));
   OUTB_reg_2_inst : DLH_X1 port map( G => n192, D => N342, Q => OUTB(2));
   OUTB_reg_1_inst : DLH_X1 port map( G => n192, D => N341, Q => OUTB(1));
   OUTB_reg_0_inst : DLH_X1 port map( G => n192, D => N340, Q => OUTB(0));
   U1905 : NAND3_X1 port map( A1 => n408, A2 => n407, A3 => WE, ZN => n1775);
   U1906 : NAND3_X1 port map( A1 => WE, A2 => n407, A3 => ADD_WR(3), ZN => 
                           n1783);
   U1907 : NAND3_X1 port map( A1 => WE, A2 => n408, A3 => ADD_WR(4), ZN => 
                           n1785);
   U1908 : NAND3_X1 port map( A1 => n410, A2 => n409, A3 => n411, ZN => n1784);
   U1909 : NAND3_X1 port map( A1 => n410, A2 => n409, A3 => ADD_WR(0), ZN => 
                           n1776);
   U1910 : NAND3_X1 port map( A1 => n411, A2 => n409, A3 => ADD_WR(1), ZN => 
                           n1777);
   U1911 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n409, A3 => ADD_WR(1), ZN 
                           => n1778);
   U1912 : NAND3_X1 port map( A1 => n411, A2 => n410, A3 => ADD_WR(2), ZN => 
                           n1779);
   U1913 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n410, A3 => ADD_WR(2), ZN 
                           => n1780);
   U1914 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n411, A3 => ADD_WR(2), ZN 
                           => n1781);
   U1915 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => WE, A3 => ADD_WR(4), ZN =>
                           n1786);
   U1916 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n1782);
   U3 : NOR2_X1 port map( A1 => n2152, A2 => ADD_RDB(1), ZN => n1130);
   U4 : NOR2_X1 port map( A1 => n2155, A2 => ADD_RDA(1), ZN => n1754);
   U5 : BUF_X1 port map( A => n542, Z => n163);
   U6 : BUF_X1 port map( A => n566, Z => n118);
   U7 : BUF_X1 port map( A => n576, Z => n94);
   U8 : BUF_X1 port map( A => n542, Z => n164);
   U9 : BUF_X1 port map( A => n566, Z => n119);
   U10 : BUF_X1 port map( A => n576, Z => n95);
   U11 : BUF_X1 port map( A => n542, Z => n165);
   U12 : BUF_X1 port map( A => n566, Z => n120);
   U13 : BUF_X1 port map( A => n576, Z => n96);
   U14 : BUF_X1 port map( A => n549, Z => n145);
   U15 : BUF_X1 port map( A => n549, Z => n146);
   U16 : BUF_X1 port map( A => n549, Z => n147);
   U17 : BUF_X1 port map( A => n536, Z => n178);
   U18 : BUF_X1 port map( A => n541, Z => n166);
   U19 : BUF_X1 port map( A => n546, Z => n154);
   U20 : BUF_X1 port map( A => n551, Z => n142);
   U21 : BUF_X1 port map( A => n570, Z => n109);
   U22 : BUF_X1 port map( A => n565, Z => n121);
   U23 : BUF_X1 port map( A => n575, Z => n97);
   U24 : BUF_X1 port map( A => n560, Z => n133);
   U25 : BUF_X1 port map( A => n536, Z => n179);
   U26 : BUF_X1 port map( A => n541, Z => n167);
   U27 : BUF_X1 port map( A => n546, Z => n155);
   U28 : BUF_X1 port map( A => n551, Z => n143);
   U29 : BUF_X1 port map( A => n570, Z => n110);
   U30 : BUF_X1 port map( A => n565, Z => n122);
   U31 : BUF_X1 port map( A => n575, Z => n98);
   U32 : BUF_X1 port map( A => n560, Z => n134);
   U33 : BUF_X1 port map( A => n533, Z => n184);
   U34 : BUF_X1 port map( A => n538, Z => n172);
   U35 : BUF_X1 port map( A => n543, Z => n160);
   U36 : BUF_X1 port map( A => n548, Z => n148);
   U37 : BUF_X1 port map( A => n567, Z => n115);
   U38 : BUF_X1 port map( A => n562, Z => n127);
   U39 : BUF_X1 port map( A => n572, Z => n103);
   U40 : BUF_X1 port map( A => n533, Z => n185);
   U41 : BUF_X1 port map( A => n538, Z => n173);
   U42 : BUF_X1 port map( A => n543, Z => n161);
   U43 : BUF_X1 port map( A => n548, Z => n149);
   U44 : BUF_X1 port map( A => n567, Z => n116);
   U45 : BUF_X1 port map( A => n562, Z => n128);
   U46 : BUF_X1 port map( A => n572, Z => n104);
   U47 : BUF_X1 port map( A => n537, Z => n175);
   U48 : BUF_X1 port map( A => n547, Z => n151);
   U49 : BUF_X1 port map( A => n552, Z => n139);
   U50 : BUF_X1 port map( A => n571, Z => n106);
   U51 : BUF_X1 port map( A => n561, Z => n130);
   U52 : BUF_X1 port map( A => n537, Z => n176);
   U53 : BUF_X1 port map( A => n547, Z => n152);
   U54 : BUF_X1 port map( A => n552, Z => n140);
   U55 : BUF_X1 port map( A => n571, Z => n107);
   U56 : BUF_X1 port map( A => n561, Z => n131);
   U57 : BUF_X1 port map( A => n1173, Z => n52);
   U58 : BUF_X1 port map( A => n1173, Z => n53);
   U59 : BUF_X1 port map( A => n533, Z => n186);
   U60 : BUF_X1 port map( A => n538, Z => n174);
   U61 : BUF_X1 port map( A => n567, Z => n117);
   U62 : BUF_X1 port map( A => n562, Z => n129);
   U63 : BUF_X1 port map( A => n572, Z => n105);
   U64 : BUF_X1 port map( A => n536, Z => n180);
   U65 : BUF_X1 port map( A => n541, Z => n168);
   U66 : BUF_X1 port map( A => n546, Z => n156);
   U67 : BUF_X1 port map( A => n551, Z => n144);
   U68 : BUF_X1 port map( A => n570, Z => n111);
   U69 : BUF_X1 port map( A => n565, Z => n123);
   U70 : BUF_X1 port map( A => n575, Z => n99);
   U71 : BUF_X1 port map( A => n560, Z => n135);
   U72 : BUF_X1 port map( A => n543, Z => n162);
   U73 : BUF_X1 port map( A => n548, Z => n150);
   U74 : BUF_X1 port map( A => n557, Z => n136);
   U75 : BUF_X1 port map( A => n557, Z => n137);
   U76 : BUF_X1 port map( A => n537, Z => n177);
   U77 : BUF_X1 port map( A => n547, Z => n153);
   U78 : BUF_X1 port map( A => n552, Z => n141);
   U79 : BUF_X1 port map( A => n571, Z => n108);
   U80 : BUF_X1 port map( A => n561, Z => n132);
   U81 : BUF_X1 port map( A => n534, Z => n181);
   U82 : BUF_X1 port map( A => n539, Z => n169);
   U83 : BUF_X1 port map( A => n544, Z => n157);
   U84 : BUF_X1 port map( A => n568, Z => n112);
   U85 : BUF_X1 port map( A => n563, Z => n124);
   U86 : BUF_X1 port map( A => n573, Z => n100);
   U87 : BUF_X1 port map( A => n534, Z => n182);
   U88 : BUF_X1 port map( A => n539, Z => n170);
   U89 : BUF_X1 port map( A => n544, Z => n158);
   U90 : BUF_X1 port map( A => n568, Z => n113);
   U91 : BUF_X1 port map( A => n563, Z => n125);
   U92 : BUF_X1 port map( A => n573, Z => n101);
   U93 : BUF_X1 port map( A => n1166, Z => n71);
   U94 : BUF_X1 port map( A => n1190, Z => n26);
   U95 : BUF_X1 port map( A => n1200, Z => n2);
   U96 : BUF_X1 port map( A => n1166, Z => n70);
   U97 : BUF_X1 port map( A => n1190, Z => n25);
   U98 : BUF_X1 port map( A => n1200, Z => n1);
   U99 : BUF_X1 port map( A => n1173, Z => n54);
   U100 : BUF_X1 port map( A => n557, Z => n138);
   U101 : BUF_X1 port map( A => n534, Z => n183);
   U102 : BUF_X1 port map( A => n539, Z => n171);
   U103 : BUF_X1 port map( A => n568, Z => n114);
   U104 : BUF_X1 port map( A => n563, Z => n126);
   U105 : BUF_X1 port map( A => n573, Z => n102);
   U106 : BUF_X1 port map( A => n544, Z => n159);
   U107 : BUF_X1 port map( A => n1166, Z => n72);
   U108 : BUF_X1 port map( A => n1190, Z => n27);
   U109 : BUF_X1 port map( A => n1200, Z => n3);
   U110 : NAND2_X1 port map( A1 => n1133, A2 => n1129, ZN => n549);
   U111 : AND2_X1 port map( A1 => n1124, A2 => n1129, ZN => n542);
   U112 : AND2_X1 port map( A1 => n1142, A2 => n1129, ZN => n566);
   U113 : AND2_X1 port map( A1 => n1147, A2 => n1129, ZN => n576);
   U114 : INV_X1 port map( A => n406, ZN => n390);
   U115 : INV_X1 port map( A => n406, ZN => n389);
   U116 : INV_X1 port map( A => n406, ZN => n393);
   U117 : INV_X1 port map( A => n406, ZN => n392);
   U118 : INV_X1 port map( A => n406, ZN => n391);
   U119 : NOR2_X1 port map( A1 => n2152, A2 => n2151, ZN => n1129);
   U120 : BUF_X1 port map( A => n1181, Z => n43);
   U121 : BUF_X1 port map( A => n1181, Z => n44);
   U122 : BUF_X1 port map( A => n1158, Z => n88);
   U123 : BUF_X1 port map( A => n1163, Z => n76);
   U124 : BUF_X1 port map( A => n1168, Z => n64);
   U125 : BUF_X1 port map( A => n1187, Z => n31);
   U126 : BUF_X1 port map( A => n1192, Z => n19);
   U127 : BUF_X1 port map( A => n1197, Z => n7);
   U128 : BUF_X1 port map( A => n1158, Z => n89);
   U129 : BUF_X1 port map( A => n1163, Z => n77);
   U130 : BUF_X1 port map( A => n1168, Z => n65);
   U131 : BUF_X1 port map( A => n1187, Z => n32);
   U132 : BUF_X1 port map( A => n1192, Z => n20);
   U133 : BUF_X1 port map( A => n1197, Z => n8);
   U134 : BUF_X1 port map( A => n1160, Z => n85);
   U135 : BUF_X1 port map( A => n1165, Z => n73);
   U136 : BUF_X1 port map( A => n1170, Z => n61);
   U137 : BUF_X1 port map( A => n1175, Z => n49);
   U138 : BUF_X1 port map( A => n1189, Z => n28);
   U139 : BUF_X1 port map( A => n1194, Z => n16);
   U140 : BUF_X1 port map( A => n1184, Z => n40);
   U141 : BUF_X1 port map( A => n1199, Z => n4);
   U142 : BUF_X1 port map( A => n1160, Z => n86);
   U143 : BUF_X1 port map( A => n1165, Z => n74);
   U144 : BUF_X1 port map( A => n1170, Z => n62);
   U145 : BUF_X1 port map( A => n1175, Z => n50);
   U146 : BUF_X1 port map( A => n1189, Z => n29);
   U147 : BUF_X1 port map( A => n1194, Z => n17);
   U148 : BUF_X1 port map( A => n1184, Z => n41);
   U149 : BUF_X1 port map( A => n1199, Z => n5);
   U150 : BUF_X1 port map( A => n1157, Z => n91);
   U151 : BUF_X1 port map( A => n1162, Z => n79);
   U152 : BUF_X1 port map( A => n1167, Z => n67);
   U153 : BUF_X1 port map( A => n1172, Z => n55);
   U154 : BUF_X1 port map( A => n1186, Z => n34);
   U155 : BUF_X1 port map( A => n1191, Z => n22);
   U156 : BUF_X1 port map( A => n1196, Z => n10);
   U157 : BUF_X1 port map( A => n1157, Z => n92);
   U158 : BUF_X1 port map( A => n1162, Z => n80);
   U159 : BUF_X1 port map( A => n1167, Z => n68);
   U160 : BUF_X1 port map( A => n1172, Z => n56);
   U161 : BUF_X1 port map( A => n1186, Z => n35);
   U162 : BUF_X1 port map( A => n1191, Z => n23);
   U163 : BUF_X1 port map( A => n1196, Z => n11);
   U164 : BUF_X1 port map( A => n1181, Z => n45);
   U165 : BUF_X1 port map( A => n1161, Z => n83);
   U166 : BUF_X1 port map( A => n1171, Z => n59);
   U167 : BUF_X1 port map( A => n1176, Z => n47);
   U168 : BUF_X1 port map( A => n1195, Z => n14);
   U169 : BUF_X1 port map( A => n1185, Z => n38);
   U170 : BUF_X1 port map( A => n1161, Z => n82);
   U171 : BUF_X1 port map( A => n1171, Z => n58);
   U172 : BUF_X1 port map( A => n1176, Z => n46);
   U173 : BUF_X1 port map( A => n1195, Z => n13);
   U174 : BUF_X1 port map( A => n1185, Z => n37);
   U175 : BUF_X1 port map( A => n1158, Z => n90);
   U176 : BUF_X1 port map( A => n1163, Z => n78);
   U177 : BUF_X1 port map( A => n1168, Z => n66);
   U178 : BUF_X1 port map( A => n1187, Z => n33);
   U179 : BUF_X1 port map( A => n1192, Z => n21);
   U180 : BUF_X1 port map( A => n1197, Z => n9);
   U181 : BUF_X1 port map( A => n1160, Z => n87);
   U182 : BUF_X1 port map( A => n1165, Z => n75);
   U183 : BUF_X1 port map( A => n1170, Z => n63);
   U184 : BUF_X1 port map( A => n1175, Z => n51);
   U185 : BUF_X1 port map( A => n1189, Z => n30);
   U186 : BUF_X1 port map( A => n1194, Z => n18);
   U187 : BUF_X1 port map( A => n1184, Z => n42);
   U188 : BUF_X1 port map( A => n1199, Z => n6);
   U189 : BUF_X1 port map( A => n1157, Z => n93);
   U190 : BUF_X1 port map( A => n1162, Z => n81);
   U191 : BUF_X1 port map( A => n1167, Z => n69);
   U192 : BUF_X1 port map( A => n1172, Z => n57);
   U193 : BUF_X1 port map( A => n1186, Z => n36);
   U194 : BUF_X1 port map( A => n1191, Z => n24);
   U195 : BUF_X1 port map( A => n1196, Z => n12);
   U196 : BUF_X1 port map( A => n1176, Z => n48);
   U197 : BUF_X1 port map( A => n1161, Z => n84);
   U198 : BUF_X1 port map( A => n1171, Z => n60);
   U199 : BUF_X1 port map( A => n1195, Z => n15);
   U200 : BUF_X1 port map( A => n1185, Z => n39);
   U201 : NAND2_X1 port map( A1 => n1127, A2 => n1134, ZN => n543);
   U202 : NAND2_X1 port map( A1 => n1127, A2 => n1133, ZN => n544);
   U203 : NAND2_X1 port map( A1 => n1129, A2 => n1134, ZN => n548);
   U204 : NAND2_X1 port map( A1 => n1126, A2 => n1130, ZN => n538);
   U205 : NAND2_X1 port map( A1 => n1124, A2 => n1130, ZN => n539);
   U206 : NAND2_X1 port map( A1 => n1143, A2 => n1130, ZN => n562);
   U207 : NAND2_X1 port map( A1 => n1142, A2 => n1130, ZN => n563);
   U208 : NAND2_X1 port map( A1 => n1148, A2 => n1130, ZN => n572);
   U209 : NAND2_X1 port map( A1 => n1147, A2 => n1130, ZN => n573);
   U210 : NAND2_X1 port map( A1 => n1126, A2 => n1127, ZN => n533);
   U211 : NAND2_X1 port map( A1 => n1124, A2 => n1127, ZN => n534);
   U212 : NAND2_X1 port map( A1 => n1148, A2 => n1127, ZN => n567);
   U213 : NAND2_X1 port map( A1 => n1147, A2 => n1127, ZN => n568);
   U214 : NAND2_X1 port map( A1 => n1143, A2 => n1127, ZN => n557);
   U215 : AND2_X1 port map( A1 => n1136, A2 => n2150, ZN => n1133);
   U216 : NAND2_X1 port map( A1 => n1757, A2 => n1753, ZN => n1173);
   U217 : AND2_X1 port map( A1 => n1150, A2 => n2150, ZN => n1147);
   U218 : AND2_X1 port map( A1 => n1131, A2 => n2150, ZN => n1124);
   U219 : AND2_X1 port map( A1 => n1130, A2 => n1133, ZN => n552);
   U220 : AND2_X1 port map( A1 => n1130, A2 => n1134, ZN => n551);
   U221 : AND2_X1 port map( A1 => n1125, A2 => n1133, ZN => n547);
   U222 : AND2_X1 port map( A1 => n1125, A2 => n1134, ZN => n546);
   U223 : AND2_X1 port map( A1 => n1126, A2 => n1129, ZN => n541);
   U224 : AND2_X1 port map( A1 => n1143, A2 => n1129, ZN => n565);
   U225 : AND2_X1 port map( A1 => n1148, A2 => n1129, ZN => n575);
   U226 : AND2_X1 port map( A1 => n1748, A2 => n1753, ZN => n1166);
   U227 : AND2_X1 port map( A1 => n1766, A2 => n1753, ZN => n1190);
   U228 : AND2_X1 port map( A1 => n1771, A2 => n1753, ZN => n1200);
   U229 : AND2_X1 port map( A1 => n1124, A2 => n1125, ZN => n537);
   U230 : AND2_X1 port map( A1 => n1126, A2 => n1125, ZN => n536);
   U231 : AND2_X1 port map( A1 => n1147, A2 => n1125, ZN => n571);
   U232 : AND2_X1 port map( A1 => n1148, A2 => n1125, ZN => n570);
   U233 : AND2_X1 port map( A1 => n1142, A2 => n1125, ZN => n561);
   U234 : AND2_X1 port map( A1 => n1143, A2 => n1125, ZN => n560);
   U235 : AND2_X1 port map( A1 => n1145, A2 => n2150, ZN => n1142);
   U236 : BUF_X1 port map( A => n386, Z => n406);
   U237 : BUF_X1 port map( A => n385, Z => n405);
   U238 : BUF_X1 port map( A => n385, Z => n404);
   U239 : BUF_X1 port map( A => n385, Z => n403);
   U240 : BUF_X1 port map( A => n384, Z => n402);
   U241 : BUF_X1 port map( A => n384, Z => n401);
   U242 : BUF_X1 port map( A => n384, Z => n400);
   U243 : BUF_X1 port map( A => n383, Z => n399);
   U244 : BUF_X1 port map( A => n383, Z => n397);
   U245 : BUF_X1 port map( A => n382, Z => n396);
   U246 : BUF_X1 port map( A => n382, Z => n395);
   U247 : BUF_X1 port map( A => n382, Z => n394);
   U248 : BUF_X1 port map( A => n383, Z => n398);
   U249 : NOR2_X1 port map( A1 => ADD_RDB(1), A2 => ADD_RDB(2), ZN => n1127);
   U250 : NOR2_X1 port map( A1 => n2155, A2 => n2156, ZN => n1753);
   U251 : NOR2_X1 port map( A1 => n2151, A2 => ADD_RDB(2), ZN => n1125);
   U252 : NAND2_X1 port map( A1 => n1751, A2 => n1757, ZN => n1168);
   U253 : NAND2_X1 port map( A1 => n1751, A2 => n1758, ZN => n1167);
   U254 : NAND2_X1 port map( A1 => n1753, A2 => n1758, ZN => n1172);
   U255 : NAND2_X1 port map( A1 => n1750, A2 => n1754, ZN => n1162);
   U256 : NAND2_X1 port map( A1 => n1748, A2 => n1754, ZN => n1163);
   U257 : NAND2_X1 port map( A1 => n1767, A2 => n1754, ZN => n1186);
   U258 : NAND2_X1 port map( A1 => n1766, A2 => n1754, ZN => n1187);
   U259 : NAND2_X1 port map( A1 => n1772, A2 => n1754, ZN => n1196);
   U260 : NAND2_X1 port map( A1 => n1771, A2 => n1754, ZN => n1197);
   U261 : NAND2_X1 port map( A1 => n1750, A2 => n1751, ZN => n1157);
   U262 : NAND2_X1 port map( A1 => n1748, A2 => n1751, ZN => n1158);
   U263 : NAND2_X1 port map( A1 => n1771, A2 => n1751, ZN => n1192);
   U264 : NAND2_X1 port map( A1 => n1772, A2 => n1751, ZN => n1191);
   U265 : NAND2_X1 port map( A1 => n1767, A2 => n1751, ZN => n1181);
   U266 : AND2_X1 port map( A1 => ADD_RDB(0), A2 => n1136, ZN => n1134);
   U267 : AND2_X1 port map( A1 => n1760, A2 => n2157, ZN => n1757);
   U268 : NOR2_X1 port map( A1 => ADD_RDB(3), A2 => ADD_RDB(4), ZN => n1145);
   U269 : NOR2_X1 port map( A1 => n2153, A2 => ADD_RDB(4), ZN => n1150);
   U270 : AND2_X1 port map( A1 => n1131, A2 => ADD_RDB(0), ZN => n1126);
   U271 : AND2_X1 port map( A1 => n1150, A2 => ADD_RDB(0), ZN => n1148);
   U272 : AND2_X1 port map( A1 => n1145, A2 => ADD_RDB(0), ZN => n1143);
   U273 : AND2_X1 port map( A1 => n1774, A2 => n2157, ZN => n1771);
   U274 : AND2_X1 port map( A1 => n1755, A2 => n2157, ZN => n1748);
   U275 : AND2_X1 port map( A1 => n1754, A2 => n1757, ZN => n1176);
   U276 : AND2_X1 port map( A1 => n1754, A2 => n1758, ZN => n1175);
   U277 : AND2_X1 port map( A1 => n1749, A2 => n1757, ZN => n1171);
   U278 : AND2_X1 port map( A1 => n1749, A2 => n1758, ZN => n1170);
   U279 : AND2_X1 port map( A1 => n1750, A2 => n1753, ZN => n1165);
   U280 : AND2_X1 port map( A1 => n1767, A2 => n1753, ZN => n1189);
   U281 : AND2_X1 port map( A1 => n1772, A2 => n1753, ZN => n1199);
   U282 : AND2_X1 port map( A1 => n1750, A2 => n1749, ZN => n1160);
   U283 : AND2_X1 port map( A1 => n1748, A2 => n1749, ZN => n1161);
   U284 : AND2_X1 port map( A1 => n1771, A2 => n1749, ZN => n1195);
   U285 : AND2_X1 port map( A1 => n1772, A2 => n1749, ZN => n1194);
   U286 : AND2_X1 port map( A1 => n1766, A2 => n1749, ZN => n1185);
   U287 : AND2_X1 port map( A1 => n1767, A2 => n1749, ZN => n1184);
   U288 : INV_X1 port map( A => ADD_RDB(0), ZN => n2150);
   U289 : AND2_X1 port map( A1 => n1769, A2 => n2157, ZN => n1766);
   U290 : INV_X1 port map( A => ADD_RDB(1), ZN => n2151);
   U291 : INV_X1 port map( A => ADD_RDB(2), ZN => n2152);
   U292 : AND2_X1 port map( A1 => ADD_RDB(4), A2 => ADD_RDB(3), ZN => n1136);
   U293 : AND2_X1 port map( A1 => ADD_RDB(4), A2 => n2153, ZN => n1131);
   U294 : INV_X1 port map( A => ADD_RDB(3), ZN => n2153);
   U295 : BUF_X1 port map( A => N298, Z => n214);
   U296 : BUF_X1 port map( A => N298, Z => n215);
   U297 : BUF_X1 port map( A => N299, Z => n211);
   U298 : BUF_X1 port map( A => N299, Z => n212);
   U299 : BUF_X1 port map( A => N300, Z => n208);
   U300 : BUF_X1 port map( A => N300, Z => n209);
   U301 : BUF_X1 port map( A => N301, Z => n205);
   U302 : BUF_X1 port map( A => N301, Z => n206);
   U303 : BUF_X1 port map( A => N302, Z => n202);
   U304 : BUF_X1 port map( A => N302, Z => n203);
   U305 : BUF_X1 port map( A => N303, Z => n199);
   U306 : BUF_X1 port map( A => N303, Z => n200);
   U307 : BUF_X1 port map( A => N304, Z => n196);
   U308 : BUF_X1 port map( A => N304, Z => n197);
   U309 : BUF_X1 port map( A => N305, Z => n193);
   U310 : BUF_X1 port map( A => N305, Z => n194);
   U311 : BUF_X1 port map( A => N243, Z => n379);
   U312 : BUF_X1 port map( A => N243, Z => n380);
   U313 : BUF_X1 port map( A => N276, Z => n280_port);
   U314 : BUF_X1 port map( A => N276, Z => n281_port);
   U315 : BUF_X1 port map( A => N277, Z => n277_port);
   U316 : BUF_X1 port map( A => N277, Z => n278_port);
   U317 : BUF_X1 port map( A => N278, Z => n274_port);
   U318 : BUF_X1 port map( A => N278, Z => n275_port);
   U319 : BUF_X1 port map( A => N279, Z => n271_port);
   U320 : BUF_X1 port map( A => N279, Z => n272_port);
   U321 : BUF_X1 port map( A => N280, Z => n268_port);
   U322 : BUF_X1 port map( A => N280, Z => n269_port);
   U323 : BUF_X1 port map( A => N281, Z => n265_port);
   U324 : BUF_X1 port map( A => N281, Z => n266_port);
   U325 : BUF_X1 port map( A => N282, Z => n262_port);
   U326 : BUF_X1 port map( A => N282, Z => n263_port);
   U327 : BUF_X1 port map( A => N283, Z => n259_port);
   U328 : BUF_X1 port map( A => N283, Z => n260_port);
   U329 : BUF_X1 port map( A => N284, Z => n256_port);
   U330 : BUF_X1 port map( A => N284, Z => n257_port);
   U331 : BUF_X1 port map( A => N285, Z => n253_port);
   U332 : BUF_X1 port map( A => N285, Z => n254_port);
   U333 : BUF_X1 port map( A => N286, Z => n250_port);
   U334 : BUF_X1 port map( A => N286, Z => n251_port);
   U335 : BUF_X1 port map( A => N287, Z => n247_port);
   U336 : BUF_X1 port map( A => N287, Z => n248_port);
   U337 : BUF_X1 port map( A => N288, Z => n244_port);
   U338 : BUF_X1 port map( A => N288, Z => n245_port);
   U339 : BUF_X1 port map( A => N289, Z => n241);
   U340 : BUF_X1 port map( A => N289, Z => n242);
   U341 : BUF_X1 port map( A => N290, Z => n238);
   U342 : BUF_X1 port map( A => N290, Z => n239);
   U343 : BUF_X1 port map( A => N291, Z => n235);
   U344 : BUF_X1 port map( A => N291, Z => n236);
   U345 : BUF_X1 port map( A => N292, Z => n232);
   U346 : BUF_X1 port map( A => N292, Z => n233);
   U347 : BUF_X1 port map( A => N293, Z => n229);
   U348 : BUF_X1 port map( A => N293, Z => n230);
   U349 : BUF_X1 port map( A => N294, Z => n226);
   U350 : BUF_X1 port map( A => N294, Z => n227);
   U351 : BUF_X1 port map( A => N295, Z => n223);
   U352 : BUF_X1 port map( A => N295, Z => n224);
   U353 : BUF_X1 port map( A => N296, Z => n220);
   U354 : BUF_X1 port map( A => N296, Z => n221);
   U355 : BUF_X1 port map( A => N297, Z => n217);
   U356 : BUF_X1 port map( A => N297, Z => n218);
   U357 : BUF_X1 port map( A => N298, Z => n216);
   U358 : BUF_X1 port map( A => N299, Z => n213);
   U359 : BUF_X1 port map( A => N300, Z => n210);
   U360 : BUF_X1 port map( A => N301, Z => n207);
   U361 : BUF_X1 port map( A => N302, Z => n204);
   U362 : BUF_X1 port map( A => N303, Z => n201);
   U363 : BUF_X1 port map( A => N304, Z => n198);
   U364 : BUF_X1 port map( A => N305, Z => n195);
   U365 : BUF_X1 port map( A => N243, Z => n381);
   U366 : BUF_X1 port map( A => N276, Z => n282_port);
   U367 : BUF_X1 port map( A => N277, Z => n279_port);
   U368 : BUF_X1 port map( A => N278, Z => n276_port);
   U369 : BUF_X1 port map( A => N279, Z => n273_port);
   U370 : BUF_X1 port map( A => N280, Z => n270_port);
   U371 : BUF_X1 port map( A => N281, Z => n267_port);
   U372 : BUF_X1 port map( A => N282, Z => n264_port);
   U373 : BUF_X1 port map( A => N283, Z => n261_port);
   U374 : BUF_X1 port map( A => N284, Z => n258_port);
   U375 : BUF_X1 port map( A => N285, Z => n255_port);
   U376 : BUF_X1 port map( A => N286, Z => n252_port);
   U377 : BUF_X1 port map( A => N287, Z => n249_port);
   U378 : BUF_X1 port map( A => N288, Z => n246_port);
   U379 : BUF_X1 port map( A => N289, Z => n243_port);
   U380 : BUF_X1 port map( A => N290, Z => n240);
   U381 : BUF_X1 port map( A => N291, Z => n237);
   U382 : BUF_X1 port map( A => N292, Z => n234);
   U383 : BUF_X1 port map( A => N293, Z => n231);
   U384 : BUF_X1 port map( A => N294, Z => n228);
   U385 : BUF_X1 port map( A => N295, Z => n225);
   U386 : BUF_X1 port map( A => N296, Z => n222);
   U387 : BUF_X1 port map( A => N297, Z => n219);
   U388 : BUF_X1 port map( A => n387, Z => n385);
   U389 : BUF_X1 port map( A => n387, Z => n384);
   U390 : BUF_X1 port map( A => n388, Z => n382);
   U391 : BUF_X1 port map( A => n388, Z => n383);
   U392 : BUF_X1 port map( A => n387, Z => n386);
   U393 : NOR2_X1 port map( A1 => ADD_RDA(1), A2 => ADD_RDA(2), ZN => n1751);
   U394 : NOR2_X1 port map( A1 => n2156, A2 => ADD_RDA(2), ZN => n1749);
   U395 : AND2_X1 port map( A1 => ADD_RDA(0), A2 => n1760, ZN => n1758);
   U396 : NOR2_X1 port map( A1 => ADD_RDA(3), A2 => ADD_RDA(4), ZN => n1769);
   U397 : AOI21_X1 port map( B1 => n1117, B2 => n1118, A => n391, ZN => N340);
   U398 : NOR4_X1 port map( A1 => n1137, A2 => n1138, A3 => n1139, A4 => n1140,
                           ZN => n1117);
   U399 : NOR4_X1 port map( A1 => n1119, A2 => n1120, A3 => n1121, A4 => n1122,
                           ZN => n1118);
   U400 : OAI21_X1 port map( B1 => n136, B2 => n443, A => n1141, ZN => n1140);
   U401 : AOI21_X1 port map( B1 => n1099, B2 => n1100, A => n391, ZN => N341);
   U402 : NOR4_X1 port map( A1 => n1109, A2 => n1110, A3 => n1111, A4 => n1112,
                           ZN => n1099);
   U403 : NOR4_X1 port map( A1 => n1101, A2 => n1102, A3 => n1103, A4 => n1104,
                           ZN => n1100);
   U404 : OAI21_X1 port map( B1 => n136, B2 => n442, A => n1113, ZN => n1112);
   U405 : AOI21_X1 port map( B1 => n1081, B2 => n1082, A => n391, ZN => N342);
   U406 : NOR4_X1 port map( A1 => n1091, A2 => n1092, A3 => n1093, A4 => n1094,
                           ZN => n1081);
   U407 : NOR4_X1 port map( A1 => n1083, A2 => n1084, A3 => n1085, A4 => n1086,
                           ZN => n1082);
   U408 : OAI21_X1 port map( B1 => n136, B2 => n441, A => n1095, ZN => n1094);
   U409 : AOI21_X1 port map( B1 => n1063, B2 => n1064, A => n391, ZN => N343);
   U410 : NOR4_X1 port map( A1 => n1073, A2 => n1074, A3 => n1075, A4 => n1076,
                           ZN => n1063);
   U411 : NOR4_X1 port map( A1 => n1065, A2 => n1066, A3 => n1067, A4 => n1068,
                           ZN => n1064);
   U412 : OAI21_X1 port map( B1 => n136, B2 => n440, A => n1077, ZN => n1076);
   U413 : AOI21_X1 port map( B1 => n1045, B2 => n1046, A => n391, ZN => N344);
   U414 : NOR4_X1 port map( A1 => n1055, A2 => n1056, A3 => n1057, A4 => n1058,
                           ZN => n1045);
   U415 : NOR4_X1 port map( A1 => n1047, A2 => n1048, A3 => n1049, A4 => n1050,
                           ZN => n1046);
   U416 : OAI21_X1 port map( B1 => n136, B2 => n439, A => n1059, ZN => n1058);
   U417 : AOI21_X1 port map( B1 => n1027, B2 => n1028, A => n391, ZN => N345);
   U418 : NOR4_X1 port map( A1 => n1037, A2 => n1038, A3 => n1039, A4 => n1040,
                           ZN => n1027);
   U419 : NOR4_X1 port map( A1 => n1029, A2 => n1030, A3 => n1031, A4 => n1032,
                           ZN => n1028);
   U420 : OAI21_X1 port map( B1 => n136, B2 => n438, A => n1041, ZN => n1040);
   U421 : AOI21_X1 port map( B1 => n1009, B2 => n1010, A => n391, ZN => N346);
   U422 : NOR4_X1 port map( A1 => n1019, A2 => n1020, A3 => n1021, A4 => n1022,
                           ZN => n1009);
   U423 : NOR4_X1 port map( A1 => n1011, A2 => n1012, A3 => n1013, A4 => n1014,
                           ZN => n1010);
   U424 : OAI21_X1 port map( B1 => n136, B2 => n437, A => n1023, ZN => n1022);
   U425 : AOI21_X1 port map( B1 => n991, B2 => n992, A => n391, ZN => N347);
   U426 : NOR4_X1 port map( A1 => n1001, A2 => n1002, A3 => n1003, A4 => n1004,
                           ZN => n991);
   U427 : NOR4_X1 port map( A1 => n993, A2 => n994, A3 => n995, A4 => n996, ZN 
                           => n992);
   U428 : OAI21_X1 port map( B1 => n136, B2 => n436, A => n1005, ZN => n1004);
   U429 : AOI21_X1 port map( B1 => n973, B2 => n974, A => n390, ZN => N348);
   U430 : NOR4_X1 port map( A1 => n983, A2 => n984, A3 => n985, A4 => n986, ZN 
                           => n973);
   U431 : NOR4_X1 port map( A1 => n975, A2 => n976, A3 => n977, A4 => n978, ZN 
                           => n974);
   U432 : OAI21_X1 port map( B1 => n136, B2 => n435, A => n987, ZN => n986);
   U433 : AOI21_X1 port map( B1 => n955, B2 => n956, A => n390, ZN => N349);
   U434 : NOR4_X1 port map( A1 => n965, A2 => n966, A3 => n967, A4 => n968, ZN 
                           => n955);
   U435 : NOR4_X1 port map( A1 => n957, A2 => n958, A3 => n959, A4 => n960, ZN 
                           => n956);
   U436 : OAI21_X1 port map( B1 => n136, B2 => n434, A => n969, ZN => n968);
   U437 : AOI21_X1 port map( B1 => n937, B2 => n938, A => n390, ZN => N350);
   U438 : NOR4_X1 port map( A1 => n947, A2 => n948, A3 => n949, A4 => n950, ZN 
                           => n937);
   U439 : NOR4_X1 port map( A1 => n939, A2 => n940, A3 => n941, A4 => n942, ZN 
                           => n938);
   U440 : OAI21_X1 port map( B1 => n136, B2 => n433, A => n951, ZN => n950);
   U441 : AOI21_X1 port map( B1 => n919, B2 => n920, A => n390, ZN => N351);
   U442 : NOR4_X1 port map( A1 => n929, A2 => n930, A3 => n931, A4 => n932, ZN 
                           => n919);
   U443 : NOR4_X1 port map( A1 => n921, A2 => n922, A3 => n923, A4 => n924, ZN 
                           => n920);
   U444 : OAI21_X1 port map( B1 => n136, B2 => n432, A => n933, ZN => n932);
   U445 : AOI21_X1 port map( B1 => n901, B2 => n902, A => n390, ZN => N352);
   U446 : NOR4_X1 port map( A1 => n911, A2 => n912, A3 => n913, A4 => n914, ZN 
                           => n901);
   U447 : NOR4_X1 port map( A1 => n903, A2 => n904, A3 => n905, A4 => n906, ZN 
                           => n902);
   U448 : OAI21_X1 port map( B1 => n137, B2 => n431, A => n915, ZN => n914);
   U449 : AOI21_X1 port map( B1 => n883, B2 => n884, A => n390, ZN => N353);
   U450 : NOR4_X1 port map( A1 => n893, A2 => n894, A3 => n895, A4 => n896, ZN 
                           => n883);
   U451 : NOR4_X1 port map( A1 => n885, A2 => n886, A3 => n887, A4 => n888, ZN 
                           => n884);
   U452 : OAI21_X1 port map( B1 => n137, B2 => n430, A => n897, ZN => n896);
   U453 : AOI21_X1 port map( B1 => n865, B2 => n866, A => n390, ZN => N354);
   U454 : NOR4_X1 port map( A1 => n875, A2 => n876, A3 => n877, A4 => n878, ZN 
                           => n865);
   U455 : NOR4_X1 port map( A1 => n867, A2 => n868, A3 => n869, A4 => n870, ZN 
                           => n866);
   U456 : OAI21_X1 port map( B1 => n137, B2 => n429, A => n879, ZN => n878);
   U457 : AOI21_X1 port map( B1 => n847, B2 => n848, A => n390, ZN => N355);
   U458 : NOR4_X1 port map( A1 => n857, A2 => n858, A3 => n859, A4 => n860, ZN 
                           => n847);
   U459 : NOR4_X1 port map( A1 => n849, A2 => n850, A3 => n851, A4 => n852, ZN 
                           => n848);
   U460 : OAI21_X1 port map( B1 => n137, B2 => n428, A => n861, ZN => n860);
   U461 : AOI21_X1 port map( B1 => n829, B2 => n830, A => n390, ZN => N356);
   U462 : NOR4_X1 port map( A1 => n839, A2 => n840, A3 => n841, A4 => n842, ZN 
                           => n829);
   U463 : NOR4_X1 port map( A1 => n831, A2 => n832, A3 => n833, A4 => n834, ZN 
                           => n830);
   U464 : OAI21_X1 port map( B1 => n137, B2 => n427, A => n843, ZN => n842);
   U465 : AOI21_X1 port map( B1 => n811, B2 => n812, A => n390, ZN => N357);
   U466 : NOR4_X1 port map( A1 => n821, A2 => n822, A3 => n823, A4 => n824, ZN 
                           => n811);
   U467 : NOR4_X1 port map( A1 => n813, A2 => n814, A3 => n815, A4 => n816, ZN 
                           => n812);
   U468 : OAI21_X1 port map( B1 => n137, B2 => n426, A => n825, ZN => n824);
   U469 : AOI21_X1 port map( B1 => n793, B2 => n794, A => n390, ZN => N358);
   U470 : NOR4_X1 port map( A1 => n803, A2 => n804, A3 => n805, A4 => n806, ZN 
                           => n793);
   U471 : NOR4_X1 port map( A1 => n795, A2 => n796, A3 => n797, A4 => n798, ZN 
                           => n794);
   U472 : OAI21_X1 port map( B1 => n137, B2 => n425, A => n807, ZN => n806);
   U473 : AOI21_X1 port map( B1 => n775, B2 => n776, A => n390, ZN => N359);
   U474 : NOR4_X1 port map( A1 => n785, A2 => n786, A3 => n787, A4 => n788, ZN 
                           => n775);
   U475 : NOR4_X1 port map( A1 => n777, A2 => n778, A3 => n779, A4 => n780, ZN 
                           => n776);
   U476 : OAI21_X1 port map( B1 => n137, B2 => n424, A => n789, ZN => n788);
   U477 : AOI21_X1 port map( B1 => n757, B2 => n758, A => n389, ZN => N360);
   U478 : NOR4_X1 port map( A1 => n767, A2 => n768, A3 => n769, A4 => n770, ZN 
                           => n757);
   U479 : NOR4_X1 port map( A1 => n759, A2 => n760, A3 => n761, A4 => n762, ZN 
                           => n758);
   U480 : OAI21_X1 port map( B1 => n137, B2 => n423, A => n771, ZN => n770);
   U481 : AOI21_X1 port map( B1 => n739, B2 => n740, A => n389, ZN => N361);
   U482 : NOR4_X1 port map( A1 => n749, A2 => n750, A3 => n751, A4 => n752, ZN 
                           => n739);
   U483 : NOR4_X1 port map( A1 => n741, A2 => n742, A3 => n743, A4 => n744, ZN 
                           => n740);
   U484 : OAI21_X1 port map( B1 => n137, B2 => n422, A => n753, ZN => n752);
   U485 : AOI21_X1 port map( B1 => n721, B2 => n722, A => n389, ZN => N362);
   U486 : NOR4_X1 port map( A1 => n731, A2 => n732, A3 => n733, A4 => n734, ZN 
                           => n721);
   U487 : NOR4_X1 port map( A1 => n723, A2 => n724, A3 => n725, A4 => n726, ZN 
                           => n722);
   U488 : OAI21_X1 port map( B1 => n137, B2 => n421, A => n735, ZN => n734);
   U489 : AOI21_X1 port map( B1 => n703, B2 => n704, A => n389, ZN => N363);
   U490 : NOR4_X1 port map( A1 => n713, A2 => n714, A3 => n715, A4 => n716, ZN 
                           => n703);
   U491 : NOR4_X1 port map( A1 => n705, A2 => n706, A3 => n707, A4 => n708, ZN 
                           => n704);
   U492 : OAI21_X1 port map( B1 => n137, B2 => n420, A => n717, ZN => n716);
   U493 : AOI21_X1 port map( B1 => n685, B2 => n686, A => n389, ZN => N364);
   U494 : NOR4_X1 port map( A1 => n695, A2 => n696, A3 => n697, A4 => n698, ZN 
                           => n685);
   U495 : NOR4_X1 port map( A1 => n687, A2 => n688, A3 => n689, A4 => n690, ZN 
                           => n686);
   U496 : OAI21_X1 port map( B1 => n138, B2 => n419, A => n699, ZN => n698);
   U497 : AOI21_X1 port map( B1 => n667, B2 => n668, A => n389, ZN => N365);
   U498 : NOR4_X1 port map( A1 => n677, A2 => n678, A3 => n679, A4 => n680, ZN 
                           => n667);
   U499 : NOR4_X1 port map( A1 => n669, A2 => n670, A3 => n671, A4 => n672, ZN 
                           => n668);
   U500 : OAI21_X1 port map( B1 => n138, B2 => n418, A => n681, ZN => n680);
   U501 : AOI21_X1 port map( B1 => n649, B2 => n650, A => n389, ZN => N366);
   U502 : NOR4_X1 port map( A1 => n659, A2 => n660, A3 => n661, A4 => n662, ZN 
                           => n649);
   U503 : NOR4_X1 port map( A1 => n651, A2 => n652, A3 => n653, A4 => n654, ZN 
                           => n650);
   U504 : OAI21_X1 port map( B1 => n138, B2 => n417, A => n663, ZN => n662);
   U505 : AOI21_X1 port map( B1 => n631, B2 => n632, A => n389, ZN => N367);
   U506 : NOR4_X1 port map( A1 => n641, A2 => n642, A3 => n643, A4 => n644, ZN 
                           => n631);
   U507 : NOR4_X1 port map( A1 => n633, A2 => n634, A3 => n635, A4 => n636, ZN 
                           => n632);
   U508 : OAI21_X1 port map( B1 => n138, B2 => n416, A => n645, ZN => n644);
   U509 : AOI21_X1 port map( B1 => n613, B2 => n614, A => n389, ZN => N368);
   U510 : NOR4_X1 port map( A1 => n623, A2 => n624, A3 => n625, A4 => n626, ZN 
                           => n613);
   U511 : NOR4_X1 port map( A1 => n615, A2 => n616, A3 => n617, A4 => n618, ZN 
                           => n614);
   U512 : OAI21_X1 port map( B1 => n138, B2 => n415, A => n627, ZN => n626);
   U513 : AOI21_X1 port map( B1 => n595, B2 => n596, A => n389, ZN => N369);
   U514 : NOR4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, ZN 
                           => n595);
   U515 : NOR4_X1 port map( A1 => n597, A2 => n598, A3 => n599, A4 => n600, ZN 
                           => n596);
   U516 : OAI21_X1 port map( B1 => n138, B2 => n414, A => n609, ZN => n608);
   U517 : AOI21_X1 port map( B1 => n577, B2 => n578, A => n389, ZN => N370);
   U518 : NOR4_X1 port map( A1 => n587, A2 => n588, A3 => n589, A4 => n590, ZN 
                           => n577);
   U519 : NOR4_X1 port map( A1 => n579, A2 => n580, A3 => n581, A4 => n582, ZN 
                           => n578);
   U520 : OAI21_X1 port map( B1 => n138, B2 => n413, A => n591, ZN => n590);
   U521 : AOI21_X1 port map( B1 => n527, B2 => n528, A => n389, ZN => N371);
   U522 : NOR4_X1 port map( A1 => n553, A2 => n554, A3 => n555, A4 => n556, ZN 
                           => n527);
   U523 : NOR4_X1 port map( A1 => n529, A2 => n530, A3 => n531, A4 => n532, ZN 
                           => n528);
   U524 : OAI21_X1 port map( B1 => n138, B2 => n412, A => n559, ZN => n556);
   U525 : AOI21_X1 port map( B1 => n1669, B2 => n1670, A => n393, ZN => N312);
   U526 : NOR4_X1 port map( A1 => n1679, A2 => n1680, A3 => n1681, A4 => n1682,
                           ZN => n1669);
   U527 : NOR4_X1 port map( A1 => n1671, A2 => n1672, A3 => n1673, A4 => n1674,
                           ZN => n1670);
   U528 : OAI221_X1 port map( B1 => n1889, B2 => n10, C1 => n1857, C2 => n7, A 
                           => n1686, ZN => n1679);
   U529 : AOI21_X1 port map( B1 => n1651, B2 => n1652, A => n393, ZN => N313);
   U530 : NOR4_X1 port map( A1 => n1661, A2 => n1662, A3 => n1663, A4 => n1664,
                           ZN => n1651);
   U531 : NOR4_X1 port map( A1 => n1653, A2 => n1654, A3 => n1655, A4 => n1656,
                           ZN => n1652);
   U532 : OAI221_X1 port map( B1 => n1888, B2 => n10, C1 => n1856, C2 => n7, A 
                           => n1668, ZN => n1661);
   U533 : AOI21_X1 port map( B1 => n1633, B2 => n1634, A => n393, ZN => N314);
   U534 : NOR4_X1 port map( A1 => n1643, A2 => n1644, A3 => n1645, A4 => n1646,
                           ZN => n1633);
   U535 : NOR4_X1 port map( A1 => n1635, A2 => n1636, A3 => n1637, A4 => n1638,
                           ZN => n1634);
   U536 : OAI221_X1 port map( B1 => n1887, B2 => n10, C1 => n1855, C2 => n7, A 
                           => n1650, ZN => n1643);
   U537 : AOI21_X1 port map( B1 => n1615, B2 => n1616, A => n393, ZN => N315);
   U538 : NOR4_X1 port map( A1 => n1625, A2 => n1626, A3 => n1627, A4 => n1628,
                           ZN => n1615);
   U539 : NOR4_X1 port map( A1 => n1617, A2 => n1618, A3 => n1619, A4 => n1620,
                           ZN => n1616);
   U540 : OAI221_X1 port map( B1 => n1886, B2 => n10, C1 => n1854, C2 => n7, A 
                           => n1632, ZN => n1625);
   U541 : AOI21_X1 port map( B1 => n1597, B2 => n1598, A => n393, ZN => N316);
   U542 : NOR4_X1 port map( A1 => n1607, A2 => n1608, A3 => n1609, A4 => n1610,
                           ZN => n1597);
   U543 : NOR4_X1 port map( A1 => n1599, A2 => n1600, A3 => n1601, A4 => n1602,
                           ZN => n1598);
   U544 : OAI221_X1 port map( B1 => n1885, B2 => n10, C1 => n1853, C2 => n7, A 
                           => n1614, ZN => n1607);
   U545 : AOI21_X1 port map( B1 => n1579, B2 => n1580, A => n393, ZN => N317);
   U546 : NOR4_X1 port map( A1 => n1589, A2 => n1590, A3 => n1591, A4 => n1592,
                           ZN => n1579);
   U547 : NOR4_X1 port map( A1 => n1581, A2 => n1582, A3 => n1583, A4 => n1584,
                           ZN => n1580);
   U548 : OAI221_X1 port map( B1 => n1884, B2 => n10, C1 => n1852, C2 => n7, A 
                           => n1596, ZN => n1589);
   U549 : AOI21_X1 port map( B1 => n1561, B2 => n1562, A => n393, ZN => N318);
   U550 : NOR4_X1 port map( A1 => n1571, A2 => n1572, A3 => n1573, A4 => n1574,
                           ZN => n1561);
   U551 : NOR4_X1 port map( A1 => n1563, A2 => n1564, A3 => n1565, A4 => n1566,
                           ZN => n1562);
   U552 : OAI221_X1 port map( B1 => n1883, B2 => n10, C1 => n1851, C2 => n7, A 
                           => n1578, ZN => n1571);
   U553 : AOI21_X1 port map( B1 => n1543, B2 => n1544, A => n393, ZN => N319);
   U554 : NOR4_X1 port map( A1 => n1553, A2 => n1554, A3 => n1555, A4 => n1556,
                           ZN => n1543);
   U555 : NOR4_X1 port map( A1 => n1545, A2 => n1546, A3 => n1547, A4 => n1548,
                           ZN => n1544);
   U556 : OAI221_X1 port map( B1 => n1882, B2 => n10, C1 => n1850, C2 => n7, A 
                           => n1560, ZN => n1553);
   U557 : AOI21_X1 port map( B1 => n1525, B2 => n1526, A => n393, ZN => N320);
   U558 : NOR4_X1 port map( A1 => n1535, A2 => n1536, A3 => n1537, A4 => n1538,
                           ZN => n1525);
   U559 : NOR4_X1 port map( A1 => n1527, A2 => n1528, A3 => n1529, A4 => n1530,
                           ZN => n1526);
   U560 : OAI221_X1 port map( B1 => n1881, B2 => n11, C1 => n1849, C2 => n8, A 
                           => n1542, ZN => n1535);
   U561 : AOI21_X1 port map( B1 => n1507, B2 => n1508, A => n393, ZN => N321);
   U562 : NOR4_X1 port map( A1 => n1517, A2 => n1518, A3 => n1519, A4 => n1520,
                           ZN => n1507);
   U563 : NOR4_X1 port map( A1 => n1509, A2 => n1510, A3 => n1511, A4 => n1512,
                           ZN => n1508);
   U564 : OAI221_X1 port map( B1 => n1880, B2 => n11, C1 => n1848, C2 => n8, A 
                           => n1524, ZN => n1517);
   U565 : AOI21_X1 port map( B1 => n1489, B2 => n1490, A => n393, ZN => N322);
   U566 : NOR4_X1 port map( A1 => n1499, A2 => n1500, A3 => n1501, A4 => n1502,
                           ZN => n1489);
   U567 : NOR4_X1 port map( A1 => n1491, A2 => n1492, A3 => n1493, A4 => n1494,
                           ZN => n1490);
   U568 : OAI221_X1 port map( B1 => n1879, B2 => n11, C1 => n1847, C2 => n8, A 
                           => n1506, ZN => n1499);
   U569 : AOI21_X1 port map( B1 => n1471, B2 => n1472, A => n393, ZN => N323);
   U570 : NOR4_X1 port map( A1 => n1481, A2 => n1482, A3 => n1483, A4 => n1484,
                           ZN => n1471);
   U571 : NOR4_X1 port map( A1 => n1473, A2 => n1474, A3 => n1475, A4 => n1476,
                           ZN => n1472);
   U572 : OAI221_X1 port map( B1 => n1878, B2 => n11, C1 => n1846, C2 => n8, A 
                           => n1488, ZN => n1481);
   U573 : AOI21_X1 port map( B1 => n1453, B2 => n1454, A => n392, ZN => N324);
   U574 : NOR4_X1 port map( A1 => n1463, A2 => n1464, A3 => n1465, A4 => n1466,
                           ZN => n1453);
   U575 : NOR4_X1 port map( A1 => n1455, A2 => n1456, A3 => n1457, A4 => n1458,
                           ZN => n1454);
   U576 : OAI221_X1 port map( B1 => n1877, B2 => n11, C1 => n1845, C2 => n8, A 
                           => n1470, ZN => n1463);
   U577 : AOI21_X1 port map( B1 => n1435, B2 => n1436, A => n392, ZN => N325);
   U578 : NOR4_X1 port map( A1 => n1445, A2 => n1446, A3 => n1447, A4 => n1448,
                           ZN => n1435);
   U579 : NOR4_X1 port map( A1 => n1437, A2 => n1438, A3 => n1439, A4 => n1440,
                           ZN => n1436);
   U580 : OAI221_X1 port map( B1 => n1876, B2 => n11, C1 => n1844, C2 => n8, A 
                           => n1452, ZN => n1445);
   U581 : AOI21_X1 port map( B1 => n1417, B2 => n1418, A => n392, ZN => N326);
   U582 : NOR4_X1 port map( A1 => n1427, A2 => n1428, A3 => n1429, A4 => n1430,
                           ZN => n1417);
   U583 : NOR4_X1 port map( A1 => n1419, A2 => n1420, A3 => n1421, A4 => n1422,
                           ZN => n1418);
   U584 : OAI221_X1 port map( B1 => n1875, B2 => n11, C1 => n1843, C2 => n8, A 
                           => n1434, ZN => n1427);
   U585 : AOI21_X1 port map( B1 => n1399, B2 => n1400, A => n392, ZN => N327);
   U586 : NOR4_X1 port map( A1 => n1409, A2 => n1410, A3 => n1411, A4 => n1412,
                           ZN => n1399);
   U587 : NOR4_X1 port map( A1 => n1401, A2 => n1402, A3 => n1403, A4 => n1404,
                           ZN => n1400);
   U588 : OAI221_X1 port map( B1 => n1874, B2 => n11, C1 => n1842, C2 => n8, A 
                           => n1416, ZN => n1409);
   U589 : AOI21_X1 port map( B1 => n1381, B2 => n1382, A => n392, ZN => N328);
   U590 : NOR4_X1 port map( A1 => n1391, A2 => n1392, A3 => n1393, A4 => n1394,
                           ZN => n1381);
   U591 : NOR4_X1 port map( A1 => n1383, A2 => n1384, A3 => n1385, A4 => n1386,
                           ZN => n1382);
   U592 : OAI221_X1 port map( B1 => n1873, B2 => n11, C1 => n1841, C2 => n8, A 
                           => n1398, ZN => n1391);
   U593 : AOI21_X1 port map( B1 => n1363, B2 => n1364, A => n392, ZN => N329);
   U594 : NOR4_X1 port map( A1 => n1373, A2 => n1374, A3 => n1375, A4 => n1376,
                           ZN => n1363);
   U595 : NOR4_X1 port map( A1 => n1365, A2 => n1366, A3 => n1367, A4 => n1368,
                           ZN => n1364);
   U596 : OAI221_X1 port map( B1 => n1872, B2 => n11, C1 => n1840, C2 => n8, A 
                           => n1380, ZN => n1373);
   U597 : AOI21_X1 port map( B1 => n1345, B2 => n1346, A => n392, ZN => N330);
   U598 : NOR4_X1 port map( A1 => n1355, A2 => n1356, A3 => n1357, A4 => n1358,
                           ZN => n1345);
   U599 : NOR4_X1 port map( A1 => n1347, A2 => n1348, A3 => n1349, A4 => n1350,
                           ZN => n1346);
   U600 : OAI221_X1 port map( B1 => n1871, B2 => n11, C1 => n1839, C2 => n8, A 
                           => n1362, ZN => n1355);
   U601 : AOI21_X1 port map( B1 => n1327, B2 => n1328, A => n392, ZN => N331);
   U602 : NOR4_X1 port map( A1 => n1337, A2 => n1338, A3 => n1339, A4 => n1340,
                           ZN => n1327);
   U603 : NOR4_X1 port map( A1 => n1329, A2 => n1330, A3 => n1331, A4 => n1332,
                           ZN => n1328);
   U604 : OAI221_X1 port map( B1 => n1870, B2 => n11, C1 => n1838, C2 => n8, A 
                           => n1344, ZN => n1337);
   U605 : AOI21_X1 port map( B1 => n1309, B2 => n1310, A => n392, ZN => N332);
   U606 : NOR4_X1 port map( A1 => n1319, A2 => n1320, A3 => n1321, A4 => n1322,
                           ZN => n1309);
   U607 : NOR4_X1 port map( A1 => n1311, A2 => n1312, A3 => n1313, A4 => n1314,
                           ZN => n1310);
   U608 : OAI221_X1 port map( B1 => n1869, B2 => n12, C1 => n1837, C2 => n9, A 
                           => n1326, ZN => n1319);
   U609 : AOI21_X1 port map( B1 => n1291, B2 => n1292, A => n392, ZN => N333);
   U610 : NOR4_X1 port map( A1 => n1301, A2 => n1302, A3 => n1303, A4 => n1304,
                           ZN => n1291);
   U611 : NOR4_X1 port map( A1 => n1293, A2 => n1294, A3 => n1295, A4 => n1296,
                           ZN => n1292);
   U612 : OAI221_X1 port map( B1 => n1868, B2 => n12, C1 => n1836, C2 => n9, A 
                           => n1308, ZN => n1301);
   U613 : AOI21_X1 port map( B1 => n1273, B2 => n1274, A => n392, ZN => N334);
   U614 : NOR4_X1 port map( A1 => n1283, A2 => n1284, A3 => n1285, A4 => n1286,
                           ZN => n1273);
   U615 : NOR4_X1 port map( A1 => n1275, A2 => n1276, A3 => n1277, A4 => n1278,
                           ZN => n1274);
   U616 : OAI221_X1 port map( B1 => n1867, B2 => n12, C1 => n1835, C2 => n9, A 
                           => n1290, ZN => n1283);
   U617 : AOI21_X1 port map( B1 => n1255, B2 => n1256, A => n392, ZN => N335);
   U618 : NOR4_X1 port map( A1 => n1265, A2 => n1266, A3 => n1267, A4 => n1268,
                           ZN => n1255);
   U619 : NOR4_X1 port map( A1 => n1257, A2 => n1258, A3 => n1259, A4 => n1260,
                           ZN => n1256);
   U620 : OAI221_X1 port map( B1 => n1866, B2 => n12, C1 => n1834, C2 => n9, A 
                           => n1272, ZN => n1265);
   U621 : AOI21_X1 port map( B1 => n1237, B2 => n1238, A => n391, ZN => N336);
   U622 : NOR4_X1 port map( A1 => n1247, A2 => n1248, A3 => n1249, A4 => n1250,
                           ZN => n1237);
   U623 : NOR4_X1 port map( A1 => n1239, A2 => n1240, A3 => n1241, A4 => n1242,
                           ZN => n1238);
   U624 : OAI221_X1 port map( B1 => n1865, B2 => n12, C1 => n1833, C2 => n9, A 
                           => n1254, ZN => n1247);
   U625 : AOI21_X1 port map( B1 => n1219, B2 => n1220, A => n391, ZN => N337);
   U626 : NOR4_X1 port map( A1 => n1229, A2 => n1230, A3 => n1231, A4 => n1232,
                           ZN => n1219);
   U627 : NOR4_X1 port map( A1 => n1221, A2 => n1222, A3 => n1223, A4 => n1224,
                           ZN => n1220);
   U628 : OAI221_X1 port map( B1 => n1864, B2 => n12, C1 => n1832, C2 => n9, A 
                           => n1236, ZN => n1229);
   U629 : AOI21_X1 port map( B1 => n1201, B2 => n1202, A => n391, ZN => N338);
   U630 : NOR4_X1 port map( A1 => n1211, A2 => n1212, A3 => n1213, A4 => n1214,
                           ZN => n1201);
   U631 : NOR4_X1 port map( A1 => n1203, A2 => n1204, A3 => n1205, A4 => n1206,
                           ZN => n1202);
   U632 : OAI221_X1 port map( B1 => n1863, B2 => n12, C1 => n1831, C2 => n9, A 
                           => n1218, ZN => n1211);
   U633 : AOI21_X1 port map( B1 => n1151, B2 => n1152, A => n391, ZN => N339);
   U634 : NOR4_X1 port map( A1 => n1177, A2 => n1178, A3 => n1179, A4 => n1180,
                           ZN => n1151);
   U635 : NOR4_X1 port map( A1 => n1153, A2 => n1154, A3 => n1155, A4 => n1156,
                           ZN => n1152);
   U636 : OAI221_X1 port map( B1 => n1862, B2 => n12, C1 => n1830, C2 => n9, A 
                           => n1198, ZN => n1177);
   U637 : NOR2_X1 port map( A1 => n2154, A2 => ADD_RDA(4), ZN => n1774);
   U638 : AND2_X1 port map( A1 => n1755, A2 => ADD_RDA(0), ZN => n1750);
   U639 : AND2_X1 port map( A1 => n1774, A2 => ADD_RDA(0), ZN => n1772);
   U640 : AND2_X1 port map( A1 => n1769, A2 => ADD_RDA(0), ZN => n1767);
   U641 : AOI21_X1 port map( B1 => n1741, B2 => n1742, A => n390, ZN => N308);
   U642 : NOR4_X1 port map( A1 => n1761, A2 => n1762, A3 => n1763, A4 => n1764,
                           ZN => n1741);
   U643 : NOR4_X1 port map( A1 => n1743, A2 => n1744, A3 => n1745, A4 => n1746,
                           ZN => n1742);
   U644 : OAI221_X1 port map( B1 => n1893, B2 => n10, C1 => n1861, C2 => n7, A 
                           => n1773, ZN => n1761);
   U645 : AOI21_X1 port map( B1 => n1723, B2 => n1724, A => n389, ZN => N309);
   U646 : NOR4_X1 port map( A1 => n1733, A2 => n1734, A3 => n1735, A4 => n1736,
                           ZN => n1723);
   U647 : NOR4_X1 port map( A1 => n1725, A2 => n1726, A3 => n1727, A4 => n1728,
                           ZN => n1724);
   U648 : OAI221_X1 port map( B1 => n1892, B2 => n10, C1 => n1860, C2 => n7, A 
                           => n1740, ZN => n1733);
   U649 : AOI21_X1 port map( B1 => n1705, B2 => n1706, A => n393, ZN => N310);
   U650 : NOR4_X1 port map( A1 => n1715, A2 => n1716, A3 => n1717, A4 => n1718,
                           ZN => n1705);
   U651 : NOR4_X1 port map( A1 => n1707, A2 => n1708, A3 => n1709, A4 => n1710,
                           ZN => n1706);
   U652 : OAI221_X1 port map( B1 => n1891, B2 => n10, C1 => n1859, C2 => n7, A 
                           => n1722, ZN => n1715);
   U653 : AOI21_X1 port map( B1 => n1687, B2 => n1688, A => n392, ZN => N311);
   U654 : NOR4_X1 port map( A1 => n1697, A2 => n1698, A3 => n1699, A4 => n1700,
                           ZN => n1687);
   U655 : NOR4_X1 port map( A1 => n1689, A2 => n1690, A3 => n1691, A4 => n1692,
                           ZN => n1688);
   U656 : OAI221_X1 port map( B1 => n1890, B2 => n10, C1 => n1858, C2 => n7, A 
                           => n1704, ZN => n1697);
   U657 : INV_X1 port map( A => ADD_RDA(0), ZN => n2157);
   U658 : INV_X1 port map( A => ADD_RDA(1), ZN => n2156);
   U659 : INV_X1 port map( A => ADD_RDA(2), ZN => n2155);
   U660 : INV_X1 port map( A => ADD_RDA(3), ZN => n2154);
   U661 : AND2_X1 port map( A1 => ADD_RDA(4), A2 => ADD_RDA(3), ZN => n1760);
   U662 : AND2_X1 port map( A1 => ADD_RDA(4), A2 => n2154, ZN => n1755);
   U663 : OAI21_X1 port map( B1 => n1783, B2 => n1784, A => n395, ZN => N298);
   U664 : OAI21_X1 port map( B1 => n1775, B2 => n1782, A => n395, ZN => N299);
   U665 : OAI21_X1 port map( B1 => n1775, B2 => n1781, A => n395, ZN => N300);
   U666 : OAI21_X1 port map( B1 => n1775, B2 => n1780, A => n394, ZN => N301);
   U667 : OAI21_X1 port map( B1 => n1775, B2 => n1779, A => n394, ZN => N302);
   U668 : OAI21_X1 port map( B1 => n1775, B2 => n1778, A => n394, ZN => N303);
   U669 : OAI21_X1 port map( B1 => n1775, B2 => n1777, A => n394, ZN => N304);
   U670 : OAI21_X1 port map( B1 => n1775, B2 => n1776, A => n398, ZN => N305);
   U671 : OAI21_X1 port map( B1 => n1782, B2 => n1786, A => n395, ZN => N243);
   U672 : OAI21_X1 port map( B1 => n1781, B2 => n1786, A => n401, ZN => N276);
   U673 : OAI21_X1 port map( B1 => n1780, B2 => n1786, A => n401, ZN => N277);
   U674 : OAI21_X1 port map( B1 => n1779, B2 => n1786, A => n401, ZN => N278);
   U675 : OAI21_X1 port map( B1 => n1778, B2 => n1786, A => n400, ZN => N279);
   U676 : OAI21_X1 port map( B1 => n1777, B2 => n1786, A => n400, ZN => N280);
   U677 : OAI21_X1 port map( B1 => n1776, B2 => n1786, A => n400, ZN => N281);
   U678 : OAI21_X1 port map( B1 => n1784, B2 => n1786, A => n400, ZN => N282);
   U679 : OAI21_X1 port map( B1 => n1782, B2 => n1785, A => n399, ZN => N283);
   U680 : OAI21_X1 port map( B1 => n1781, B2 => n1785, A => n399, ZN => N284);
   U681 : OAI21_X1 port map( B1 => n1780, B2 => n1785, A => n399, ZN => N285);
   U682 : OAI21_X1 port map( B1 => n1779, B2 => n1785, A => n399, ZN => N286);
   U683 : OAI21_X1 port map( B1 => n1778, B2 => n1785, A => n398, ZN => N287);
   U684 : OAI21_X1 port map( B1 => n1777, B2 => n1785, A => n398, ZN => N288);
   U685 : OAI21_X1 port map( B1 => n1776, B2 => n1785, A => n398, ZN => N289);
   U686 : OAI21_X1 port map( B1 => n1784, B2 => n1785, A => n397, ZN => N290);
   U687 : OAI21_X1 port map( B1 => n1782, B2 => n1783, A => n397, ZN => N291);
   U688 : OAI21_X1 port map( B1 => n1781, B2 => n1783, A => n397, ZN => N292);
   U689 : OAI21_X1 port map( B1 => n1780, B2 => n1783, A => n397, ZN => N293);
   U690 : OAI21_X1 port map( B1 => n1779, B2 => n1783, A => n396, ZN => N294);
   U691 : OAI21_X1 port map( B1 => n1778, B2 => n1783, A => n396, ZN => N295);
   U692 : OAI21_X1 port map( B1 => n1777, B2 => n1783, A => n396, ZN => N296);
   U693 : OAI21_X1 port map( B1 => n1776, B2 => n1783, A => n396, ZN => N297);
   U694 : BUF_X1 port map( A => N244, Z => n377);
   U695 : BUF_X1 port map( A => N245, Z => n374);
   U696 : BUF_X1 port map( A => N246, Z => n371_port);
   U697 : BUF_X1 port map( A => N247, Z => n368_port);
   U698 : BUF_X1 port map( A => N248, Z => n365_port);
   U699 : BUF_X1 port map( A => N249, Z => n362_port);
   U700 : BUF_X1 port map( A => N250, Z => n359_port);
   U701 : BUF_X1 port map( A => N251, Z => n356_port);
   U702 : BUF_X1 port map( A => N252, Z => n353_port);
   U703 : BUF_X1 port map( A => N253, Z => n350_port);
   U704 : BUF_X1 port map( A => N254, Z => n347_port);
   U705 : BUF_X1 port map( A => N255, Z => n344_port);
   U706 : BUF_X1 port map( A => N256, Z => n341_port);
   U707 : BUF_X1 port map( A => N257, Z => n338_port);
   U708 : BUF_X1 port map( A => N258, Z => n335_port);
   U709 : BUF_X1 port map( A => N259, Z => n332_port);
   U710 : BUF_X1 port map( A => N260, Z => n329_port);
   U711 : BUF_X1 port map( A => N261, Z => n326_port);
   U712 : BUF_X1 port map( A => N262, Z => n323_port);
   U713 : BUF_X1 port map( A => N263, Z => n320_port);
   U714 : BUF_X1 port map( A => N264, Z => n317_port);
   U715 : BUF_X1 port map( A => N265, Z => n314_port);
   U716 : BUF_X1 port map( A => N266, Z => n311_port);
   U717 : BUF_X1 port map( A => N267, Z => n308_port);
   U718 : BUF_X1 port map( A => N268, Z => n305_port);
   U719 : BUF_X1 port map( A => N269, Z => n302_port);
   U720 : BUF_X1 port map( A => N270, Z => n299_port);
   U721 : BUF_X1 port map( A => N271, Z => n296_port);
   U722 : BUF_X1 port map( A => N272, Z => n293_port);
   U723 : BUF_X1 port map( A => N273, Z => n290_port);
   U724 : BUF_X1 port map( A => N274, Z => n287_port);
   U725 : BUF_X1 port map( A => N275, Z => n284_port);
   U726 : BUF_X1 port map( A => N244, Z => n376);
   U727 : BUF_X1 port map( A => N245, Z => n373);
   U728 : BUF_X1 port map( A => N246, Z => n370_port);
   U729 : BUF_X1 port map( A => N247, Z => n367_port);
   U730 : BUF_X1 port map( A => N248, Z => n364_port);
   U731 : BUF_X1 port map( A => N249, Z => n361_port);
   U732 : BUF_X1 port map( A => N250, Z => n358_port);
   U733 : BUF_X1 port map( A => N251, Z => n355_port);
   U734 : BUF_X1 port map( A => N252, Z => n352_port);
   U735 : BUF_X1 port map( A => N253, Z => n349_port);
   U736 : BUF_X1 port map( A => N254, Z => n346_port);
   U737 : BUF_X1 port map( A => N255, Z => n343_port);
   U738 : BUF_X1 port map( A => N256, Z => n340_port);
   U739 : BUF_X1 port map( A => N257, Z => n337_port);
   U740 : BUF_X1 port map( A => N258, Z => n334_port);
   U741 : BUF_X1 port map( A => N259, Z => n331_port);
   U742 : BUF_X1 port map( A => N260, Z => n328_port);
   U743 : BUF_X1 port map( A => N261, Z => n325_port);
   U744 : BUF_X1 port map( A => N262, Z => n322_port);
   U745 : BUF_X1 port map( A => N263, Z => n319_port);
   U746 : BUF_X1 port map( A => N264, Z => n316_port);
   U747 : BUF_X1 port map( A => N265, Z => n313_port);
   U748 : BUF_X1 port map( A => N266, Z => n310_port);
   U749 : BUF_X1 port map( A => N267, Z => n307_port);
   U750 : BUF_X1 port map( A => N268, Z => n304_port);
   U751 : BUF_X1 port map( A => N269, Z => n301_port);
   U752 : BUF_X1 port map( A => N270, Z => n298_port);
   U753 : BUF_X1 port map( A => N271, Z => n295_port);
   U754 : BUF_X1 port map( A => N272, Z => n292_port);
   U755 : BUF_X1 port map( A => N273, Z => n289_port);
   U756 : BUF_X1 port map( A => N274, Z => n286_port);
   U757 : BUF_X1 port map( A => N275, Z => n283_port);
   U758 : BUF_X1 port map( A => N244, Z => n378);
   U759 : BUF_X1 port map( A => N245, Z => n375);
   U760 : BUF_X1 port map( A => N246, Z => n372);
   U761 : BUF_X1 port map( A => N247, Z => n369_port);
   U762 : BUF_X1 port map( A => N248, Z => n366_port);
   U763 : BUF_X1 port map( A => N249, Z => n363_port);
   U764 : BUF_X1 port map( A => N250, Z => n360_port);
   U765 : BUF_X1 port map( A => N251, Z => n357_port);
   U766 : BUF_X1 port map( A => N252, Z => n354_port);
   U767 : BUF_X1 port map( A => N253, Z => n351_port);
   U768 : BUF_X1 port map( A => N254, Z => n348_port);
   U769 : BUF_X1 port map( A => N255, Z => n345_port);
   U770 : BUF_X1 port map( A => N256, Z => n342_port);
   U771 : BUF_X1 port map( A => N257, Z => n339_port);
   U772 : BUF_X1 port map( A => N258, Z => n336_port);
   U773 : BUF_X1 port map( A => N259, Z => n333_port);
   U774 : BUF_X1 port map( A => N260, Z => n330_port);
   U775 : BUF_X1 port map( A => N261, Z => n327_port);
   U776 : BUF_X1 port map( A => N262, Z => n324_port);
   U777 : BUF_X1 port map( A => N263, Z => n321_port);
   U778 : BUF_X1 port map( A => N264, Z => n318_port);
   U779 : BUF_X1 port map( A => N265, Z => n315_port);
   U780 : BUF_X1 port map( A => N266, Z => n312_port);
   U781 : BUF_X1 port map( A => N267, Z => n309_port);
   U782 : BUF_X1 port map( A => N268, Z => n306);
   U783 : BUF_X1 port map( A => N269, Z => n303_port);
   U784 : BUF_X1 port map( A => N270, Z => n300_port);
   U785 : BUF_X1 port map( A => N271, Z => n297_port);
   U786 : BUF_X1 port map( A => N272, Z => n294_port);
   U787 : BUF_X1 port map( A => N273, Z => n291_port);
   U788 : BUF_X1 port map( A => N274, Z => n288_port);
   U789 : BUF_X1 port map( A => N275, Z => n285_port);
   U790 : BUF_X1 port map( A => RESET, Z => n387);
   U791 : BUF_X1 port map( A => RESET, Z => n388);
   U792 : OAI221_X1 port map( B1 => n1933, B2 => n93, C1 => n1901, C2 => n90, A
                           => n1315, ZN => n1314);
   U793 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_24_port, B1 => n82, 
                           B2 => REGISTERS_18_24_port, ZN => n1315);
   U794 : OAI221_X1 port map( B1 => n1932, B2 => n93, C1 => n1900, C2 => n90, A
                           => n1297, ZN => n1296);
   U795 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_25_port, B1 => n82, 
                           B2 => REGISTERS_18_25_port, ZN => n1297);
   U796 : OAI221_X1 port map( B1 => n1931, B2 => n93, C1 => n1899, C2 => n90, A
                           => n1279, ZN => n1278);
   U797 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_26_port, B1 => n82, 
                           B2 => REGISTERS_18_26_port, ZN => n1279);
   U798 : OAI221_X1 port map( B1 => n1930, B2 => n93, C1 => n1898, C2 => n90, A
                           => n1261, ZN => n1260);
   U799 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_27_port, B1 => n82, 
                           B2 => REGISTERS_18_27_port, ZN => n1261);
   U800 : OAI221_X1 port map( B1 => n1929, B2 => n93, C1 => n1897, C2 => n90, A
                           => n1243, ZN => n1242);
   U801 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_28_port, B1 => n82, 
                           B2 => REGISTERS_18_28_port, ZN => n1243);
   U802 : OAI221_X1 port map( B1 => n1928, B2 => n93, C1 => n1896, C2 => n90, A
                           => n1225, ZN => n1224);
   U803 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_29_port, B1 => n82, 
                           B2 => REGISTERS_18_29_port, ZN => n1225);
   U804 : OAI221_X1 port map( B1 => n1927, B2 => n93, C1 => n1895, C2 => n90, A
                           => n1207, ZN => n1206);
   U805 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_30_port, B1 => n82, 
                           B2 => REGISTERS_18_30_port, ZN => n1207);
   U806 : OAI221_X1 port map( B1 => n1926, B2 => n93, C1 => n1894, C2 => n90, A
                           => n1159, ZN => n1156);
   U807 : AOI22_X1 port map( A1 => n87, A2 => REGISTERS_19_31_port, B1 => n82, 
                           B2 => REGISTERS_18_31_port, ZN => n1159);
   U808 : OAI221_X1 port map( B1 => n1997, B2 => n81, C1 => n1965, C2 => n78, A
                           => n1316, ZN => n1313);
   U809 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_24_port, B1 => n70, 
                           B2 => REGISTERS_22_24_port, ZN => n1316);
   U810 : OAI221_X1 port map( B1 => n483, B2 => n36, C1 => n451, C2 => n33, A 
                           => n1324, ZN => n1321);
   U811 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_24_port, B1 => n25, 
                           B2 => REGISTERS_6_24_port, ZN => n1324);
   U812 : OAI221_X1 port map( B1 => n1996, B2 => n81, C1 => n1964, C2 => n78, A
                           => n1298, ZN => n1295);
   U813 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_25_port, B1 => n70, 
                           B2 => REGISTERS_22_25_port, ZN => n1298);
   U814 : OAI221_X1 port map( B1 => n482, B2 => n36, C1 => n450, C2 => n33, A 
                           => n1306, ZN => n1303);
   U815 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_25_port, B1 => n25, 
                           B2 => REGISTERS_6_25_port, ZN => n1306);
   U816 : OAI221_X1 port map( B1 => n1995, B2 => n81, C1 => n1963, C2 => n78, A
                           => n1280, ZN => n1277);
   U817 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_26_port, B1 => n70, 
                           B2 => REGISTERS_22_26_port, ZN => n1280);
   U818 : OAI221_X1 port map( B1 => n481, B2 => n36, C1 => n449, C2 => n33, A 
                           => n1288, ZN => n1285);
   U819 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_26_port, B1 => n25, 
                           B2 => REGISTERS_6_26_port, ZN => n1288);
   U820 : OAI221_X1 port map( B1 => n1994, B2 => n81, C1 => n1962, C2 => n78, A
                           => n1262, ZN => n1259);
   U821 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_27_port, B1 => n70, 
                           B2 => REGISTERS_22_27_port, ZN => n1262);
   U822 : OAI221_X1 port map( B1 => n480, B2 => n36, C1 => n448, C2 => n33, A 
                           => n1270, ZN => n1267);
   U823 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_27_port, B1 => n25, 
                           B2 => REGISTERS_6_27_port, ZN => n1270);
   U824 : OAI221_X1 port map( B1 => n1993, B2 => n81, C1 => n1961, C2 => n78, A
                           => n1244, ZN => n1241);
   U825 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_28_port, B1 => n70, 
                           B2 => REGISTERS_22_28_port, ZN => n1244);
   U826 : OAI221_X1 port map( B1 => n479, B2 => n36, C1 => n447, C2 => n33, A 
                           => n1252, ZN => n1249);
   U827 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_28_port, B1 => n25, 
                           B2 => REGISTERS_6_28_port, ZN => n1252);
   U828 : OAI221_X1 port map( B1 => n1992, B2 => n81, C1 => n1960, C2 => n78, A
                           => n1226, ZN => n1223);
   U829 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_29_port, B1 => n70, 
                           B2 => REGISTERS_22_29_port, ZN => n1226);
   U830 : OAI221_X1 port map( B1 => n478, B2 => n36, C1 => n446, C2 => n33, A 
                           => n1234, ZN => n1231);
   U831 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_29_port, B1 => n25, 
                           B2 => REGISTERS_6_29_port, ZN => n1234);
   U832 : OAI221_X1 port map( B1 => n1991, B2 => n81, C1 => n1959, C2 => n78, A
                           => n1208, ZN => n1205);
   U833 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_30_port, B1 => n70, 
                           B2 => REGISTERS_22_30_port, ZN => n1208);
   U834 : OAI221_X1 port map( B1 => n477, B2 => n36, C1 => n445, C2 => n33, A 
                           => n1216, ZN => n1213);
   U835 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_30_port, B1 => n25, 
                           B2 => REGISTERS_6_30_port, ZN => n1216);
   U836 : OAI221_X1 port map( B1 => n1990, B2 => n81, C1 => n1958, C2 => n78, A
                           => n1164, ZN => n1155);
   U837 : AOI22_X1 port map( A1 => n75, A2 => REGISTERS_23_31_port, B1 => n70, 
                           B2 => REGISTERS_22_31_port, ZN => n1164);
   U838 : OAI221_X1 port map( B1 => n476, B2 => n36, C1 => n444, C2 => n33, A 
                           => n1188, ZN => n1179);
   U839 : AOI22_X1 port map( A1 => n30, A2 => REGISTERS_7_31_port, B1 => n25, 
                           B2 => REGISTERS_6_31_port, ZN => n1188);
   U840 : OAI221_X1 port map( B1 => n499, B2 => n34, C1 => n467, C2 => n31, A 
                           => n1612, ZN => n1609);
   U841 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_8_port, B1 => n26, B2
                           => REGISTERS_6_8_port, ZN => n1612);
   U842 : OAI221_X1 port map( B1 => n498, B2 => n34, C1 => n466, C2 => n31, A 
                           => n1594, ZN => n1591);
   U843 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_9_port, B1 => n26, B2
                           => REGISTERS_6_9_port, ZN => n1594);
   U844 : OAI221_X1 port map( B1 => n497, B2 => n34, C1 => n465, C2 => n31, A 
                           => n1576, ZN => n1573);
   U845 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_10_port, B1 => n26, 
                           B2 => REGISTERS_6_10_port, ZN => n1576);
   U846 : OAI221_X1 port map( B1 => n496, B2 => n34, C1 => n464, C2 => n31, A 
                           => n1558, ZN => n1555);
   U847 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_11_port, B1 => n26, 
                           B2 => REGISTERS_6_11_port, ZN => n1558);
   U848 : OAI221_X1 port map( B1 => n495, B2 => n35, C1 => n463, C2 => n32, A 
                           => n1540, ZN => n1537);
   U849 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_12_port, B1 => n26, 
                           B2 => REGISTERS_6_12_port, ZN => n1540);
   U850 : OAI221_X1 port map( B1 => n494, B2 => n35, C1 => n462, C2 => n32, A 
                           => n1522, ZN => n1519);
   U851 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_13_port, B1 => n26, 
                           B2 => REGISTERS_6_13_port, ZN => n1522);
   U852 : OAI221_X1 port map( B1 => n493, B2 => n35, C1 => n461, C2 => n32, A 
                           => n1504, ZN => n1501);
   U853 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_14_port, B1 => n26, 
                           B2 => REGISTERS_6_14_port, ZN => n1504);
   U854 : OAI221_X1 port map( B1 => n492, B2 => n35, C1 => n460, C2 => n32, A 
                           => n1486, ZN => n1483);
   U855 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_15_port, B1 => n26, 
                           B2 => REGISTERS_6_15_port, ZN => n1486);
   U856 : OAI221_X1 port map( B1 => n491, B2 => n35, C1 => n459, C2 => n32, A 
                           => n1468, ZN => n1465);
   U857 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_16_port, B1 => n26, 
                           B2 => REGISTERS_6_16_port, ZN => n1468);
   U858 : OAI221_X1 port map( B1 => n490, B2 => n35, C1 => n458, C2 => n32, A 
                           => n1450, ZN => n1447);
   U859 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_17_port, B1 => n26, 
                           B2 => REGISTERS_6_17_port, ZN => n1450);
   U860 : OAI221_X1 port map( B1 => n489, B2 => n35, C1 => n457, C2 => n32, A 
                           => n1432, ZN => n1429);
   U861 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_18_port, B1 => n26, 
                           B2 => REGISTERS_6_18_port, ZN => n1432);
   U862 : OAI221_X1 port map( B1 => n488, B2 => n35, C1 => n456, C2 => n32, A 
                           => n1414, ZN => n1411);
   U863 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_19_port, B1 => n26, 
                           B2 => REGISTERS_6_19_port, ZN => n1414);
   U864 : OAI221_X1 port map( B1 => n487, B2 => n35, C1 => n455, C2 => n32, A 
                           => n1396, ZN => n1393);
   U865 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_20_port, B1 => n25, 
                           B2 => REGISTERS_6_20_port, ZN => n1396);
   U866 : OAI221_X1 port map( B1 => n486, B2 => n35, C1 => n454, C2 => n32, A 
                           => n1378, ZN => n1375);
   U867 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_21_port, B1 => n25, 
                           B2 => REGISTERS_6_21_port, ZN => n1378);
   U868 : OAI221_X1 port map( B1 => n485, B2 => n35, C1 => n453, C2 => n32, A 
                           => n1360, ZN => n1357);
   U869 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_22_port, B1 => n25, 
                           B2 => REGISTERS_6_22_port, ZN => n1360);
   U870 : OAI221_X1 port map( B1 => n484, B2 => n35, C1 => n452, C2 => n32, A 
                           => n1342, ZN => n1339);
   U871 : AOI22_X1 port map( A1 => n29, A2 => REGISTERS_7_23_port, B1 => n25, 
                           B2 => REGISTERS_6_23_port, ZN => n1342);
   U872 : OAI221_X1 port map( B1 => n186, B2 => n1933, C1 => n183, C2 => n1901,
                           A => n691, ZN => n690);
   U873 : AOI22_X1 port map( A1 => REGISTERS_19_24_port, A2 => n180, B1 => 
                           REGISTERS_18_24_port, B2 => n177, ZN => n691);
   U874 : OAI221_X1 port map( B1 => n174, B2 => n1997, C1 => n171, C2 => n1965,
                           A => n692, ZN => n689);
   U875 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n168, B1 => 
                           REGISTERS_22_24_port, B2 => n165, ZN => n692);
   U876 : OAI221_X1 port map( B1 => n162, B2 => n2061, C1 => n159, C2 => n2029,
                           A => n693, ZN => n688);
   U877 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n156, B1 => 
                           REGISTERS_26_24_port, B2 => n153, ZN => n693);
   U878 : OAI221_X1 port map( B1 => n150, B2 => n2125, C1 => n147, C2 => n2093,
                           A => n694, ZN => n687);
   U879 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n144, B1 => 
                           REGISTERS_28_24_port, B2 => n141, ZN => n694);
   U880 : OAI221_X1 port map( B1 => n117, B2 => n1805, C1 => n114, C2 => n515, 
                           A => n701, ZN => n696);
   U881 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n111, B1 => 
                           REGISTERS_10_24_port, B2 => n108, ZN => n701);
   U882 : OAI221_X1 port map( B1 => n129, B2 => n483, C1 => n126, C2 => n451, A
                           => n700, ZN => n697);
   U883 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n123, B1 => 
                           REGISTERS_6_24_port, B2 => n120, ZN => n700);
   U884 : OAI221_X1 port map( B1 => n105, B2 => n1869, C1 => n102, C2 => n1837,
                           A => n702, ZN => n695);
   U885 : AOI22_X1 port map( A1 => REGISTERS_15_24_port, A2 => n99, B1 => 
                           REGISTERS_14_24_port, B2 => n96, ZN => n702);
   U886 : OAI221_X1 port map( B1 => n186, B2 => n1932, C1 => n183, C2 => n1900,
                           A => n673, ZN => n672);
   U887 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n180, B1 => 
                           REGISTERS_18_25_port, B2 => n177, ZN => n673);
   U888 : OAI221_X1 port map( B1 => n174, B2 => n1996, C1 => n171, C2 => n1964,
                           A => n674, ZN => n671);
   U889 : AOI22_X1 port map( A1 => REGISTERS_23_25_port, A2 => n168, B1 => 
                           REGISTERS_22_25_port, B2 => n165, ZN => n674);
   U890 : OAI221_X1 port map( B1 => n162, B2 => n2060, C1 => n159, C2 => n2028,
                           A => n675, ZN => n670);
   U891 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n156, B1 => 
                           REGISTERS_26_25_port, B2 => n153, ZN => n675);
   U892 : OAI221_X1 port map( B1 => n150, B2 => n2124, C1 => n147, C2 => n2092,
                           A => n676, ZN => n669);
   U893 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n144, B1 => 
                           REGISTERS_28_25_port, B2 => n141, ZN => n676);
   U894 : OAI221_X1 port map( B1 => n117, B2 => n1804, C1 => n114, C2 => n514, 
                           A => n683, ZN => n678);
   U895 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n111, B1 => 
                           REGISTERS_10_25_port, B2 => n108, ZN => n683);
   U896 : OAI221_X1 port map( B1 => n129, B2 => n482, C1 => n126, C2 => n450, A
                           => n682, ZN => n679);
   U897 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n123, B1 => 
                           REGISTERS_6_25_port, B2 => n120, ZN => n682);
   U898 : OAI221_X1 port map( B1 => n105, B2 => n1868, C1 => n102, C2 => n1836,
                           A => n684, ZN => n677);
   U899 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n99, B1 => 
                           REGISTERS_14_25_port, B2 => n96, ZN => n684);
   U900 : OAI221_X1 port map( B1 => n186, B2 => n1931, C1 => n183, C2 => n1899,
                           A => n655, ZN => n654);
   U901 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n180, B1 => 
                           REGISTERS_18_26_port, B2 => n177, ZN => n655);
   U902 : OAI221_X1 port map( B1 => n174, B2 => n1995, C1 => n171, C2 => n1963,
                           A => n656, ZN => n653);
   U903 : AOI22_X1 port map( A1 => REGISTERS_23_26_port, A2 => n168, B1 => 
                           REGISTERS_22_26_port, B2 => n165, ZN => n656);
   U904 : OAI221_X1 port map( B1 => n162, B2 => n2059, C1 => n159, C2 => n2027,
                           A => n657, ZN => n652);
   U905 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n156, B1 => 
                           REGISTERS_26_26_port, B2 => n153, ZN => n657);
   U906 : OAI221_X1 port map( B1 => n150, B2 => n2123, C1 => n147, C2 => n2091,
                           A => n658, ZN => n651);
   U907 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n144, B1 => 
                           REGISTERS_28_26_port, B2 => n141, ZN => n658);
   U908 : OAI221_X1 port map( B1 => n117, B2 => n1803, C1 => n114, C2 => n513, 
                           A => n665, ZN => n660);
   U909 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n111, B1 => 
                           REGISTERS_10_26_port, B2 => n108, ZN => n665);
   U910 : OAI221_X1 port map( B1 => n129, B2 => n481, C1 => n126, C2 => n449, A
                           => n664, ZN => n661);
   U911 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n123, B1 => 
                           REGISTERS_6_26_port, B2 => n120, ZN => n664);
   U912 : OAI221_X1 port map( B1 => n105, B2 => n1867, C1 => n102, C2 => n1835,
                           A => n666, ZN => n659);
   U913 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n99, B1 => 
                           REGISTERS_14_26_port, B2 => n96, ZN => n666);
   U914 : OAI221_X1 port map( B1 => n186, B2 => n1930, C1 => n183, C2 => n1898,
                           A => n637, ZN => n636);
   U915 : AOI22_X1 port map( A1 => REGISTERS_19_27_port, A2 => n180, B1 => 
                           REGISTERS_18_27_port, B2 => n177, ZN => n637);
   U916 : OAI221_X1 port map( B1 => n174, B2 => n1994, C1 => n171, C2 => n1962,
                           A => n638, ZN => n635);
   U917 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n168, B1 => 
                           REGISTERS_22_27_port, B2 => n165, ZN => n638);
   U918 : OAI221_X1 port map( B1 => n162, B2 => n2058, C1 => n159, C2 => n2026,
                           A => n639, ZN => n634);
   U919 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n156, B1 => 
                           REGISTERS_26_27_port, B2 => n153, ZN => n639);
   U920 : OAI221_X1 port map( B1 => n150, B2 => n2122, C1 => n147, C2 => n2090,
                           A => n640, ZN => n633);
   U921 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n144, B1 => 
                           REGISTERS_28_27_port, B2 => n141, ZN => n640);
   U922 : OAI221_X1 port map( B1 => n117, B2 => n1802, C1 => n114, C2 => n512, 
                           A => n647, ZN => n642);
   U923 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n111, B1 => 
                           REGISTERS_10_27_port, B2 => n108, ZN => n647);
   U924 : OAI221_X1 port map( B1 => n129, B2 => n480, C1 => n126, C2 => n448, A
                           => n646, ZN => n643);
   U925 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n123, B1 => 
                           REGISTERS_6_27_port, B2 => n120, ZN => n646);
   U926 : OAI221_X1 port map( B1 => n105, B2 => n1866, C1 => n102, C2 => n1834,
                           A => n648, ZN => n641);
   U927 : AOI22_X1 port map( A1 => REGISTERS_15_27_port, A2 => n99, B1 => 
                           REGISTERS_14_27_port, B2 => n96, ZN => n648);
   U928 : OAI221_X1 port map( B1 => n186, B2 => n1929, C1 => n183, C2 => n1897,
                           A => n619, ZN => n618);
   U929 : AOI22_X1 port map( A1 => REGISTERS_19_28_port, A2 => n180, B1 => 
                           REGISTERS_18_28_port, B2 => n177, ZN => n619);
   U930 : OAI221_X1 port map( B1 => n174, B2 => n1993, C1 => n171, C2 => n1961,
                           A => n620, ZN => n617);
   U931 : AOI22_X1 port map( A1 => REGISTERS_23_28_port, A2 => n168, B1 => 
                           REGISTERS_22_28_port, B2 => n165, ZN => n620);
   U932 : OAI221_X1 port map( B1 => n162, B2 => n2057, C1 => n159, C2 => n2025,
                           A => n621, ZN => n616);
   U933 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n156, B1 => 
                           REGISTERS_26_28_port, B2 => n153, ZN => n621);
   U934 : OAI221_X1 port map( B1 => n150, B2 => n2121, C1 => n147, C2 => n2089,
                           A => n622, ZN => n615);
   U935 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n144, B1 => 
                           REGISTERS_28_28_port, B2 => n141, ZN => n622);
   U936 : OAI221_X1 port map( B1 => n117, B2 => n1801, C1 => n114, C2 => n511, 
                           A => n629, ZN => n624);
   U937 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n111, B1 => 
                           REGISTERS_10_28_port, B2 => n108, ZN => n629);
   U938 : OAI221_X1 port map( B1 => n129, B2 => n479, C1 => n126, C2 => n447, A
                           => n628, ZN => n625);
   U939 : AOI22_X1 port map( A1 => REGISTERS_7_28_port, A2 => n123, B1 => 
                           REGISTERS_6_28_port, B2 => n120, ZN => n628);
   U940 : OAI221_X1 port map( B1 => n105, B2 => n1865, C1 => n102, C2 => n1833,
                           A => n630, ZN => n623);
   U941 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n99, B1 => 
                           REGISTERS_14_28_port, B2 => n96, ZN => n630);
   U942 : OAI221_X1 port map( B1 => n186, B2 => n1928, C1 => n183, C2 => n1896,
                           A => n601, ZN => n600);
   U943 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n180, B1 => 
                           REGISTERS_18_29_port, B2 => n177, ZN => n601);
   U944 : OAI221_X1 port map( B1 => n174, B2 => n1992, C1 => n171, C2 => n1960,
                           A => n602, ZN => n599);
   U945 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n168, B1 => 
                           REGISTERS_22_29_port, B2 => n165, ZN => n602);
   U946 : OAI221_X1 port map( B1 => n162, B2 => n2056, C1 => n159, C2 => n2024,
                           A => n603, ZN => n598);
   U947 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n156, B1 => 
                           REGISTERS_26_29_port, B2 => n153, ZN => n603);
   U948 : OAI221_X1 port map( B1 => n150, B2 => n2120, C1 => n147, C2 => n2088,
                           A => n604, ZN => n597);
   U949 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n144, B1 => 
                           REGISTERS_28_29_port, B2 => n141, ZN => n604);
   U950 : OAI221_X1 port map( B1 => n117, B2 => n1800, C1 => n114, C2 => n510, 
                           A => n611, ZN => n606);
   U951 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n111, B1 => 
                           REGISTERS_10_29_port, B2 => n108, ZN => n611);
   U952 : OAI221_X1 port map( B1 => n129, B2 => n478, C1 => n126, C2 => n446, A
                           => n610, ZN => n607);
   U953 : AOI22_X1 port map( A1 => REGISTERS_7_29_port, A2 => n123, B1 => 
                           REGISTERS_6_29_port, B2 => n120, ZN => n610);
   U954 : OAI221_X1 port map( B1 => n105, B2 => n1864, C1 => n102, C2 => n1832,
                           A => n612, ZN => n605);
   U955 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n99, B1 => 
                           REGISTERS_14_29_port, B2 => n96, ZN => n612);
   U956 : OAI221_X1 port map( B1 => n186, B2 => n1927, C1 => n183, C2 => n1895,
                           A => n583, ZN => n582);
   U957 : AOI22_X1 port map( A1 => REGISTERS_19_30_port, A2 => n180, B1 => 
                           REGISTERS_18_30_port, B2 => n177, ZN => n583);
   U958 : OAI221_X1 port map( B1 => n174, B2 => n1991, C1 => n171, C2 => n1959,
                           A => n584, ZN => n581);
   U959 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n168, B1 => 
                           REGISTERS_22_30_port, B2 => n165, ZN => n584);
   U960 : OAI221_X1 port map( B1 => n162, B2 => n2055, C1 => n159, C2 => n2023,
                           A => n585, ZN => n580);
   U961 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n156, B1 => 
                           REGISTERS_26_30_port, B2 => n153, ZN => n585);
   U962 : OAI221_X1 port map( B1 => n150, B2 => n2119, C1 => n147, C2 => n2087,
                           A => n586, ZN => n579);
   U963 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n144, B1 => 
                           REGISTERS_28_30_port, B2 => n141, ZN => n586);
   U964 : OAI221_X1 port map( B1 => n117, B2 => n1799, C1 => n114, C2 => n509, 
                           A => n593, ZN => n588);
   U965 : AOI22_X1 port map( A1 => REGISTERS_11_30_port, A2 => n111, B1 => 
                           REGISTERS_10_30_port, B2 => n108, ZN => n593);
   U966 : OAI221_X1 port map( B1 => n129, B2 => n477, C1 => n126, C2 => n445, A
                           => n592, ZN => n589);
   U967 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n123, B1 => 
                           REGISTERS_6_30_port, B2 => n120, ZN => n592);
   U968 : OAI221_X1 port map( B1 => n105, B2 => n1863, C1 => n102, C2 => n1831,
                           A => n594, ZN => n587);
   U969 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n99, B1 => 
                           REGISTERS_14_30_port, B2 => n96, ZN => n594);
   U970 : OAI221_X1 port map( B1 => n186, B2 => n1926, C1 => n183, C2 => n1894,
                           A => n535, ZN => n532);
   U971 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n180, B1 => 
                           REGISTERS_18_31_port, B2 => n177, ZN => n535);
   U972 : OAI221_X1 port map( B1 => n174, B2 => n1990, C1 => n171, C2 => n1958,
                           A => n540, ZN => n531);
   U973 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n168, B1 => 
                           REGISTERS_22_31_port, B2 => n165, ZN => n540);
   U974 : OAI221_X1 port map( B1 => n162, B2 => n2054, C1 => n159, C2 => n2022,
                           A => n545, ZN => n530);
   U975 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n156, B1 => 
                           REGISTERS_26_31_port, B2 => n153, ZN => n545);
   U976 : OAI221_X1 port map( B1 => n150, B2 => n2118, C1 => n147, C2 => n2086,
                           A => n550, ZN => n529);
   U977 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n144, B1 => 
                           REGISTERS_28_31_port, B2 => n141, ZN => n550);
   U978 : OAI221_X1 port map( B1 => n117, B2 => n1798, C1 => n114, C2 => n508, 
                           A => n569, ZN => n554);
   U979 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n111, B1 => 
                           REGISTERS_10_31_port, B2 => n108, ZN => n569);
   U980 : OAI221_X1 port map( B1 => n129, B2 => n476, C1 => n126, C2 => n444, A
                           => n564, ZN => n555);
   U981 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n123, B1 => 
                           REGISTERS_6_31_port, B2 => n120, ZN => n564);
   U982 : OAI221_X1 port map( B1 => n105, B2 => n1862, C1 => n102, C2 => n1830,
                           A => n574, ZN => n553);
   U983 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n99, B1 => 
                           REGISTERS_14_31_port, B2 => n96, ZN => n574);
   U984 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_0_port, B1 => n3, B2 
                           => REGISTERS_14_0_port, ZN => n1773);
   U985 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_1_port, B1 => n3, B2 
                           => REGISTERS_14_1_port, ZN => n1740);
   U986 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_2_port, B1 => n3, B2 
                           => REGISTERS_14_2_port, ZN => n1722);
   U987 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_3_port, B1 => n3, B2 
                           => REGISTERS_14_3_port, ZN => n1704);
   U988 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_4_port, B1 => n3, B2 
                           => REGISTERS_14_4_port, ZN => n1686);
   U989 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_5_port, B1 => n3, B2 
                           => REGISTERS_14_5_port, ZN => n1668);
   U990 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_6_port, B1 => n3, B2 
                           => REGISTERS_14_6_port, ZN => n1650);
   U991 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_7_port, B1 => n3, B2 
                           => REGISTERS_14_7_port, ZN => n1632);
   U992 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_8_port, B1 => n2, B2 
                           => REGISTERS_14_8_port, ZN => n1614);
   U993 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_9_port, B1 => n2, B2 
                           => REGISTERS_14_9_port, ZN => n1596);
   U994 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_10_port, B1 => n2, B2
                           => REGISTERS_14_10_port, ZN => n1578);
   U995 : AOI22_X1 port map( A1 => n4, A2 => REGISTERS_15_11_port, B1 => n2, B2
                           => REGISTERS_14_11_port, ZN => n1560);
   U996 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_12_port, B1 => n2, B2
                           => REGISTERS_14_12_port, ZN => n1542);
   U997 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_13_port, B1 => n2, B2
                           => REGISTERS_14_13_port, ZN => n1524);
   U998 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_14_port, B1 => n2, B2
                           => REGISTERS_14_14_port, ZN => n1506);
   U999 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_15_port, B1 => n2, B2
                           => REGISTERS_14_15_port, ZN => n1488);
   U1000 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_16_port, B1 => n2, 
                           B2 => REGISTERS_14_16_port, ZN => n1470);
   U1001 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_17_port, B1 => n2, 
                           B2 => REGISTERS_14_17_port, ZN => n1452);
   U1002 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_18_port, B1 => n2, 
                           B2 => REGISTERS_14_18_port, ZN => n1434);
   U1003 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_19_port, B1 => n2, 
                           B2 => REGISTERS_14_19_port, ZN => n1416);
   U1004 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_20_port, B1 => n1, 
                           B2 => REGISTERS_14_20_port, ZN => n1398);
   U1005 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_21_port, B1 => n1, 
                           B2 => REGISTERS_14_21_port, ZN => n1380);
   U1006 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_22_port, B1 => n1, 
                           B2 => REGISTERS_14_22_port, ZN => n1362);
   U1007 : AOI22_X1 port map( A1 => n5, A2 => REGISTERS_15_23_port, B1 => n1, 
                           B2 => REGISTERS_14_23_port, ZN => n1344);
   U1008 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_24_port, B1 => n1, 
                           B2 => REGISTERS_14_24_port, ZN => n1326);
   U1009 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_25_port, B1 => n1, 
                           B2 => REGISTERS_14_25_port, ZN => n1308);
   U1010 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_26_port, B1 => n1, 
                           B2 => REGISTERS_14_26_port, ZN => n1290);
   U1011 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_27_port, B1 => n1, 
                           B2 => REGISTERS_14_27_port, ZN => n1272);
   U1012 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_28_port, B1 => n1, 
                           B2 => REGISTERS_14_28_port, ZN => n1254);
   U1013 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_29_port, B1 => n1, 
                           B2 => REGISTERS_14_29_port, ZN => n1236);
   U1014 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_30_port, B1 => n1, 
                           B2 => REGISTERS_14_30_port, ZN => n1218);
   U1015 : AOI22_X1 port map( A1 => n6, A2 => REGISTERS_15_31_port, B1 => n1, 
                           B2 => REGISTERS_14_31_port, ZN => n1198);
   U1016 : OAI221_X1 port map( B1 => n184, B2 => n1957, C1 => n181, C2 => n1925
                           , A => n1123, ZN => n1122);
   U1017 : AOI22_X1 port map( A1 => REGISTERS_19_0_port, A2 => n178, B1 => 
                           REGISTERS_18_0_port, B2 => n175, ZN => n1123);
   U1018 : OAI221_X1 port map( B1 => n172, B2 => n2021, C1 => n169, C2 => n1989
                           , A => n1128, ZN => n1121);
   U1019 : AOI22_X1 port map( A1 => REGISTERS_23_0_port, A2 => n166, B1 => 
                           REGISTERS_22_0_port, B2 => n163, ZN => n1128);
   U1020 : OAI221_X1 port map( B1 => n160, B2 => n2085, C1 => n157, C2 => n2053
                           , A => n1132, ZN => n1120);
   U1021 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n154, B1 => 
                           REGISTERS_26_0_port, B2 => n151, ZN => n1132);
   U1022 : OAI221_X1 port map( B1 => n148, B2 => n2149, C1 => n145, C2 => n2117
                           , A => n1135, ZN => n1119);
   U1023 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n142, B1 => 
                           REGISTERS_28_0_port, B2 => n139, ZN => n1135);
   U1024 : OAI221_X1 port map( B1 => n115, B2 => n1829, C1 => n112, C2 => n1797
                           , A => n1146, ZN => n1138);
   U1025 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n109, B1 => 
                           REGISTERS_10_0_port, B2 => n106, ZN => n1146);
   U1026 : OAI221_X1 port map( B1 => n127, B2 => n507, C1 => n124, C2 => n475, 
                           A => n1144, ZN => n1139);
   U1027 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n121, B1 => 
                           REGISTERS_6_0_port, B2 => n118, ZN => n1144);
   U1028 : OAI221_X1 port map( B1 => n103, B2 => n1893, C1 => n100, C2 => n1861
                           , A => n1149, ZN => n1137);
   U1029 : AOI22_X1 port map( A1 => REGISTERS_15_0_port, A2 => n97, B1 => 
                           REGISTERS_14_0_port, B2 => n94, ZN => n1149);
   U1030 : OAI221_X1 port map( B1 => n184, B2 => n1956, C1 => n181, C2 => n1924
                           , A => n1105, ZN => n1104);
   U1031 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n178, B1 => 
                           REGISTERS_18_1_port, B2 => n175, ZN => n1105);
   U1032 : OAI221_X1 port map( B1 => n172, B2 => n2020, C1 => n169, C2 => n1988
                           , A => n1106, ZN => n1103);
   U1033 : AOI22_X1 port map( A1 => REGISTERS_23_1_port, A2 => n166, B1 => 
                           REGISTERS_22_1_port, B2 => n163, ZN => n1106);
   U1034 : OAI221_X1 port map( B1 => n160, B2 => n2084, C1 => n157, C2 => n2052
                           , A => n1107, ZN => n1102);
   U1035 : AOI22_X1 port map( A1 => REGISTERS_27_1_port, A2 => n154, B1 => 
                           REGISTERS_26_1_port, B2 => n151, ZN => n1107);
   U1036 : OAI221_X1 port map( B1 => n148, B2 => n2148, C1 => n145, C2 => n2116
                           , A => n1108, ZN => n1101);
   U1037 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n142, B1 => 
                           REGISTERS_28_1_port, B2 => n139, ZN => n1108);
   U1038 : OAI221_X1 port map( B1 => n115, B2 => n1828, C1 => n112, C2 => n1796
                           , A => n1115, ZN => n1110);
   U1039 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n109, B1 => 
                           REGISTERS_10_1_port, B2 => n106, ZN => n1115);
   U1040 : OAI221_X1 port map( B1 => n127, B2 => n506, C1 => n124, C2 => n474, 
                           A => n1114, ZN => n1111);
   U1041 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n121, B1 => 
                           REGISTERS_6_1_port, B2 => n118, ZN => n1114);
   U1042 : OAI221_X1 port map( B1 => n103, B2 => n1892, C1 => n100, C2 => n1860
                           , A => n1116, ZN => n1109);
   U1043 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n97, B1 => 
                           REGISTERS_14_1_port, B2 => n94, ZN => n1116);
   U1044 : OAI221_X1 port map( B1 => n184, B2 => n1955, C1 => n181, C2 => n1923
                           , A => n1087, ZN => n1086);
   U1045 : AOI22_X1 port map( A1 => REGISTERS_19_2_port, A2 => n178, B1 => 
                           REGISTERS_18_2_port, B2 => n175, ZN => n1087);
   U1046 : OAI221_X1 port map( B1 => n172, B2 => n2019, C1 => n169, C2 => n1987
                           , A => n1088, ZN => n1085);
   U1047 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n166, B1 => 
                           REGISTERS_22_2_port, B2 => n163, ZN => n1088);
   U1048 : OAI221_X1 port map( B1 => n160, B2 => n2083, C1 => n157, C2 => n2051
                           , A => n1089, ZN => n1084);
   U1049 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n154, B1 => 
                           REGISTERS_26_2_port, B2 => n151, ZN => n1089);
   U1050 : OAI221_X1 port map( B1 => n148, B2 => n2147, C1 => n145, C2 => n2115
                           , A => n1090, ZN => n1083);
   U1051 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n142, B1 => 
                           REGISTERS_28_2_port, B2 => n139, ZN => n1090);
   U1052 : OAI221_X1 port map( B1 => n115, B2 => n1827, C1 => n112, C2 => n1795
                           , A => n1097, ZN => n1092);
   U1053 : AOI22_X1 port map( A1 => REGISTERS_11_2_port, A2 => n109, B1 => 
                           REGISTERS_10_2_port, B2 => n106, ZN => n1097);
   U1054 : OAI221_X1 port map( B1 => n127, B2 => n505, C1 => n124, C2 => n473, 
                           A => n1096, ZN => n1093);
   U1055 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n121, B1 => 
                           REGISTERS_6_2_port, B2 => n118, ZN => n1096);
   U1056 : OAI221_X1 port map( B1 => n103, B2 => n1891, C1 => n100, C2 => n1859
                           , A => n1098, ZN => n1091);
   U1057 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n97, B1 => 
                           REGISTERS_14_2_port, B2 => n94, ZN => n1098);
   U1058 : OAI221_X1 port map( B1 => n184, B2 => n1954, C1 => n181, C2 => n1922
                           , A => n1069, ZN => n1068);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n178, B1 => 
                           REGISTERS_18_3_port, B2 => n175, ZN => n1069);
   U1060 : OAI221_X1 port map( B1 => n172, B2 => n2018, C1 => n169, C2 => n1986
                           , A => n1070, ZN => n1067);
   U1061 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n166, B1 => 
                           REGISTERS_22_3_port, B2 => n163, ZN => n1070);
   U1062 : OAI221_X1 port map( B1 => n160, B2 => n2082, C1 => n157, C2 => n2050
                           , A => n1071, ZN => n1066);
   U1063 : AOI22_X1 port map( A1 => REGISTERS_27_3_port, A2 => n154, B1 => 
                           REGISTERS_26_3_port, B2 => n151, ZN => n1071);
   U1064 : OAI221_X1 port map( B1 => n148, B2 => n2146, C1 => n145, C2 => n2114
                           , A => n1072, ZN => n1065);
   U1065 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n142, B1 => 
                           REGISTERS_28_3_port, B2 => n139, ZN => n1072);
   U1066 : OAI221_X1 port map( B1 => n115, B2 => n1826, C1 => n112, C2 => n1794
                           , A => n1079, ZN => n1074);
   U1067 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n109, B1 => 
                           REGISTERS_10_3_port, B2 => n106, ZN => n1079);
   U1068 : OAI221_X1 port map( B1 => n127, B2 => n504, C1 => n124, C2 => n472, 
                           A => n1078, ZN => n1075);
   U1069 : AOI22_X1 port map( A1 => REGISTERS_7_3_port, A2 => n121, B1 => 
                           REGISTERS_6_3_port, B2 => n118, ZN => n1078);
   U1070 : OAI221_X1 port map( B1 => n103, B2 => n1890, C1 => n100, C2 => n1858
                           , A => n1080, ZN => n1073);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_15_3_port, A2 => n97, B1 => 
                           REGISTERS_14_3_port, B2 => n94, ZN => n1080);
   U1072 : OAI221_X1 port map( B1 => n184, B2 => n1953, C1 => n181, C2 => n1921
                           , A => n1051, ZN => n1050);
   U1073 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n178, B1 => 
                           REGISTERS_18_4_port, B2 => n175, ZN => n1051);
   U1074 : OAI221_X1 port map( B1 => n172, B2 => n2017, C1 => n169, C2 => n1985
                           , A => n1052, ZN => n1049);
   U1075 : AOI22_X1 port map( A1 => REGISTERS_23_4_port, A2 => n166, B1 => 
                           REGISTERS_22_4_port, B2 => n163, ZN => n1052);
   U1076 : OAI221_X1 port map( B1 => n160, B2 => n2081, C1 => n157, C2 => n2049
                           , A => n1053, ZN => n1048);
   U1077 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n154, B1 => 
                           REGISTERS_26_4_port, B2 => n151, ZN => n1053);
   U1078 : OAI221_X1 port map( B1 => n148, B2 => n2145, C1 => n145, C2 => n2113
                           , A => n1054, ZN => n1047);
   U1079 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n142, B1 => 
                           REGISTERS_28_4_port, B2 => n139, ZN => n1054);
   U1080 : OAI221_X1 port map( B1 => n115, B2 => n1825, C1 => n112, C2 => n1793
                           , A => n1061, ZN => n1056);
   U1081 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n109, B1 => 
                           REGISTERS_10_4_port, B2 => n106, ZN => n1061);
   U1082 : OAI221_X1 port map( B1 => n127, B2 => n503, C1 => n124, C2 => n471, 
                           A => n1060, ZN => n1057);
   U1083 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n121, B1 => 
                           REGISTERS_6_4_port, B2 => n118, ZN => n1060);
   U1084 : OAI221_X1 port map( B1 => n103, B2 => n1889, C1 => n100, C2 => n1857
                           , A => n1062, ZN => n1055);
   U1085 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n97, B1 => 
                           REGISTERS_14_4_port, B2 => n94, ZN => n1062);
   U1086 : OAI221_X1 port map( B1 => n184, B2 => n1952, C1 => n181, C2 => n1920
                           , A => n1033, ZN => n1032);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_19_5_port, A2 => n178, B1 => 
                           REGISTERS_18_5_port, B2 => n175, ZN => n1033);
   U1088 : OAI221_X1 port map( B1 => n172, B2 => n2016, C1 => n169, C2 => n1984
                           , A => n1034, ZN => n1031);
   U1089 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n166, B1 => 
                           REGISTERS_22_5_port, B2 => n163, ZN => n1034);
   U1090 : OAI221_X1 port map( B1 => n160, B2 => n2080, C1 => n157, C2 => n2048
                           , A => n1035, ZN => n1030);
   U1091 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n154, B1 => 
                           REGISTERS_26_5_port, B2 => n151, ZN => n1035);
   U1092 : OAI221_X1 port map( B1 => n148, B2 => n2144, C1 => n145, C2 => n2112
                           , A => n1036, ZN => n1029);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n142, B1 => 
                           REGISTERS_28_5_port, B2 => n139, ZN => n1036);
   U1094 : OAI221_X1 port map( B1 => n115, B2 => n1824, C1 => n112, C2 => n1792
                           , A => n1043, ZN => n1038);
   U1095 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n109, B1 => 
                           REGISTERS_10_5_port, B2 => n106, ZN => n1043);
   U1096 : OAI221_X1 port map( B1 => n127, B2 => n502, C1 => n124, C2 => n470, 
                           A => n1042, ZN => n1039);
   U1097 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n121, B1 => 
                           REGISTERS_6_5_port, B2 => n118, ZN => n1042);
   U1098 : OAI221_X1 port map( B1 => n103, B2 => n1888, C1 => n100, C2 => n1856
                           , A => n1044, ZN => n1037);
   U1099 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n97, B1 => 
                           REGISTERS_14_5_port, B2 => n94, ZN => n1044);
   U1100 : OAI221_X1 port map( B1 => n184, B2 => n1951, C1 => n181, C2 => n1919
                           , A => n1015, ZN => n1014);
   U1101 : AOI22_X1 port map( A1 => REGISTERS_19_6_port, A2 => n178, B1 => 
                           REGISTERS_18_6_port, B2 => n175, ZN => n1015);
   U1102 : OAI221_X1 port map( B1 => n172, B2 => n2015, C1 => n169, C2 => n1983
                           , A => n1016, ZN => n1013);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n166, B1 => 
                           REGISTERS_22_6_port, B2 => n163, ZN => n1016);
   U1104 : OAI221_X1 port map( B1 => n160, B2 => n2079, C1 => n157, C2 => n2047
                           , A => n1017, ZN => n1012);
   U1105 : AOI22_X1 port map( A1 => REGISTERS_27_6_port, A2 => n154, B1 => 
                           REGISTERS_26_6_port, B2 => n151, ZN => n1017);
   U1106 : OAI221_X1 port map( B1 => n148, B2 => n2143, C1 => n145, C2 => n2111
                           , A => n1018, ZN => n1011);
   U1107 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n142, B1 => 
                           REGISTERS_28_6_port, B2 => n139, ZN => n1018);
   U1108 : OAI221_X1 port map( B1 => n115, B2 => n1823, C1 => n112, C2 => n1791
                           , A => n1025, ZN => n1020);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n109, B1 => 
                           REGISTERS_10_6_port, B2 => n106, ZN => n1025);
   U1110 : OAI221_X1 port map( B1 => n127, B2 => n501, C1 => n124, C2 => n469, 
                           A => n1024, ZN => n1021);
   U1111 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n121, B1 => 
                           REGISTERS_6_6_port, B2 => n118, ZN => n1024);
   U1112 : OAI221_X1 port map( B1 => n103, B2 => n1887, C1 => n100, C2 => n1855
                           , A => n1026, ZN => n1019);
   U1113 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n97, B1 => 
                           REGISTERS_14_6_port, B2 => n94, ZN => n1026);
   U1114 : OAI221_X1 port map( B1 => n184, B2 => n1950, C1 => n181, C2 => n1918
                           , A => n997, ZN => n996);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_19_7_port, A2 => n178, B1 => 
                           REGISTERS_18_7_port, B2 => n175, ZN => n997);
   U1116 : OAI221_X1 port map( B1 => n172, B2 => n2014, C1 => n169, C2 => n1982
                           , A => n998, ZN => n995);
   U1117 : AOI22_X1 port map( A1 => REGISTERS_23_7_port, A2 => n166, B1 => 
                           REGISTERS_22_7_port, B2 => n163, ZN => n998);
   U1118 : OAI221_X1 port map( B1 => n160, B2 => n2078, C1 => n157, C2 => n2046
                           , A => n999, ZN => n994);
   U1119 : AOI22_X1 port map( A1 => REGISTERS_27_7_port, A2 => n154, B1 => 
                           REGISTERS_26_7_port, B2 => n151, ZN => n999);
   U1120 : OAI221_X1 port map( B1 => n148, B2 => n2142, C1 => n145, C2 => n2110
                           , A => n1000, ZN => n993);
   U1121 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n142, B1 => 
                           REGISTERS_28_7_port, B2 => n139, ZN => n1000);
   U1122 : OAI221_X1 port map( B1 => n115, B2 => n1822, C1 => n112, C2 => n1790
                           , A => n1007, ZN => n1002);
   U1123 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n109, B1 => 
                           REGISTERS_10_7_port, B2 => n106, ZN => n1007);
   U1124 : OAI221_X1 port map( B1 => n127, B2 => n500, C1 => n124, C2 => n468, 
                           A => n1006, ZN => n1003);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n121, B1 => 
                           REGISTERS_6_7_port, B2 => n118, ZN => n1006);
   U1126 : OAI221_X1 port map( B1 => n103, B2 => n1886, C1 => n100, C2 => n1854
                           , A => n1008, ZN => n1001);
   U1127 : AOI22_X1 port map( A1 => REGISTERS_15_7_port, A2 => n97, B1 => 
                           REGISTERS_14_7_port, B2 => n94, ZN => n1008);
   U1128 : OAI221_X1 port map( B1 => n184, B2 => n1949, C1 => n181, C2 => n1917
                           , A => n979, ZN => n978);
   U1129 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n178, B1 => 
                           REGISTERS_18_8_port, B2 => n175, ZN => n979);
   U1130 : OAI221_X1 port map( B1 => n172, B2 => n2013, C1 => n169, C2 => n1981
                           , A => n980, ZN => n977);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n166, B1 => 
                           REGISTERS_22_8_port, B2 => n163, ZN => n980);
   U1132 : OAI221_X1 port map( B1 => n160, B2 => n2077, C1 => n157, C2 => n2045
                           , A => n981, ZN => n976);
   U1133 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n154, B1 => 
                           REGISTERS_26_8_port, B2 => n151, ZN => n981);
   U1134 : OAI221_X1 port map( B1 => n148, B2 => n2141, C1 => n145, C2 => n2109
                           , A => n982, ZN => n975);
   U1135 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n142, B1 => 
                           REGISTERS_28_8_port, B2 => n139, ZN => n982);
   U1136 : OAI221_X1 port map( B1 => n115, B2 => n1821, C1 => n112, C2 => n1789
                           , A => n989, ZN => n984);
   U1137 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n109, B1 => 
                           REGISTERS_10_8_port, B2 => n106, ZN => n989);
   U1138 : OAI221_X1 port map( B1 => n127, B2 => n499, C1 => n124, C2 => n467, 
                           A => n988, ZN => n985);
   U1139 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n121, B1 => 
                           REGISTERS_6_8_port, B2 => n118, ZN => n988);
   U1140 : OAI221_X1 port map( B1 => n103, B2 => n1885, C1 => n100, C2 => n1853
                           , A => n990, ZN => n983);
   U1141 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n97, B1 => 
                           REGISTERS_14_8_port, B2 => n94, ZN => n990);
   U1142 : OAI221_X1 port map( B1 => n184, B2 => n1948, C1 => n181, C2 => n1916
                           , A => n961, ZN => n960);
   U1143 : AOI22_X1 port map( A1 => REGISTERS_19_9_port, A2 => n178, B1 => 
                           REGISTERS_18_9_port, B2 => n175, ZN => n961);
   U1144 : OAI221_X1 port map( B1 => n172, B2 => n2012, C1 => n169, C2 => n1980
                           , A => n962, ZN => n959);
   U1145 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n166, B1 => 
                           REGISTERS_22_9_port, B2 => n163, ZN => n962);
   U1146 : OAI221_X1 port map( B1 => n160, B2 => n2076, C1 => n157, C2 => n2044
                           , A => n963, ZN => n958);
   U1147 : AOI22_X1 port map( A1 => REGISTERS_27_9_port, A2 => n154, B1 => 
                           REGISTERS_26_9_port, B2 => n151, ZN => n963);
   U1148 : OAI221_X1 port map( B1 => n148, B2 => n2140, C1 => n145, C2 => n2108
                           , A => n964, ZN => n957);
   U1149 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n142, B1 => 
                           REGISTERS_28_9_port, B2 => n139, ZN => n964);
   U1150 : OAI221_X1 port map( B1 => n115, B2 => n1820, C1 => n112, C2 => n1788
                           , A => n971, ZN => n966);
   U1151 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n109, B1 => 
                           REGISTERS_10_9_port, B2 => n106, ZN => n971);
   U1152 : OAI221_X1 port map( B1 => n127, B2 => n498, C1 => n124, C2 => n466, 
                           A => n970, ZN => n967);
   U1153 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n121, B1 => 
                           REGISTERS_6_9_port, B2 => n118, ZN => n970);
   U1154 : OAI221_X1 port map( B1 => n103, B2 => n1884, C1 => n100, C2 => n1852
                           , A => n972, ZN => n965);
   U1155 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n97, B1 => 
                           REGISTERS_14_9_port, B2 => n94, ZN => n972);
   U1156 : OAI221_X1 port map( B1 => n184, B2 => n1947, C1 => n181, C2 => n1915
                           , A => n943, ZN => n942);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n178, B1 => 
                           REGISTERS_18_10_port, B2 => n175, ZN => n943);
   U1158 : OAI221_X1 port map( B1 => n172, B2 => n2011, C1 => n169, C2 => n1979
                           , A => n944, ZN => n941);
   U1159 : AOI22_X1 port map( A1 => REGISTERS_23_10_port, A2 => n166, B1 => 
                           REGISTERS_22_10_port, B2 => n163, ZN => n944);
   U1160 : OAI221_X1 port map( B1 => n160, B2 => n2075, C1 => n157, C2 => n2043
                           , A => n945, ZN => n940);
   U1161 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n154, B1 => 
                           REGISTERS_26_10_port, B2 => n151, ZN => n945);
   U1162 : OAI221_X1 port map( B1 => n148, B2 => n2139, C1 => n145, C2 => n2107
                           , A => n946, ZN => n939);
   U1163 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n142, B1 => 
                           REGISTERS_28_10_port, B2 => n139, ZN => n946);
   U1164 : OAI221_X1 port map( B1 => n115, B2 => n1819, C1 => n112, C2 => n1787
                           , A => n953, ZN => n948);
   U1165 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n109, B1 => 
                           REGISTERS_10_10_port, B2 => n106, ZN => n953);
   U1166 : OAI221_X1 port map( B1 => n127, B2 => n497, C1 => n124, C2 => n465, 
                           A => n952, ZN => n949);
   U1167 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n121, B1 => 
                           REGISTERS_6_10_port, B2 => n118, ZN => n952);
   U1168 : OAI221_X1 port map( B1 => n103, B2 => n1883, C1 => n100, C2 => n1851
                           , A => n954, ZN => n947);
   U1169 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n97, B1 => 
                           REGISTERS_14_10_port, B2 => n94, ZN => n954);
   U1170 : OAI221_X1 port map( B1 => n184, B2 => n1946, C1 => n181, C2 => n1914
                           , A => n925, ZN => n924);
   U1171 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n178, B1 => 
                           REGISTERS_18_11_port, B2 => n175, ZN => n925);
   U1172 : OAI221_X1 port map( B1 => n172, B2 => n2010, C1 => n169, C2 => n1978
                           , A => n926, ZN => n923);
   U1173 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n166, B1 => 
                           REGISTERS_22_11_port, B2 => n163, ZN => n926);
   U1174 : OAI221_X1 port map( B1 => n160, B2 => n2074, C1 => n157, C2 => n2042
                           , A => n927, ZN => n922);
   U1175 : AOI22_X1 port map( A1 => REGISTERS_27_11_port, A2 => n154, B1 => 
                           REGISTERS_26_11_port, B2 => n151, ZN => n927);
   U1176 : OAI221_X1 port map( B1 => n148, B2 => n2138, C1 => n145, C2 => n2106
                           , A => n928, ZN => n921);
   U1177 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n142, B1 => 
                           REGISTERS_28_11_port, B2 => n139, ZN => n928);
   U1178 : OAI221_X1 port map( B1 => n115, B2 => n1818, C1 => n112, C2 => n1182
                           , A => n935, ZN => n930);
   U1179 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n109, B1 => 
                           REGISTERS_10_11_port, B2 => n106, ZN => n935);
   U1180 : OAI221_X1 port map( B1 => n127, B2 => n496, C1 => n124, C2 => n464, 
                           A => n934, ZN => n931);
   U1181 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n121, B1 => 
                           REGISTERS_6_11_port, B2 => n118, ZN => n934);
   U1182 : OAI221_X1 port map( B1 => n103, B2 => n1882, C1 => n100, C2 => n1850
                           , A => n936, ZN => n929);
   U1183 : AOI22_X1 port map( A1 => REGISTERS_15_11_port, A2 => n97, B1 => 
                           REGISTERS_14_11_port, B2 => n94, ZN => n936);
   U1184 : OAI221_X1 port map( B1 => n185, B2 => n1945, C1 => n182, C2 => n1913
                           , A => n907, ZN => n906);
   U1185 : AOI22_X1 port map( A1 => REGISTERS_19_12_port, A2 => n179, B1 => 
                           REGISTERS_18_12_port, B2 => n176, ZN => n907);
   U1186 : OAI221_X1 port map( B1 => n173, B2 => n2009, C1 => n170, C2 => n1977
                           , A => n908, ZN => n905);
   U1187 : AOI22_X1 port map( A1 => REGISTERS_23_12_port, A2 => n167, B1 => 
                           REGISTERS_22_12_port, B2 => n164, ZN => n908);
   U1188 : OAI221_X1 port map( B1 => n161, B2 => n2073, C1 => n158, C2 => n2041
                           , A => n909, ZN => n904);
   U1189 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n155, B1 => 
                           REGISTERS_26_12_port, B2 => n152, ZN => n909);
   U1190 : OAI221_X1 port map( B1 => n149, B2 => n2137, C1 => n146, C2 => n2105
                           , A => n910, ZN => n903);
   U1191 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n143, B1 => 
                           REGISTERS_28_12_port, B2 => n140, ZN => n910);
   U1192 : OAI221_X1 port map( B1 => n116, B2 => n1817, C1 => n113, C2 => n558,
                           A => n917, ZN => n912);
   U1193 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n110, B1 => 
                           REGISTERS_10_12_port, B2 => n107, ZN => n917);
   U1194 : OAI221_X1 port map( B1 => n128, B2 => n495, C1 => n125, C2 => n463, 
                           A => n916, ZN => n913);
   U1195 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n122, B1 => 
                           REGISTERS_6_12_port, B2 => n119, ZN => n916);
   U1196 : OAI221_X1 port map( B1 => n104, B2 => n1881, C1 => n101, C2 => n1849
                           , A => n918, ZN => n911);
   U1197 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n98, B1 => 
                           REGISTERS_14_12_port, B2 => n95, ZN => n918);
   U1198 : OAI221_X1 port map( B1 => n185, B2 => n1944, C1 => n182, C2 => n1912
                           , A => n889, ZN => n888);
   U1199 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n179, B1 => 
                           REGISTERS_18_13_port, B2 => n176, ZN => n889);
   U1200 : OAI221_X1 port map( B1 => n173, B2 => n2008, C1 => n170, C2 => n1976
                           , A => n890, ZN => n887);
   U1201 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n167, B1 => 
                           REGISTERS_22_13_port, B2 => n164, ZN => n890);
   U1202 : OAI221_X1 port map( B1 => n161, B2 => n2072, C1 => n158, C2 => n2040
                           , A => n891, ZN => n886);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_27_13_port, A2 => n155, B1 => 
                           REGISTERS_26_13_port, B2 => n152, ZN => n891);
   U1204 : OAI221_X1 port map( B1 => n149, B2 => n2136, C1 => n146, C2 => n2104
                           , A => n892, ZN => n885);
   U1205 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n143, B1 => 
                           REGISTERS_28_13_port, B2 => n140, ZN => n892);
   U1206 : OAI221_X1 port map( B1 => n116, B2 => n1816, C1 => n113, C2 => n526,
                           A => n899, ZN => n894);
   U1207 : AOI22_X1 port map( A1 => REGISTERS_11_13_port, A2 => n110, B1 => 
                           REGISTERS_10_13_port, B2 => n107, ZN => n899);
   U1208 : OAI221_X1 port map( B1 => n128, B2 => n494, C1 => n125, C2 => n462, 
                           A => n898, ZN => n895);
   U1209 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n122, B1 => 
                           REGISTERS_6_13_port, B2 => n119, ZN => n898);
   U1210 : OAI221_X1 port map( B1 => n104, B2 => n1880, C1 => n101, C2 => n1848
                           , A => n900, ZN => n893);
   U1211 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n98, B1 => 
                           REGISTERS_14_13_port, B2 => n95, ZN => n900);
   U1212 : OAI221_X1 port map( B1 => n185, B2 => n1943, C1 => n182, C2 => n1911
                           , A => n871, ZN => n870);
   U1213 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n179, B1 => 
                           REGISTERS_18_14_port, B2 => n176, ZN => n871);
   U1214 : OAI221_X1 port map( B1 => n173, B2 => n2007, C1 => n170, C2 => n1975
                           , A => n872, ZN => n869);
   U1215 : AOI22_X1 port map( A1 => REGISTERS_23_14_port, A2 => n167, B1 => 
                           REGISTERS_22_14_port, B2 => n164, ZN => n872);
   U1216 : OAI221_X1 port map( B1 => n161, B2 => n2071, C1 => n158, C2 => n2039
                           , A => n873, ZN => n868);
   U1217 : AOI22_X1 port map( A1 => REGISTERS_27_14_port, A2 => n155, B1 => 
                           REGISTERS_26_14_port, B2 => n152, ZN => n873);
   U1218 : OAI221_X1 port map( B1 => n149, B2 => n2135, C1 => n146, C2 => n2103
                           , A => n874, ZN => n867);
   U1219 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n143, B1 => 
                           REGISTERS_28_14_port, B2 => n140, ZN => n874);
   U1220 : OAI221_X1 port map( B1 => n116, B2 => n1815, C1 => n113, C2 => n525,
                           A => n881, ZN => n876);
   U1221 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n110, B1 => 
                           REGISTERS_10_14_port, B2 => n107, ZN => n881);
   U1222 : OAI221_X1 port map( B1 => n128, B2 => n493, C1 => n125, C2 => n461, 
                           A => n880, ZN => n877);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n122, B1 => 
                           REGISTERS_6_14_port, B2 => n119, ZN => n880);
   U1224 : OAI221_X1 port map( B1 => n104, B2 => n1879, C1 => n101, C2 => n1847
                           , A => n882, ZN => n875);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_15_14_port, A2 => n98, B1 => 
                           REGISTERS_14_14_port, B2 => n95, ZN => n882);
   U1226 : OAI221_X1 port map( B1 => n185, B2 => n1942, C1 => n182, C2 => n1910
                           , A => n853, ZN => n852);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n179, B1 => 
                           REGISTERS_18_15_port, B2 => n176, ZN => n853);
   U1228 : OAI221_X1 port map( B1 => n173, B2 => n2006, C1 => n170, C2 => n1974
                           , A => n854, ZN => n851);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n167, B1 => 
                           REGISTERS_22_15_port, B2 => n164, ZN => n854);
   U1230 : OAI221_X1 port map( B1 => n161, B2 => n2070, C1 => n158, C2 => n2038
                           , A => n855, ZN => n850);
   U1231 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n155, B1 => 
                           REGISTERS_26_15_port, B2 => n152, ZN => n855);
   U1232 : OAI221_X1 port map( B1 => n149, B2 => n2134, C1 => n146, C2 => n2102
                           , A => n856, ZN => n849);
   U1233 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n143, B1 => 
                           REGISTERS_28_15_port, B2 => n140, ZN => n856);
   U1234 : OAI221_X1 port map( B1 => n116, B2 => n1814, C1 => n113, C2 => n524,
                           A => n863, ZN => n858);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n110, B1 => 
                           REGISTERS_10_15_port, B2 => n107, ZN => n863);
   U1236 : OAI221_X1 port map( B1 => n128, B2 => n492, C1 => n125, C2 => n460, 
                           A => n862, ZN => n859);
   U1237 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n122, B1 => 
                           REGISTERS_6_15_port, B2 => n119, ZN => n862);
   U1238 : OAI221_X1 port map( B1 => n104, B2 => n1878, C1 => n101, C2 => n1846
                           , A => n864, ZN => n857);
   U1239 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n98, B1 => 
                           REGISTERS_14_15_port, B2 => n95, ZN => n864);
   U1240 : OAI221_X1 port map( B1 => n185, B2 => n1941, C1 => n182, C2 => n1909
                           , A => n835, ZN => n834);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n179, B1 => 
                           REGISTERS_18_16_port, B2 => n176, ZN => n835);
   U1242 : OAI221_X1 port map( B1 => n173, B2 => n2005, C1 => n170, C2 => n1973
                           , A => n836, ZN => n833);
   U1243 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n167, B1 => 
                           REGISTERS_22_16_port, B2 => n164, ZN => n836);
   U1244 : OAI221_X1 port map( B1 => n161, B2 => n2069, C1 => n158, C2 => n2037
                           , A => n837, ZN => n832);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n155, B1 => 
                           REGISTERS_26_16_port, B2 => n152, ZN => n837);
   U1246 : OAI221_X1 port map( B1 => n149, B2 => n2133, C1 => n146, C2 => n2101
                           , A => n838, ZN => n831);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n143, B1 => 
                           REGISTERS_28_16_port, B2 => n140, ZN => n838);
   U1248 : OAI221_X1 port map( B1 => n116, B2 => n1813, C1 => n113, C2 => n523,
                           A => n845, ZN => n840);
   U1249 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n110, B1 => 
                           REGISTERS_10_16_port, B2 => n107, ZN => n845);
   U1250 : OAI221_X1 port map( B1 => n128, B2 => n491, C1 => n125, C2 => n459, 
                           A => n844, ZN => n841);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n122, B1 => 
                           REGISTERS_6_16_port, B2 => n119, ZN => n844);
   U1252 : OAI221_X1 port map( B1 => n104, B2 => n1877, C1 => n101, C2 => n1845
                           , A => n846, ZN => n839);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n98, B1 => 
                           REGISTERS_14_16_port, B2 => n95, ZN => n846);
   U1254 : OAI221_X1 port map( B1 => n185, B2 => n1940, C1 => n182, C2 => n1908
                           , A => n817, ZN => n816);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_19_17_port, A2 => n179, B1 => 
                           REGISTERS_18_17_port, B2 => n176, ZN => n817);
   U1256 : OAI221_X1 port map( B1 => n173, B2 => n2004, C1 => n170, C2 => n1972
                           , A => n818, ZN => n815);
   U1257 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n167, B1 => 
                           REGISTERS_22_17_port, B2 => n164, ZN => n818);
   U1258 : OAI221_X1 port map( B1 => n161, B2 => n2068, C1 => n158, C2 => n2036
                           , A => n819, ZN => n814);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_27_17_port, A2 => n155, B1 => 
                           REGISTERS_26_17_port, B2 => n152, ZN => n819);
   U1260 : OAI221_X1 port map( B1 => n149, B2 => n2132, C1 => n146, C2 => n2100
                           , A => n820, ZN => n813);
   U1261 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n143, B1 => 
                           REGISTERS_28_17_port, B2 => n140, ZN => n820);
   U1262 : OAI221_X1 port map( B1 => n116, B2 => n1812, C1 => n113, C2 => n522,
                           A => n827, ZN => n822);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n110, B1 => 
                           REGISTERS_10_17_port, B2 => n107, ZN => n827);
   U1264 : OAI221_X1 port map( B1 => n128, B2 => n490, C1 => n125, C2 => n458, 
                           A => n826, ZN => n823);
   U1265 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n122, B1 => 
                           REGISTERS_6_17_port, B2 => n119, ZN => n826);
   U1266 : OAI221_X1 port map( B1 => n104, B2 => n1876, C1 => n101, C2 => n1844
                           , A => n828, ZN => n821);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n98, B1 => 
                           REGISTERS_14_17_port, B2 => n95, ZN => n828);
   U1268 : OAI221_X1 port map( B1 => n185, B2 => n1939, C1 => n182, C2 => n1907
                           , A => n799, ZN => n798);
   U1269 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n179, B1 => 
                           REGISTERS_18_18_port, B2 => n176, ZN => n799);
   U1270 : OAI221_X1 port map( B1 => n173, B2 => n2003, C1 => n170, C2 => n1971
                           , A => n800, ZN => n797);
   U1271 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n167, B1 => 
                           REGISTERS_22_18_port, B2 => n164, ZN => n800);
   U1272 : OAI221_X1 port map( B1 => n161, B2 => n2067, C1 => n158, C2 => n2035
                           , A => n801, ZN => n796);
   U1273 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n155, B1 => 
                           REGISTERS_26_18_port, B2 => n152, ZN => n801);
   U1274 : OAI221_X1 port map( B1 => n149, B2 => n2131, C1 => n146, C2 => n2099
                           , A => n802, ZN => n795);
   U1275 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n143, B1 => 
                           REGISTERS_28_18_port, B2 => n140, ZN => n802);
   U1276 : OAI221_X1 port map( B1 => n116, B2 => n1811, C1 => n113, C2 => n521,
                           A => n809, ZN => n804);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_11_18_port, A2 => n110, B1 => 
                           REGISTERS_10_18_port, B2 => n107, ZN => n809);
   U1278 : OAI221_X1 port map( B1 => n128, B2 => n489, C1 => n125, C2 => n457, 
                           A => n808, ZN => n805);
   U1279 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n122, B1 => 
                           REGISTERS_6_18_port, B2 => n119, ZN => n808);
   U1280 : OAI221_X1 port map( B1 => n104, B2 => n1875, C1 => n101, C2 => n1843
                           , A => n810, ZN => n803);
   U1281 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n98, B1 => 
                           REGISTERS_14_18_port, B2 => n95, ZN => n810);
   U1282 : OAI221_X1 port map( B1 => n185, B2 => n1938, C1 => n182, C2 => n1906
                           , A => n781, ZN => n780);
   U1283 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n179, B1 => 
                           REGISTERS_18_19_port, B2 => n176, ZN => n781);
   U1284 : OAI221_X1 port map( B1 => n173, B2 => n2002, C1 => n170, C2 => n1970
                           , A => n782, ZN => n779);
   U1285 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n167, B1 => 
                           REGISTERS_22_19_port, B2 => n164, ZN => n782);
   U1286 : OAI221_X1 port map( B1 => n161, B2 => n2066, C1 => n158, C2 => n2034
                           , A => n783, ZN => n778);
   U1287 : AOI22_X1 port map( A1 => REGISTERS_27_19_port, A2 => n155, B1 => 
                           REGISTERS_26_19_port, B2 => n152, ZN => n783);
   U1288 : OAI221_X1 port map( B1 => n149, B2 => n2130, C1 => n146, C2 => n2098
                           , A => n784, ZN => n777);
   U1289 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n143, B1 => 
                           REGISTERS_28_19_port, B2 => n140, ZN => n784);
   U1290 : OAI221_X1 port map( B1 => n116, B2 => n1810, C1 => n113, C2 => n520,
                           A => n791, ZN => n786);
   U1291 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n110, B1 => 
                           REGISTERS_10_19_port, B2 => n107, ZN => n791);
   U1292 : OAI221_X1 port map( B1 => n128, B2 => n488, C1 => n125, C2 => n456, 
                           A => n790, ZN => n787);
   U1293 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n122, B1 => 
                           REGISTERS_6_19_port, B2 => n119, ZN => n790);
   U1294 : OAI221_X1 port map( B1 => n104, B2 => n1874, C1 => n101, C2 => n1842
                           , A => n792, ZN => n785);
   U1295 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n98, B1 => 
                           REGISTERS_14_19_port, B2 => n95, ZN => n792);
   U1296 : OAI221_X1 port map( B1 => n185, B2 => n1937, C1 => n182, C2 => n1905
                           , A => n763, ZN => n762);
   U1297 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n179, B1 => 
                           REGISTERS_18_20_port, B2 => n176, ZN => n763);
   U1298 : OAI221_X1 port map( B1 => n173, B2 => n2001, C1 => n170, C2 => n1969
                           , A => n764, ZN => n761);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_23_20_port, A2 => n167, B1 => 
                           REGISTERS_22_20_port, B2 => n164, ZN => n764);
   U1300 : OAI221_X1 port map( B1 => n161, B2 => n2065, C1 => n158, C2 => n2033
                           , A => n765, ZN => n760);
   U1301 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n155, B1 => 
                           REGISTERS_26_20_port, B2 => n152, ZN => n765);
   U1302 : OAI221_X1 port map( B1 => n149, B2 => n2129, C1 => n146, C2 => n2097
                           , A => n766, ZN => n759);
   U1303 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n143, B1 => 
                           REGISTERS_28_20_port, B2 => n140, ZN => n766);
   U1304 : OAI221_X1 port map( B1 => n116, B2 => n1809, C1 => n113, C2 => n519,
                           A => n773, ZN => n768);
   U1305 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n110, B1 => 
                           REGISTERS_10_20_port, B2 => n107, ZN => n773);
   U1306 : OAI221_X1 port map( B1 => n128, B2 => n487, C1 => n125, C2 => n455, 
                           A => n772, ZN => n769);
   U1307 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n122, B1 => 
                           REGISTERS_6_20_port, B2 => n119, ZN => n772);
   U1308 : OAI221_X1 port map( B1 => n104, B2 => n1873, C1 => n101, C2 => n1841
                           , A => n774, ZN => n767);
   U1309 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n98, B1 => 
                           REGISTERS_14_20_port, B2 => n95, ZN => n774);
   U1310 : OAI221_X1 port map( B1 => n185, B2 => n1936, C1 => n182, C2 => n1904
                           , A => n745, ZN => n744);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n179, B1 => 
                           REGISTERS_18_21_port, B2 => n176, ZN => n745);
   U1312 : OAI221_X1 port map( B1 => n173, B2 => n2000, C1 => n170, C2 => n1968
                           , A => n746, ZN => n743);
   U1313 : AOI22_X1 port map( A1 => REGISTERS_23_21_port, A2 => n167, B1 => 
                           REGISTERS_22_21_port, B2 => n164, ZN => n746);
   U1314 : OAI221_X1 port map( B1 => n161, B2 => n2064, C1 => n158, C2 => n2032
                           , A => n747, ZN => n742);
   U1315 : AOI22_X1 port map( A1 => REGISTERS_27_21_port, A2 => n155, B1 => 
                           REGISTERS_26_21_port, B2 => n152, ZN => n747);
   U1316 : OAI221_X1 port map( B1 => n149, B2 => n2128, C1 => n146, C2 => n2096
                           , A => n748, ZN => n741);
   U1317 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n143, B1 => 
                           REGISTERS_28_21_port, B2 => n140, ZN => n748);
   U1318 : OAI221_X1 port map( B1 => n116, B2 => n1808, C1 => n113, C2 => n518,
                           A => n755, ZN => n750);
   U1319 : AOI22_X1 port map( A1 => REGISTERS_11_21_port, A2 => n110, B1 => 
                           REGISTERS_10_21_port, B2 => n107, ZN => n755);
   U1320 : OAI221_X1 port map( B1 => n128, B2 => n486, C1 => n125, C2 => n454, 
                           A => n754, ZN => n751);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n122, B1 => 
                           REGISTERS_6_21_port, B2 => n119, ZN => n754);
   U1322 : OAI221_X1 port map( B1 => n104, B2 => n1872, C1 => n101, C2 => n1840
                           , A => n756, ZN => n749);
   U1323 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n98, B1 => 
                           REGISTERS_14_21_port, B2 => n95, ZN => n756);
   U1324 : OAI221_X1 port map( B1 => n185, B2 => n1935, C1 => n182, C2 => n1903
                           , A => n727, ZN => n726);
   U1325 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n179, B1 => 
                           REGISTERS_18_22_port, B2 => n176, ZN => n727);
   U1326 : OAI221_X1 port map( B1 => n173, B2 => n1999, C1 => n170, C2 => n1967
                           , A => n728, ZN => n725);
   U1327 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n167, B1 => 
                           REGISTERS_22_22_port, B2 => n164, ZN => n728);
   U1328 : OAI221_X1 port map( B1 => n161, B2 => n2063, C1 => n158, C2 => n2031
                           , A => n729, ZN => n724);
   U1329 : AOI22_X1 port map( A1 => REGISTERS_27_22_port, A2 => n155, B1 => 
                           REGISTERS_26_22_port, B2 => n152, ZN => n729);
   U1330 : OAI221_X1 port map( B1 => n149, B2 => n2127, C1 => n146, C2 => n2095
                           , A => n730, ZN => n723);
   U1331 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n143, B1 => 
                           REGISTERS_28_22_port, B2 => n140, ZN => n730);
   U1332 : OAI221_X1 port map( B1 => n116, B2 => n1807, C1 => n113, C2 => n517,
                           A => n737, ZN => n732);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n110, B1 => 
                           REGISTERS_10_22_port, B2 => n107, ZN => n737);
   U1334 : OAI221_X1 port map( B1 => n128, B2 => n485, C1 => n125, C2 => n453, 
                           A => n736, ZN => n733);
   U1335 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n122, B1 => 
                           REGISTERS_6_22_port, B2 => n119, ZN => n736);
   U1336 : OAI221_X1 port map( B1 => n104, B2 => n1871, C1 => n101, C2 => n1839
                           , A => n738, ZN => n731);
   U1337 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n98, B1 => 
                           REGISTERS_14_22_port, B2 => n95, ZN => n738);
   U1338 : OAI221_X1 port map( B1 => n185, B2 => n1934, C1 => n182, C2 => n1902
                           , A => n709, ZN => n708);
   U1339 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n179, B1 => 
                           REGISTERS_18_23_port, B2 => n176, ZN => n709);
   U1340 : OAI221_X1 port map( B1 => n173, B2 => n1998, C1 => n170, C2 => n1966
                           , A => n710, ZN => n707);
   U1341 : AOI22_X1 port map( A1 => REGISTERS_23_23_port, A2 => n167, B1 => 
                           REGISTERS_22_23_port, B2 => n164, ZN => n710);
   U1342 : OAI221_X1 port map( B1 => n161, B2 => n2062, C1 => n158, C2 => n2030
                           , A => n711, ZN => n706);
   U1343 : AOI22_X1 port map( A1 => REGISTERS_27_23_port, A2 => n155, B1 => 
                           REGISTERS_26_23_port, B2 => n152, ZN => n711);
   U1344 : OAI221_X1 port map( B1 => n149, B2 => n2126, C1 => n146, C2 => n2094
                           , A => n712, ZN => n705);
   U1345 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n143, B1 => 
                           REGISTERS_28_23_port, B2 => n140, ZN => n712);
   U1346 : OAI221_X1 port map( B1 => n116, B2 => n1806, C1 => n113, C2 => n516,
                           A => n719, ZN => n714);
   U1347 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n110, B1 => 
                           REGISTERS_10_23_port, B2 => n107, ZN => n719);
   U1348 : OAI221_X1 port map( B1 => n128, B2 => n484, C1 => n125, C2 => n452, 
                           A => n718, ZN => n715);
   U1349 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n122, B1 => 
                           REGISTERS_6_23_port, B2 => n119, ZN => n718);
   U1350 : OAI221_X1 port map( B1 => n104, B2 => n1870, C1 => n101, C2 => n1838
                           , A => n720, ZN => n713);
   U1351 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n98, B1 => 
                           REGISTERS_14_23_port, B2 => n95, ZN => n720);
   U1352 : OAI221_X1 port map( B1 => n1957, B2 => n91, C1 => n1925, C2 => n88, 
                           A => n1747, ZN => n1746);
   U1353 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_0_port, B1 => n84, 
                           B2 => REGISTERS_18_0_port, ZN => n1747);
   U1354 : OAI221_X1 port map( B1 => n2021, B2 => n79, C1 => n1989, C2 => n76, 
                           A => n1752, ZN => n1745);
   U1355 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_0_port, B1 => n72, 
                           B2 => REGISTERS_22_0_port, ZN => n1752);
   U1356 : OAI221_X1 port map( B1 => n2085, B2 => n67, C1 => n2053, C2 => n64, 
                           A => n1756, ZN => n1744);
   U1357 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_0_port, B1 => n60, 
                           B2 => REGISTERS_26_0_port, ZN => n1756);
   U1358 : OAI221_X1 port map( B1 => n2149, B2 => n55, C1 => n2117, C2 => n52, 
                           A => n1759, ZN => n1743);
   U1359 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_0_port, B1 => n48, 
                           B2 => REGISTERS_28_0_port, ZN => n1759);
   U1360 : OAI221_X1 port map( B1 => n507, B2 => n34, C1 => n475, C2 => n31, A 
                           => n1768, ZN => n1763);
   U1361 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_0_port, B1 => n27, 
                           B2 => REGISTERS_6_0_port, ZN => n1768);
   U1362 : OAI221_X1 port map( B1 => n1829, B2 => n22, C1 => n1797, C2 => n19, 
                           A => n1770, ZN => n1762);
   U1363 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_0_port, B1 => n15, 
                           B2 => REGISTERS_10_0_port, ZN => n1770);
   U1364 : OAI221_X1 port map( B1 => n1956, B2 => n91, C1 => n1924, C2 => n88, 
                           A => n1729, ZN => n1728);
   U1365 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_1_port, B1 => n84, 
                           B2 => REGISTERS_18_1_port, ZN => n1729);
   U1366 : OAI221_X1 port map( B1 => n2020, B2 => n79, C1 => n1988, C2 => n76, 
                           A => n1730, ZN => n1727);
   U1367 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_1_port, B1 => n72, 
                           B2 => REGISTERS_22_1_port, ZN => n1730);
   U1368 : OAI221_X1 port map( B1 => n2084, B2 => n67, C1 => n2052, C2 => n64, 
                           A => n1731, ZN => n1726);
   U1369 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_1_port, B1 => n60, 
                           B2 => REGISTERS_26_1_port, ZN => n1731);
   U1370 : OAI221_X1 port map( B1 => n2148, B2 => n55, C1 => n2116, C2 => n52, 
                           A => n1732, ZN => n1725);
   U1371 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_1_port, B1 => n48, 
                           B2 => REGISTERS_28_1_port, ZN => n1732);
   U1372 : OAI221_X1 port map( B1 => n506, B2 => n34, C1 => n474, C2 => n31, A 
                           => n1738, ZN => n1735);
   U1373 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_1_port, B1 => n27, 
                           B2 => REGISTERS_6_1_port, ZN => n1738);
   U1374 : OAI221_X1 port map( B1 => n1828, B2 => n22, C1 => n1796, C2 => n19, 
                           A => n1739, ZN => n1734);
   U1375 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_1_port, B1 => n15, 
                           B2 => REGISTERS_10_1_port, ZN => n1739);
   U1376 : OAI221_X1 port map( B1 => n1955, B2 => n91, C1 => n1923, C2 => n88, 
                           A => n1711, ZN => n1710);
   U1377 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_2_port, B1 => n84, 
                           B2 => REGISTERS_18_2_port, ZN => n1711);
   U1378 : OAI221_X1 port map( B1 => n2019, B2 => n79, C1 => n1987, C2 => n76, 
                           A => n1712, ZN => n1709);
   U1379 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_2_port, B1 => n72, 
                           B2 => REGISTERS_22_2_port, ZN => n1712);
   U1380 : OAI221_X1 port map( B1 => n2083, B2 => n67, C1 => n2051, C2 => n64, 
                           A => n1713, ZN => n1708);
   U1381 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_2_port, B1 => n60, 
                           B2 => REGISTERS_26_2_port, ZN => n1713);
   U1382 : OAI221_X1 port map( B1 => n2147, B2 => n55, C1 => n2115, C2 => n52, 
                           A => n1714, ZN => n1707);
   U1383 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_2_port, B1 => n48, 
                           B2 => REGISTERS_28_2_port, ZN => n1714);
   U1384 : OAI221_X1 port map( B1 => n505, B2 => n34, C1 => n473, C2 => n31, A 
                           => n1720, ZN => n1717);
   U1385 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_2_port, B1 => n27, 
                           B2 => REGISTERS_6_2_port, ZN => n1720);
   U1386 : OAI221_X1 port map( B1 => n1827, B2 => n22, C1 => n1795, C2 => n19, 
                           A => n1721, ZN => n1716);
   U1387 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_2_port, B1 => n15, 
                           B2 => REGISTERS_10_2_port, ZN => n1721);
   U1388 : OAI221_X1 port map( B1 => n1954, B2 => n91, C1 => n1922, C2 => n88, 
                           A => n1693, ZN => n1692);
   U1389 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_3_port, B1 => n84, 
                           B2 => REGISTERS_18_3_port, ZN => n1693);
   U1390 : OAI221_X1 port map( B1 => n2018, B2 => n79, C1 => n1986, C2 => n76, 
                           A => n1694, ZN => n1691);
   U1391 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_3_port, B1 => n72, 
                           B2 => REGISTERS_22_3_port, ZN => n1694);
   U1392 : OAI221_X1 port map( B1 => n2082, B2 => n67, C1 => n2050, C2 => n64, 
                           A => n1695, ZN => n1690);
   U1393 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_3_port, B1 => n60, 
                           B2 => REGISTERS_26_3_port, ZN => n1695);
   U1394 : OAI221_X1 port map( B1 => n2146, B2 => n55, C1 => n2114, C2 => n52, 
                           A => n1696, ZN => n1689);
   U1395 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_3_port, B1 => n48, 
                           B2 => REGISTERS_28_3_port, ZN => n1696);
   U1396 : OAI221_X1 port map( B1 => n504, B2 => n34, C1 => n472, C2 => n31, A 
                           => n1702, ZN => n1699);
   U1397 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_3_port, B1 => n27, 
                           B2 => REGISTERS_6_3_port, ZN => n1702);
   U1398 : OAI221_X1 port map( B1 => n1826, B2 => n22, C1 => n1794, C2 => n19, 
                           A => n1703, ZN => n1698);
   U1399 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_3_port, B1 => n15, 
                           B2 => REGISTERS_10_3_port, ZN => n1703);
   U1400 : OAI221_X1 port map( B1 => n1953, B2 => n91, C1 => n1921, C2 => n88, 
                           A => n1675, ZN => n1674);
   U1401 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_4_port, B1 => n84, 
                           B2 => REGISTERS_18_4_port, ZN => n1675);
   U1402 : OAI221_X1 port map( B1 => n2017, B2 => n79, C1 => n1985, C2 => n76, 
                           A => n1676, ZN => n1673);
   U1403 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_4_port, B1 => n72, 
                           B2 => REGISTERS_22_4_port, ZN => n1676);
   U1404 : OAI221_X1 port map( B1 => n2081, B2 => n67, C1 => n2049, C2 => n64, 
                           A => n1677, ZN => n1672);
   U1405 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_4_port, B1 => n60, 
                           B2 => REGISTERS_26_4_port, ZN => n1677);
   U1406 : OAI221_X1 port map( B1 => n2145, B2 => n55, C1 => n2113, C2 => n52, 
                           A => n1678, ZN => n1671);
   U1407 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_4_port, B1 => n48, 
                           B2 => REGISTERS_28_4_port, ZN => n1678);
   U1408 : OAI221_X1 port map( B1 => n503, B2 => n34, C1 => n471, C2 => n31, A 
                           => n1684, ZN => n1681);
   U1409 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_4_port, B1 => n27, 
                           B2 => REGISTERS_6_4_port, ZN => n1684);
   U1410 : OAI221_X1 port map( B1 => n1825, B2 => n22, C1 => n1793, C2 => n19, 
                           A => n1685, ZN => n1680);
   U1411 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_4_port, B1 => n15, 
                           B2 => REGISTERS_10_4_port, ZN => n1685);
   U1412 : OAI221_X1 port map( B1 => n1952, B2 => n91, C1 => n1920, C2 => n88, 
                           A => n1657, ZN => n1656);
   U1413 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_5_port, B1 => n84, 
                           B2 => REGISTERS_18_5_port, ZN => n1657);
   U1414 : OAI221_X1 port map( B1 => n2016, B2 => n79, C1 => n1984, C2 => n76, 
                           A => n1658, ZN => n1655);
   U1415 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_5_port, B1 => n72, 
                           B2 => REGISTERS_22_5_port, ZN => n1658);
   U1416 : OAI221_X1 port map( B1 => n2080, B2 => n67, C1 => n2048, C2 => n64, 
                           A => n1659, ZN => n1654);
   U1417 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_5_port, B1 => n60, 
                           B2 => REGISTERS_26_5_port, ZN => n1659);
   U1418 : OAI221_X1 port map( B1 => n2144, B2 => n55, C1 => n2112, C2 => n52, 
                           A => n1660, ZN => n1653);
   U1419 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_5_port, B1 => n48, 
                           B2 => REGISTERS_28_5_port, ZN => n1660);
   U1420 : OAI221_X1 port map( B1 => n502, B2 => n34, C1 => n470, C2 => n31, A 
                           => n1666, ZN => n1663);
   U1421 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_5_port, B1 => n27, 
                           B2 => REGISTERS_6_5_port, ZN => n1666);
   U1422 : OAI221_X1 port map( B1 => n1824, B2 => n22, C1 => n1792, C2 => n19, 
                           A => n1667, ZN => n1662);
   U1423 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_5_port, B1 => n15, 
                           B2 => REGISTERS_10_5_port, ZN => n1667);
   U1424 : OAI221_X1 port map( B1 => n1951, B2 => n91, C1 => n1919, C2 => n88, 
                           A => n1639, ZN => n1638);
   U1425 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_6_port, B1 => n84, 
                           B2 => REGISTERS_18_6_port, ZN => n1639);
   U1426 : OAI221_X1 port map( B1 => n2015, B2 => n79, C1 => n1983, C2 => n76, 
                           A => n1640, ZN => n1637);
   U1427 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_6_port, B1 => n72, 
                           B2 => REGISTERS_22_6_port, ZN => n1640);
   U1428 : OAI221_X1 port map( B1 => n2079, B2 => n67, C1 => n2047, C2 => n64, 
                           A => n1641, ZN => n1636);
   U1429 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_6_port, B1 => n60, 
                           B2 => REGISTERS_26_6_port, ZN => n1641);
   U1430 : OAI221_X1 port map( B1 => n2143, B2 => n55, C1 => n2111, C2 => n52, 
                           A => n1642, ZN => n1635);
   U1431 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_6_port, B1 => n48, 
                           B2 => REGISTERS_28_6_port, ZN => n1642);
   U1432 : OAI221_X1 port map( B1 => n501, B2 => n34, C1 => n469, C2 => n31, A 
                           => n1648, ZN => n1645);
   U1433 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_6_port, B1 => n27, 
                           B2 => REGISTERS_6_6_port, ZN => n1648);
   U1434 : OAI221_X1 port map( B1 => n1823, B2 => n22, C1 => n1791, C2 => n19, 
                           A => n1649, ZN => n1644);
   U1435 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_6_port, B1 => n15, 
                           B2 => REGISTERS_10_6_port, ZN => n1649);
   U1436 : OAI221_X1 port map( B1 => n1950, B2 => n91, C1 => n1918, C2 => n88, 
                           A => n1621, ZN => n1620);
   U1437 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_7_port, B1 => n84, 
                           B2 => REGISTERS_18_7_port, ZN => n1621);
   U1438 : OAI221_X1 port map( B1 => n2014, B2 => n79, C1 => n1982, C2 => n76, 
                           A => n1622, ZN => n1619);
   U1439 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_7_port, B1 => n72, 
                           B2 => REGISTERS_22_7_port, ZN => n1622);
   U1440 : OAI221_X1 port map( B1 => n2078, B2 => n67, C1 => n2046, C2 => n64, 
                           A => n1623, ZN => n1618);
   U1441 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_7_port, B1 => n60, 
                           B2 => REGISTERS_26_7_port, ZN => n1623);
   U1442 : OAI221_X1 port map( B1 => n2142, B2 => n55, C1 => n2110, C2 => n52, 
                           A => n1624, ZN => n1617);
   U1443 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_7_port, B1 => n48, 
                           B2 => REGISTERS_28_7_port, ZN => n1624);
   U1444 : OAI221_X1 port map( B1 => n500, B2 => n34, C1 => n468, C2 => n31, A 
                           => n1630, ZN => n1627);
   U1445 : AOI22_X1 port map( A1 => n28, A2 => REGISTERS_7_7_port, B1 => n27, 
                           B2 => REGISTERS_6_7_port, ZN => n1630);
   U1446 : OAI221_X1 port map( B1 => n1822, B2 => n22, C1 => n1790, C2 => n19, 
                           A => n1631, ZN => n1626);
   U1447 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_7_port, B1 => n15, 
                           B2 => REGISTERS_10_7_port, ZN => n1631);
   U1448 : OAI221_X1 port map( B1 => n1949, B2 => n91, C1 => n1917, C2 => n88, 
                           A => n1603, ZN => n1602);
   U1449 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_8_port, B1 => n83, 
                           B2 => REGISTERS_18_8_port, ZN => n1603);
   U1450 : OAI221_X1 port map( B1 => n2013, B2 => n79, C1 => n1981, C2 => n76, 
                           A => n1604, ZN => n1601);
   U1451 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_8_port, B1 => n71, 
                           B2 => REGISTERS_22_8_port, ZN => n1604);
   U1452 : OAI221_X1 port map( B1 => n2077, B2 => n67, C1 => n2045, C2 => n64, 
                           A => n1605, ZN => n1600);
   U1453 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_8_port, B1 => n59, 
                           B2 => REGISTERS_26_8_port, ZN => n1605);
   U1454 : OAI221_X1 port map( B1 => n2141, B2 => n55, C1 => n2109, C2 => n52, 
                           A => n1606, ZN => n1599);
   U1455 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_8_port, B1 => n47, 
                           B2 => REGISTERS_28_8_port, ZN => n1606);
   U1456 : OAI221_X1 port map( B1 => n1821, B2 => n22, C1 => n1789, C2 => n19, 
                           A => n1613, ZN => n1608);
   U1457 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_8_port, B1 => n14, 
                           B2 => REGISTERS_10_8_port, ZN => n1613);
   U1458 : OAI221_X1 port map( B1 => n1948, B2 => n91, C1 => n1916, C2 => n88, 
                           A => n1585, ZN => n1584);
   U1459 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_9_port, B1 => n83, 
                           B2 => REGISTERS_18_9_port, ZN => n1585);
   U1460 : OAI221_X1 port map( B1 => n2012, B2 => n79, C1 => n1980, C2 => n76, 
                           A => n1586, ZN => n1583);
   U1461 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_9_port, B1 => n71, 
                           B2 => REGISTERS_22_9_port, ZN => n1586);
   U1462 : OAI221_X1 port map( B1 => n2076, B2 => n67, C1 => n2044, C2 => n64, 
                           A => n1587, ZN => n1582);
   U1463 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_9_port, B1 => n59, 
                           B2 => REGISTERS_26_9_port, ZN => n1587);
   U1464 : OAI221_X1 port map( B1 => n2140, B2 => n55, C1 => n2108, C2 => n52, 
                           A => n1588, ZN => n1581);
   U1465 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_9_port, B1 => n47, 
                           B2 => REGISTERS_28_9_port, ZN => n1588);
   U1466 : OAI221_X1 port map( B1 => n1820, B2 => n22, C1 => n1788, C2 => n19, 
                           A => n1595, ZN => n1590);
   U1467 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_9_port, B1 => n14, 
                           B2 => REGISTERS_10_9_port, ZN => n1595);
   U1468 : OAI221_X1 port map( B1 => n1947, B2 => n91, C1 => n1915, C2 => n88, 
                           A => n1567, ZN => n1566);
   U1469 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_10_port, B1 => n83,
                           B2 => REGISTERS_18_10_port, ZN => n1567);
   U1470 : OAI221_X1 port map( B1 => n2011, B2 => n79, C1 => n1979, C2 => n76, 
                           A => n1568, ZN => n1565);
   U1471 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_10_port, B1 => n71,
                           B2 => REGISTERS_22_10_port, ZN => n1568);
   U1472 : OAI221_X1 port map( B1 => n2075, B2 => n67, C1 => n2043, C2 => n64, 
                           A => n1569, ZN => n1564);
   U1473 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_10_port, B1 => n59,
                           B2 => REGISTERS_26_10_port, ZN => n1569);
   U1474 : OAI221_X1 port map( B1 => n2139, B2 => n55, C1 => n2107, C2 => n52, 
                           A => n1570, ZN => n1563);
   U1475 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_10_port, B1 => n47,
                           B2 => REGISTERS_28_10_port, ZN => n1570);
   U1476 : OAI221_X1 port map( B1 => n1819, B2 => n22, C1 => n1787, C2 => n19, 
                           A => n1577, ZN => n1572);
   U1477 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_10_port, B1 => n14,
                           B2 => REGISTERS_10_10_port, ZN => n1577);
   U1478 : OAI221_X1 port map( B1 => n1946, B2 => n91, C1 => n1914, C2 => n88, 
                           A => n1549, ZN => n1548);
   U1479 : AOI22_X1 port map( A1 => n85, A2 => REGISTERS_19_11_port, B1 => n83,
                           B2 => REGISTERS_18_11_port, ZN => n1549);
   U1480 : OAI221_X1 port map( B1 => n2010, B2 => n79, C1 => n1978, C2 => n76, 
                           A => n1550, ZN => n1547);
   U1481 : AOI22_X1 port map( A1 => n73, A2 => REGISTERS_23_11_port, B1 => n71,
                           B2 => REGISTERS_22_11_port, ZN => n1550);
   U1482 : OAI221_X1 port map( B1 => n2074, B2 => n67, C1 => n2042, C2 => n64, 
                           A => n1551, ZN => n1546);
   U1483 : AOI22_X1 port map( A1 => n61, A2 => REGISTERS_27_11_port, B1 => n59,
                           B2 => REGISTERS_26_11_port, ZN => n1551);
   U1484 : OAI221_X1 port map( B1 => n2138, B2 => n55, C1 => n2106, C2 => n52, 
                           A => n1552, ZN => n1545);
   U1485 : AOI22_X1 port map( A1 => n49, A2 => REGISTERS_29_11_port, B1 => n47,
                           B2 => REGISTERS_28_11_port, ZN => n1552);
   U1486 : OAI221_X1 port map( B1 => n1818, B2 => n22, C1 => n1182, C2 => n19, 
                           A => n1559, ZN => n1554);
   U1487 : AOI22_X1 port map( A1 => n16, A2 => REGISTERS_11_11_port, B1 => n14,
                           B2 => REGISTERS_10_11_port, ZN => n1559);
   U1488 : OAI221_X1 port map( B1 => n1945, B2 => n92, C1 => n1913, C2 => n89, 
                           A => n1531, ZN => n1530);
   U1489 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_12_port, B1 => n83,
                           B2 => REGISTERS_18_12_port, ZN => n1531);
   U1490 : OAI221_X1 port map( B1 => n2009, B2 => n80, C1 => n1977, C2 => n77, 
                           A => n1532, ZN => n1529);
   U1491 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_12_port, B1 => n71,
                           B2 => REGISTERS_22_12_port, ZN => n1532);
   U1492 : OAI221_X1 port map( B1 => n2073, B2 => n68, C1 => n2041, C2 => n65, 
                           A => n1533, ZN => n1528);
   U1493 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_12_port, B1 => n59,
                           B2 => REGISTERS_26_12_port, ZN => n1533);
   U1494 : OAI221_X1 port map( B1 => n2137, B2 => n56, C1 => n2105, C2 => n53, 
                           A => n1534, ZN => n1527);
   U1495 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_12_port, B1 => n47,
                           B2 => REGISTERS_28_12_port, ZN => n1534);
   U1496 : OAI221_X1 port map( B1 => n1817, B2 => n23, C1 => n558, C2 => n20, A
                           => n1541, ZN => n1536);
   U1497 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_12_port, B1 => n14,
                           B2 => REGISTERS_10_12_port, ZN => n1541);
   U1498 : OAI221_X1 port map( B1 => n1944, B2 => n92, C1 => n1912, C2 => n89, 
                           A => n1513, ZN => n1512);
   U1499 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_13_port, B1 => n83,
                           B2 => REGISTERS_18_13_port, ZN => n1513);
   U1500 : OAI221_X1 port map( B1 => n2008, B2 => n80, C1 => n1976, C2 => n77, 
                           A => n1514, ZN => n1511);
   U1501 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_13_port, B1 => n71,
                           B2 => REGISTERS_22_13_port, ZN => n1514);
   U1502 : OAI221_X1 port map( B1 => n2072, B2 => n68, C1 => n2040, C2 => n65, 
                           A => n1515, ZN => n1510);
   U1503 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_13_port, B1 => n59,
                           B2 => REGISTERS_26_13_port, ZN => n1515);
   U1504 : OAI221_X1 port map( B1 => n2136, B2 => n56, C1 => n2104, C2 => n53, 
                           A => n1516, ZN => n1509);
   U1505 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_13_port, B1 => n47,
                           B2 => REGISTERS_28_13_port, ZN => n1516);
   U1506 : OAI221_X1 port map( B1 => n1816, B2 => n23, C1 => n526, C2 => n20, A
                           => n1523, ZN => n1518);
   U1507 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_13_port, B1 => n14,
                           B2 => REGISTERS_10_13_port, ZN => n1523);
   U1508 : OAI221_X1 port map( B1 => n1943, B2 => n92, C1 => n1911, C2 => n89, 
                           A => n1495, ZN => n1494);
   U1509 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_14_port, B1 => n83,
                           B2 => REGISTERS_18_14_port, ZN => n1495);
   U1510 : OAI221_X1 port map( B1 => n2007, B2 => n80, C1 => n1975, C2 => n77, 
                           A => n1496, ZN => n1493);
   U1511 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_14_port, B1 => n71,
                           B2 => REGISTERS_22_14_port, ZN => n1496);
   U1512 : OAI221_X1 port map( B1 => n2071, B2 => n68, C1 => n2039, C2 => n65, 
                           A => n1497, ZN => n1492);
   U1513 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_14_port, B1 => n59,
                           B2 => REGISTERS_26_14_port, ZN => n1497);
   U1514 : OAI221_X1 port map( B1 => n2135, B2 => n56, C1 => n2103, C2 => n53, 
                           A => n1498, ZN => n1491);
   U1515 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_14_port, B1 => n47,
                           B2 => REGISTERS_28_14_port, ZN => n1498);
   U1516 : OAI221_X1 port map( B1 => n1815, B2 => n23, C1 => n525, C2 => n20, A
                           => n1505, ZN => n1500);
   U1517 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_14_port, B1 => n14,
                           B2 => REGISTERS_10_14_port, ZN => n1505);
   U1518 : OAI221_X1 port map( B1 => n1942, B2 => n92, C1 => n1910, C2 => n89, 
                           A => n1477, ZN => n1476);
   U1519 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_15_port, B1 => n83,
                           B2 => REGISTERS_18_15_port, ZN => n1477);
   U1520 : OAI221_X1 port map( B1 => n2006, B2 => n80, C1 => n1974, C2 => n77, 
                           A => n1478, ZN => n1475);
   U1521 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_15_port, B1 => n71,
                           B2 => REGISTERS_22_15_port, ZN => n1478);
   U1522 : OAI221_X1 port map( B1 => n2070, B2 => n68, C1 => n2038, C2 => n65, 
                           A => n1479, ZN => n1474);
   U1523 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_15_port, B1 => n59,
                           B2 => REGISTERS_26_15_port, ZN => n1479);
   U1524 : OAI221_X1 port map( B1 => n2134, B2 => n56, C1 => n2102, C2 => n53, 
                           A => n1480, ZN => n1473);
   U1525 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_15_port, B1 => n47,
                           B2 => REGISTERS_28_15_port, ZN => n1480);
   U1526 : OAI221_X1 port map( B1 => n1814, B2 => n23, C1 => n524, C2 => n20, A
                           => n1487, ZN => n1482);
   U1527 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_15_port, B1 => n14,
                           B2 => REGISTERS_10_15_port, ZN => n1487);
   U1528 : OAI221_X1 port map( B1 => n1941, B2 => n92, C1 => n1909, C2 => n89, 
                           A => n1459, ZN => n1458);
   U1529 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_16_port, B1 => n83,
                           B2 => REGISTERS_18_16_port, ZN => n1459);
   U1530 : OAI221_X1 port map( B1 => n2005, B2 => n80, C1 => n1973, C2 => n77, 
                           A => n1460, ZN => n1457);
   U1531 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_16_port, B1 => n71,
                           B2 => REGISTERS_22_16_port, ZN => n1460);
   U1532 : OAI221_X1 port map( B1 => n2069, B2 => n68, C1 => n2037, C2 => n65, 
                           A => n1461, ZN => n1456);
   U1533 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_16_port, B1 => n59,
                           B2 => REGISTERS_26_16_port, ZN => n1461);
   U1534 : OAI221_X1 port map( B1 => n2133, B2 => n56, C1 => n2101, C2 => n53, 
                           A => n1462, ZN => n1455);
   U1535 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_16_port, B1 => n47,
                           B2 => REGISTERS_28_16_port, ZN => n1462);
   U1536 : OAI221_X1 port map( B1 => n1813, B2 => n23, C1 => n523, C2 => n20, A
                           => n1469, ZN => n1464);
   U1537 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_16_port, B1 => n14,
                           B2 => REGISTERS_10_16_port, ZN => n1469);
   U1538 : OAI221_X1 port map( B1 => n1940, B2 => n92, C1 => n1908, C2 => n89, 
                           A => n1441, ZN => n1440);
   U1539 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_17_port, B1 => n83,
                           B2 => REGISTERS_18_17_port, ZN => n1441);
   U1540 : OAI221_X1 port map( B1 => n2004, B2 => n80, C1 => n1972, C2 => n77, 
                           A => n1442, ZN => n1439);
   U1541 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_17_port, B1 => n71,
                           B2 => REGISTERS_22_17_port, ZN => n1442);
   U1542 : OAI221_X1 port map( B1 => n2068, B2 => n68, C1 => n2036, C2 => n65, 
                           A => n1443, ZN => n1438);
   U1543 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_17_port, B1 => n59,
                           B2 => REGISTERS_26_17_port, ZN => n1443);
   U1544 : OAI221_X1 port map( B1 => n2132, B2 => n56, C1 => n2100, C2 => n53, 
                           A => n1444, ZN => n1437);
   U1545 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_17_port, B1 => n47,
                           B2 => REGISTERS_28_17_port, ZN => n1444);
   U1546 : OAI221_X1 port map( B1 => n1812, B2 => n23, C1 => n522, C2 => n20, A
                           => n1451, ZN => n1446);
   U1547 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_17_port, B1 => n14,
                           B2 => REGISTERS_10_17_port, ZN => n1451);
   U1548 : OAI221_X1 port map( B1 => n1939, B2 => n92, C1 => n1907, C2 => n89, 
                           A => n1423, ZN => n1422);
   U1549 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_18_port, B1 => n83,
                           B2 => REGISTERS_18_18_port, ZN => n1423);
   U1550 : OAI221_X1 port map( B1 => n2003, B2 => n80, C1 => n1971, C2 => n77, 
                           A => n1424, ZN => n1421);
   U1551 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_18_port, B1 => n71,
                           B2 => REGISTERS_22_18_port, ZN => n1424);
   U1552 : OAI221_X1 port map( B1 => n2067, B2 => n68, C1 => n2035, C2 => n65, 
                           A => n1425, ZN => n1420);
   U1553 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_18_port, B1 => n59,
                           B2 => REGISTERS_26_18_port, ZN => n1425);
   U1554 : OAI221_X1 port map( B1 => n2131, B2 => n56, C1 => n2099, C2 => n53, 
                           A => n1426, ZN => n1419);
   U1555 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_18_port, B1 => n47,
                           B2 => REGISTERS_28_18_port, ZN => n1426);
   U1556 : OAI221_X1 port map( B1 => n1811, B2 => n23, C1 => n521, C2 => n20, A
                           => n1433, ZN => n1428);
   U1557 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_18_port, B1 => n14,
                           B2 => REGISTERS_10_18_port, ZN => n1433);
   U1558 : OAI221_X1 port map( B1 => n1938, B2 => n92, C1 => n1906, C2 => n89, 
                           A => n1405, ZN => n1404);
   U1559 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_19_port, B1 => n83,
                           B2 => REGISTERS_18_19_port, ZN => n1405);
   U1560 : OAI221_X1 port map( B1 => n2002, B2 => n80, C1 => n1970, C2 => n77, 
                           A => n1406, ZN => n1403);
   U1561 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_19_port, B1 => n71,
                           B2 => REGISTERS_22_19_port, ZN => n1406);
   U1562 : OAI221_X1 port map( B1 => n2066, B2 => n68, C1 => n2034, C2 => n65, 
                           A => n1407, ZN => n1402);
   U1563 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_19_port, B1 => n59,
                           B2 => REGISTERS_26_19_port, ZN => n1407);
   U1564 : OAI221_X1 port map( B1 => n2130, B2 => n56, C1 => n2098, C2 => n53, 
                           A => n1408, ZN => n1401);
   U1565 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_19_port, B1 => n47,
                           B2 => REGISTERS_28_19_port, ZN => n1408);
   U1566 : OAI221_X1 port map( B1 => n1810, B2 => n23, C1 => n520, C2 => n20, A
                           => n1415, ZN => n1410);
   U1567 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_19_port, B1 => n14,
                           B2 => REGISTERS_10_19_port, ZN => n1415);
   U1568 : OAI221_X1 port map( B1 => n1937, B2 => n92, C1 => n1905, C2 => n89, 
                           A => n1387, ZN => n1386);
   U1569 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_20_port, B1 => n82,
                           B2 => REGISTERS_18_20_port, ZN => n1387);
   U1570 : OAI221_X1 port map( B1 => n2001, B2 => n80, C1 => n1969, C2 => n77, 
                           A => n1388, ZN => n1385);
   U1571 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_20_port, B1 => n70,
                           B2 => REGISTERS_22_20_port, ZN => n1388);
   U1572 : OAI221_X1 port map( B1 => n2065, B2 => n68, C1 => n2033, C2 => n65, 
                           A => n1389, ZN => n1384);
   U1573 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_20_port, B1 => n58,
                           B2 => REGISTERS_26_20_port, ZN => n1389);
   U1574 : OAI221_X1 port map( B1 => n2129, B2 => n56, C1 => n2097, C2 => n53, 
                           A => n1390, ZN => n1383);
   U1575 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_20_port, B1 => n46,
                           B2 => REGISTERS_28_20_port, ZN => n1390);
   U1576 : OAI221_X1 port map( B1 => n1809, B2 => n23, C1 => n519, C2 => n20, A
                           => n1397, ZN => n1392);
   U1577 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_20_port, B1 => n13,
                           B2 => REGISTERS_10_20_port, ZN => n1397);
   U1578 : OAI221_X1 port map( B1 => n1936, B2 => n92, C1 => n1904, C2 => n89, 
                           A => n1369, ZN => n1368);
   U1579 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_21_port, B1 => n82,
                           B2 => REGISTERS_18_21_port, ZN => n1369);
   U1580 : OAI221_X1 port map( B1 => n2000, B2 => n80, C1 => n1968, C2 => n77, 
                           A => n1370, ZN => n1367);
   U1581 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_21_port, B1 => n70,
                           B2 => REGISTERS_22_21_port, ZN => n1370);
   U1582 : OAI221_X1 port map( B1 => n2064, B2 => n68, C1 => n2032, C2 => n65, 
                           A => n1371, ZN => n1366);
   U1583 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_21_port, B1 => n58,
                           B2 => REGISTERS_26_21_port, ZN => n1371);
   U1584 : OAI221_X1 port map( B1 => n2128, B2 => n56, C1 => n2096, C2 => n53, 
                           A => n1372, ZN => n1365);
   U1585 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_21_port, B1 => n46,
                           B2 => REGISTERS_28_21_port, ZN => n1372);
   U1586 : OAI221_X1 port map( B1 => n1808, B2 => n23, C1 => n518, C2 => n20, A
                           => n1379, ZN => n1374);
   U1587 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_21_port, B1 => n13,
                           B2 => REGISTERS_10_21_port, ZN => n1379);
   U1588 : OAI221_X1 port map( B1 => n1935, B2 => n92, C1 => n1903, C2 => n89, 
                           A => n1351, ZN => n1350);
   U1589 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_22_port, B1 => n82,
                           B2 => REGISTERS_18_22_port, ZN => n1351);
   U1590 : OAI221_X1 port map( B1 => n1999, B2 => n80, C1 => n1967, C2 => n77, 
                           A => n1352, ZN => n1349);
   U1591 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_22_port, B1 => n70,
                           B2 => REGISTERS_22_22_port, ZN => n1352);
   U1592 : OAI221_X1 port map( B1 => n2063, B2 => n68, C1 => n2031, C2 => n65, 
                           A => n1353, ZN => n1348);
   U1593 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_22_port, B1 => n58,
                           B2 => REGISTERS_26_22_port, ZN => n1353);
   U1594 : OAI221_X1 port map( B1 => n2127, B2 => n56, C1 => n2095, C2 => n53, 
                           A => n1354, ZN => n1347);
   U1595 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_22_port, B1 => n46,
                           B2 => REGISTERS_28_22_port, ZN => n1354);
   U1596 : OAI221_X1 port map( B1 => n1807, B2 => n23, C1 => n517, C2 => n20, A
                           => n1361, ZN => n1356);
   U1597 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_22_port, B1 => n13,
                           B2 => REGISTERS_10_22_port, ZN => n1361);
   U1598 : OAI221_X1 port map( B1 => n1934, B2 => n92, C1 => n1902, C2 => n89, 
                           A => n1333, ZN => n1332);
   U1599 : AOI22_X1 port map( A1 => n86, A2 => REGISTERS_19_23_port, B1 => n82,
                           B2 => REGISTERS_18_23_port, ZN => n1333);
   U1600 : OAI221_X1 port map( B1 => n1998, B2 => n80, C1 => n1966, C2 => n77, 
                           A => n1334, ZN => n1331);
   U1601 : AOI22_X1 port map( A1 => n74, A2 => REGISTERS_23_23_port, B1 => n70,
                           B2 => REGISTERS_22_23_port, ZN => n1334);
   U1602 : OAI221_X1 port map( B1 => n2062, B2 => n68, C1 => n2030, C2 => n65, 
                           A => n1335, ZN => n1330);
   U1603 : AOI22_X1 port map( A1 => n62, A2 => REGISTERS_27_23_port, B1 => n58,
                           B2 => REGISTERS_26_23_port, ZN => n1335);
   U1604 : OAI221_X1 port map( B1 => n2126, B2 => n56, C1 => n2094, C2 => n53, 
                           A => n1336, ZN => n1329);
   U1605 : AOI22_X1 port map( A1 => n50, A2 => REGISTERS_29_23_port, B1 => n46,
                           B2 => REGISTERS_28_23_port, ZN => n1336);
   U1606 : OAI221_X1 port map( B1 => n1806, B2 => n23, C1 => n516, C2 => n20, A
                           => n1343, ZN => n1338);
   U1607 : AOI22_X1 port map( A1 => n17, A2 => REGISTERS_11_23_port, B1 => n13,
                           B2 => REGISTERS_10_23_port, ZN => n1343);
   U1608 : OAI221_X1 port map( B1 => n2061, B2 => n69, C1 => n2029, C2 => n66, 
                           A => n1317, ZN => n1312);
   U1609 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_24_port, B1 => n58,
                           B2 => REGISTERS_26_24_port, ZN => n1317);
   U1610 : OAI221_X1 port map( B1 => n2125, B2 => n57, C1 => n2093, C2 => n54, 
                           A => n1318, ZN => n1311);
   U1611 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_24_port, B1 => n46,
                           B2 => REGISTERS_28_24_port, ZN => n1318);
   U1612 : OAI221_X1 port map( B1 => n1805, B2 => n24, C1 => n515, C2 => n21, A
                           => n1325, ZN => n1320);
   U1613 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_24_port, B1 => n13,
                           B2 => REGISTERS_10_24_port, ZN => n1325);
   U1614 : OAI221_X1 port map( B1 => n2060, B2 => n69, C1 => n2028, C2 => n66, 
                           A => n1299, ZN => n1294);
   U1615 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_25_port, B1 => n58,
                           B2 => REGISTERS_26_25_port, ZN => n1299);
   U1616 : OAI221_X1 port map( B1 => n2124, B2 => n57, C1 => n2092, C2 => n54, 
                           A => n1300, ZN => n1293);
   U1617 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_25_port, B1 => n46,
                           B2 => REGISTERS_28_25_port, ZN => n1300);
   U1618 : OAI221_X1 port map( B1 => n1804, B2 => n24, C1 => n514, C2 => n21, A
                           => n1307, ZN => n1302);
   U1619 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_25_port, B1 => n13,
                           B2 => REGISTERS_10_25_port, ZN => n1307);
   U1620 : OAI221_X1 port map( B1 => n2059, B2 => n69, C1 => n2027, C2 => n66, 
                           A => n1281, ZN => n1276);
   U1621 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_26_port, B1 => n58,
                           B2 => REGISTERS_26_26_port, ZN => n1281);
   U1622 : OAI221_X1 port map( B1 => n2123, B2 => n57, C1 => n2091, C2 => n54, 
                           A => n1282, ZN => n1275);
   U1623 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_26_port, B1 => n46,
                           B2 => REGISTERS_28_26_port, ZN => n1282);
   U1624 : OAI221_X1 port map( B1 => n1803, B2 => n24, C1 => n513, C2 => n21, A
                           => n1289, ZN => n1284);
   U1625 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_26_port, B1 => n13,
                           B2 => REGISTERS_10_26_port, ZN => n1289);
   U1626 : OAI221_X1 port map( B1 => n2058, B2 => n69, C1 => n2026, C2 => n66, 
                           A => n1263, ZN => n1258);
   U1627 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_27_port, B1 => n58,
                           B2 => REGISTERS_26_27_port, ZN => n1263);
   U1628 : OAI221_X1 port map( B1 => n2122, B2 => n57, C1 => n2090, C2 => n54, 
                           A => n1264, ZN => n1257);
   U1629 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_27_port, B1 => n46,
                           B2 => REGISTERS_28_27_port, ZN => n1264);
   U1630 : OAI221_X1 port map( B1 => n1802, B2 => n24, C1 => n512, C2 => n21, A
                           => n1271, ZN => n1266);
   U1631 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_27_port, B1 => n13,
                           B2 => REGISTERS_10_27_port, ZN => n1271);
   U1632 : OAI221_X1 port map( B1 => n2057, B2 => n69, C1 => n2025, C2 => n66, 
                           A => n1245, ZN => n1240);
   U1633 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_28_port, B1 => n58,
                           B2 => REGISTERS_26_28_port, ZN => n1245);
   U1634 : OAI221_X1 port map( B1 => n2121, B2 => n57, C1 => n2089, C2 => n54, 
                           A => n1246, ZN => n1239);
   U1635 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_28_port, B1 => n46,
                           B2 => REGISTERS_28_28_port, ZN => n1246);
   U1636 : OAI221_X1 port map( B1 => n1801, B2 => n24, C1 => n511, C2 => n21, A
                           => n1253, ZN => n1248);
   U1637 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_28_port, B1 => n13,
                           B2 => REGISTERS_10_28_port, ZN => n1253);
   U1638 : OAI221_X1 port map( B1 => n2056, B2 => n69, C1 => n2024, C2 => n66, 
                           A => n1227, ZN => n1222);
   U1639 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_29_port, B1 => n58,
                           B2 => REGISTERS_26_29_port, ZN => n1227);
   U1640 : OAI221_X1 port map( B1 => n2120, B2 => n57, C1 => n2088, C2 => n54, 
                           A => n1228, ZN => n1221);
   U1641 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_29_port, B1 => n46,
                           B2 => REGISTERS_28_29_port, ZN => n1228);
   U1642 : OAI221_X1 port map( B1 => n1800, B2 => n24, C1 => n510, C2 => n21, A
                           => n1235, ZN => n1230);
   U1643 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_29_port, B1 => n13,
                           B2 => REGISTERS_10_29_port, ZN => n1235);
   U1644 : OAI221_X1 port map( B1 => n2055, B2 => n69, C1 => n2023, C2 => n66, 
                           A => n1209, ZN => n1204);
   U1645 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_30_port, B1 => n58,
                           B2 => REGISTERS_26_30_port, ZN => n1209);
   U1646 : OAI221_X1 port map( B1 => n2119, B2 => n57, C1 => n2087, C2 => n54, 
                           A => n1210, ZN => n1203);
   U1647 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_30_port, B1 => n46,
                           B2 => REGISTERS_28_30_port, ZN => n1210);
   U1648 : OAI221_X1 port map( B1 => n1799, B2 => n24, C1 => n509, C2 => n21, A
                           => n1217, ZN => n1212);
   U1649 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_30_port, B1 => n13,
                           B2 => REGISTERS_10_30_port, ZN => n1217);
   U1650 : OAI221_X1 port map( B1 => n2054, B2 => n69, C1 => n2022, C2 => n66, 
                           A => n1169, ZN => n1154);
   U1651 : AOI22_X1 port map( A1 => n63, A2 => REGISTERS_27_31_port, B1 => n58,
                           B2 => REGISTERS_26_31_port, ZN => n1169);
   U1652 : OAI221_X1 port map( B1 => n2118, B2 => n57, C1 => n2086, C2 => n54, 
                           A => n1174, ZN => n1153);
   U1653 : AOI22_X1 port map( A1 => n51, A2 => REGISTERS_29_31_port, B1 => n46,
                           B2 => REGISTERS_28_31_port, ZN => n1174);
   U1654 : OAI221_X1 port map( B1 => n1798, B2 => n24, C1 => n508, C2 => n21, A
                           => n1193, ZN => n1178);
   U1655 : AOI22_X1 port map( A1 => n18, A2 => REGISTERS_11_31_port, B1 => n13,
                           B2 => REGISTERS_10_31_port, ZN => n1193);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n135, B1 => 
                           REGISTERS_2_24_port, B2 => n132, ZN => n699);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n135, B1 => 
                           REGISTERS_2_25_port, B2 => n132, ZN => n681);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n135, B1 => 
                           REGISTERS_2_26_port, B2 => n132, ZN => n663);
   U1659 : AOI22_X1 port map( A1 => REGISTERS_3_27_port, A2 => n135, B1 => 
                           REGISTERS_2_27_port, B2 => n132, ZN => n645);
   U1660 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n135, B1 => 
                           REGISTERS_2_28_port, B2 => n132, ZN => n627);
   U1661 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n135, B1 => 
                           REGISTERS_2_29_port, B2 => n132, ZN => n609);
   U1662 : AOI22_X1 port map( A1 => REGISTERS_3_30_port, A2 => n135, B1 => 
                           REGISTERS_2_30_port, B2 => n132, ZN => n591);
   U1663 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n135, B1 => 
                           REGISTERS_2_31_port, B2 => n132, ZN => n559);
   U1664 : AOI22_X1 port map( A1 => REGISTERS_3_0_port, A2 => n133, B1 => 
                           REGISTERS_2_0_port, B2 => n130, ZN => n1141);
   U1665 : AOI22_X1 port map( A1 => REGISTERS_3_1_port, A2 => n133, B1 => 
                           REGISTERS_2_1_port, B2 => n130, ZN => n1113);
   U1666 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n133, B1 => 
                           REGISTERS_2_2_port, B2 => n130, ZN => n1095);
   U1667 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n133, B1 => 
                           REGISTERS_2_3_port, B2 => n130, ZN => n1077);
   U1668 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n133, B1 => 
                           REGISTERS_2_4_port, B2 => n130, ZN => n1059);
   U1669 : AOI22_X1 port map( A1 => REGISTERS_3_5_port, A2 => n133, B1 => 
                           REGISTERS_2_5_port, B2 => n130, ZN => n1041);
   U1670 : AOI22_X1 port map( A1 => REGISTERS_3_6_port, A2 => n133, B1 => 
                           REGISTERS_2_6_port, B2 => n130, ZN => n1023);
   U1671 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n133, B1 => 
                           REGISTERS_2_7_port, B2 => n130, ZN => n1005);
   U1672 : AOI22_X1 port map( A1 => REGISTERS_3_8_port, A2 => n133, B1 => 
                           REGISTERS_2_8_port, B2 => n130, ZN => n987);
   U1673 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n133, B1 => 
                           REGISTERS_2_9_port, B2 => n130, ZN => n969);
   U1674 : AOI22_X1 port map( A1 => REGISTERS_3_10_port, A2 => n133, B1 => 
                           REGISTERS_2_10_port, B2 => n130, ZN => n951);
   U1675 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n133, B1 => 
                           REGISTERS_2_11_port, B2 => n130, ZN => n933);
   U1676 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n134, B1 => 
                           REGISTERS_2_12_port, B2 => n131, ZN => n915);
   U1677 : AOI22_X1 port map( A1 => REGISTERS_3_13_port, A2 => n134, B1 => 
                           REGISTERS_2_13_port, B2 => n131, ZN => n897);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n134, B1 => 
                           REGISTERS_2_14_port, B2 => n131, ZN => n879);
   U1679 : AOI22_X1 port map( A1 => REGISTERS_3_15_port, A2 => n134, B1 => 
                           REGISTERS_2_15_port, B2 => n131, ZN => n861);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n134, B1 => 
                           REGISTERS_2_16_port, B2 => n131, ZN => n843);
   U1681 : AOI22_X1 port map( A1 => REGISTERS_3_17_port, A2 => n134, B1 => 
                           REGISTERS_2_17_port, B2 => n131, ZN => n825);
   U1682 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n134, B1 => 
                           REGISTERS_2_18_port, B2 => n131, ZN => n807);
   U1683 : AOI22_X1 port map( A1 => REGISTERS_3_19_port, A2 => n134, B1 => 
                           REGISTERS_2_19_port, B2 => n131, ZN => n789);
   U1684 : AOI22_X1 port map( A1 => REGISTERS_3_20_port, A2 => n134, B1 => 
                           REGISTERS_2_20_port, B2 => n131, ZN => n771);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_3_21_port, A2 => n134, B1 => 
                           REGISTERS_2_21_port, B2 => n131, ZN => n753);
   U1686 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n134, B1 => 
                           REGISTERS_2_22_port, B2 => n131, ZN => n735);
   U1687 : AOI22_X1 port map( A1 => REGISTERS_3_23_port, A2 => n134, B1 => 
                           REGISTERS_2_23_port, B2 => n131, ZN => n717);
   U1688 : OAI21_X1 port map( B1 => n419, B2 => n45, A => n1323, ZN => n1322);
   U1689 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_24_port, B1 => n37, 
                           B2 => REGISTERS_2_24_port, ZN => n1323);
   U1690 : OAI21_X1 port map( B1 => n418, B2 => n45, A => n1305, ZN => n1304);
   U1691 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_25_port, B1 => n37, 
                           B2 => REGISTERS_2_25_port, ZN => n1305);
   U1692 : OAI21_X1 port map( B1 => n417, B2 => n45, A => n1287, ZN => n1286);
   U1693 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_26_port, B1 => n37, 
                           B2 => REGISTERS_2_26_port, ZN => n1287);
   U1694 : OAI21_X1 port map( B1 => n416, B2 => n45, A => n1269, ZN => n1268);
   U1695 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_27_port, B1 => n37, 
                           B2 => REGISTERS_2_27_port, ZN => n1269);
   U1696 : OAI21_X1 port map( B1 => n415, B2 => n45, A => n1251, ZN => n1250);
   U1697 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_28_port, B1 => n37, 
                           B2 => REGISTERS_2_28_port, ZN => n1251);
   U1698 : OAI21_X1 port map( B1 => n414, B2 => n45, A => n1233, ZN => n1232);
   U1699 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_29_port, B1 => n37, 
                           B2 => REGISTERS_2_29_port, ZN => n1233);
   U1700 : OAI21_X1 port map( B1 => n413, B2 => n45, A => n1215, ZN => n1214);
   U1701 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_30_port, B1 => n37, 
                           B2 => REGISTERS_2_30_port, ZN => n1215);
   U1702 : OAI21_X1 port map( B1 => n412, B2 => n45, A => n1183, ZN => n1180);
   U1703 : AOI22_X1 port map( A1 => n42, A2 => REGISTERS_3_31_port, B1 => n37, 
                           B2 => REGISTERS_2_31_port, ZN => n1183);
   U1704 : OAI21_X1 port map( B1 => n443, B2 => n43, A => n1765, ZN => n1764);
   U1705 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_0_port, B1 => n39, 
                           B2 => REGISTERS_2_0_port, ZN => n1765);
   U1706 : OAI21_X1 port map( B1 => n442, B2 => n43, A => n1737, ZN => n1736);
   U1707 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_1_port, B1 => n39, 
                           B2 => REGISTERS_2_1_port, ZN => n1737);
   U1708 : OAI21_X1 port map( B1 => n441, B2 => n43, A => n1719, ZN => n1718);
   U1709 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_2_port, B1 => n39, 
                           B2 => REGISTERS_2_2_port, ZN => n1719);
   U1710 : OAI21_X1 port map( B1 => n440, B2 => n43, A => n1701, ZN => n1700);
   U1711 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_3_port, B1 => n39, 
                           B2 => REGISTERS_2_3_port, ZN => n1701);
   U1712 : OAI21_X1 port map( B1 => n439, B2 => n43, A => n1683, ZN => n1682);
   U1713 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_4_port, B1 => n39, 
                           B2 => REGISTERS_2_4_port, ZN => n1683);
   U1714 : OAI21_X1 port map( B1 => n438, B2 => n43, A => n1665, ZN => n1664);
   U1715 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_5_port, B1 => n39, 
                           B2 => REGISTERS_2_5_port, ZN => n1665);
   U1716 : OAI21_X1 port map( B1 => n437, B2 => n43, A => n1647, ZN => n1646);
   U1717 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_6_port, B1 => n39, 
                           B2 => REGISTERS_2_6_port, ZN => n1647);
   U1718 : OAI21_X1 port map( B1 => n436, B2 => n43, A => n1629, ZN => n1628);
   U1719 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_7_port, B1 => n39, 
                           B2 => REGISTERS_2_7_port, ZN => n1629);
   U1720 : OAI21_X1 port map( B1 => n435, B2 => n43, A => n1611, ZN => n1610);
   U1721 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_8_port, B1 => n38, 
                           B2 => REGISTERS_2_8_port, ZN => n1611);
   U1722 : OAI21_X1 port map( B1 => n434, B2 => n43, A => n1593, ZN => n1592);
   U1723 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_9_port, B1 => n38, 
                           B2 => REGISTERS_2_9_port, ZN => n1593);
   U1724 : OAI21_X1 port map( B1 => n433, B2 => n43, A => n1575, ZN => n1574);
   U1725 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_10_port, B1 => n38, 
                           B2 => REGISTERS_2_10_port, ZN => n1575);
   U1726 : OAI21_X1 port map( B1 => n432, B2 => n43, A => n1557, ZN => n1556);
   U1727 : AOI22_X1 port map( A1 => n40, A2 => REGISTERS_3_11_port, B1 => n38, 
                           B2 => REGISTERS_2_11_port, ZN => n1557);
   U1728 : OAI21_X1 port map( B1 => n431, B2 => n44, A => n1539, ZN => n1538);
   U1729 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_12_port, B1 => n38, 
                           B2 => REGISTERS_2_12_port, ZN => n1539);
   U1730 : OAI21_X1 port map( B1 => n430, B2 => n44, A => n1521, ZN => n1520);
   U1731 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_13_port, B1 => n38, 
                           B2 => REGISTERS_2_13_port, ZN => n1521);
   U1732 : OAI21_X1 port map( B1 => n429, B2 => n44, A => n1503, ZN => n1502);
   U1733 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_14_port, B1 => n38, 
                           B2 => REGISTERS_2_14_port, ZN => n1503);
   U1734 : OAI21_X1 port map( B1 => n428, B2 => n44, A => n1485, ZN => n1484);
   U1735 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_15_port, B1 => n38, 
                           B2 => REGISTERS_2_15_port, ZN => n1485);
   U1736 : OAI21_X1 port map( B1 => n427, B2 => n44, A => n1467, ZN => n1466);
   U1737 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_16_port, B1 => n38, 
                           B2 => REGISTERS_2_16_port, ZN => n1467);
   U1738 : OAI21_X1 port map( B1 => n426, B2 => n44, A => n1449, ZN => n1448);
   U1739 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_17_port, B1 => n38, 
                           B2 => REGISTERS_2_17_port, ZN => n1449);
   U1740 : OAI21_X1 port map( B1 => n425, B2 => n44, A => n1431, ZN => n1430);
   U1741 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_18_port, B1 => n38, 
                           B2 => REGISTERS_2_18_port, ZN => n1431);
   U1742 : OAI21_X1 port map( B1 => n424, B2 => n44, A => n1413, ZN => n1412);
   U1743 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_19_port, B1 => n38, 
                           B2 => REGISTERS_2_19_port, ZN => n1413);
   U1744 : OAI21_X1 port map( B1 => n423, B2 => n44, A => n1395, ZN => n1394);
   U1745 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_20_port, B1 => n37, 
                           B2 => REGISTERS_2_20_port, ZN => n1395);
   U1746 : OAI21_X1 port map( B1 => n422, B2 => n44, A => n1377, ZN => n1376);
   U1747 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_21_port, B1 => n37, 
                           B2 => REGISTERS_2_21_port, ZN => n1377);
   U1748 : OAI21_X1 port map( B1 => n421, B2 => n44, A => n1359, ZN => n1358);
   U1749 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_22_port, B1 => n37, 
                           B2 => REGISTERS_2_22_port, ZN => n1359);
   U1750 : OAI21_X1 port map( B1 => n420, B2 => n44, A => n1341, ZN => n1340);
   U1751 : AOI22_X1 port map( A1 => n41, A2 => REGISTERS_3_23_port, B1 => n37, 
                           B2 => REGISTERS_2_23_port, ZN => n1341);
   U1752 : INV_X1 port map( A => ADD_WR(2), ZN => n409);
   U1753 : INV_X1 port map( A => ADD_WR(0), ZN => n411);
   U1754 : INV_X1 port map( A => ADD_WR(1), ZN => n410);
   U1755 : INV_X1 port map( A => ADD_WR(3), ZN => n408);
   U1756 : INV_X1 port map( A => ADD_WR(4), ZN => n407);
   U1757 : OR2_X1 port map( A1 => RE, A2 => n391, ZN => N307);
   U1758 : INV_X1 port map( A => REGISTERS_17_0_port, ZN => n1957);
   U1759 : INV_X1 port map( A => REGISTERS_21_0_port, ZN => n2021);
   U1760 : INV_X1 port map( A => REGISTERS_25_0_port, ZN => n2085);
   U1761 : INV_X1 port map( A => REGISTERS_31_0_port, ZN => n2149);
   U1762 : INV_X1 port map( A => REGISTERS_5_0_port, ZN => n507);
   U1763 : INV_X1 port map( A => REGISTERS_9_0_port, ZN => n1829);
   U1764 : INV_X1 port map( A => REGISTERS_13_0_port, ZN => n1893);
   U1765 : INV_X1 port map( A => REGISTERS_17_1_port, ZN => n1956);
   U1766 : INV_X1 port map( A => REGISTERS_21_1_port, ZN => n2020);
   U1767 : INV_X1 port map( A => REGISTERS_25_1_port, ZN => n2084);
   U1768 : INV_X1 port map( A => REGISTERS_31_1_port, ZN => n2148);
   U1769 : INV_X1 port map( A => REGISTERS_5_1_port, ZN => n506);
   U1770 : INV_X1 port map( A => REGISTERS_9_1_port, ZN => n1828);
   U1771 : INV_X1 port map( A => REGISTERS_13_1_port, ZN => n1892);
   U1772 : INV_X1 port map( A => REGISTERS_17_2_port, ZN => n1955);
   U1773 : INV_X1 port map( A => REGISTERS_21_2_port, ZN => n2019);
   U1774 : INV_X1 port map( A => REGISTERS_25_2_port, ZN => n2083);
   U1775 : INV_X1 port map( A => REGISTERS_31_2_port, ZN => n2147);
   U1776 : INV_X1 port map( A => REGISTERS_5_2_port, ZN => n505);
   U1777 : INV_X1 port map( A => REGISTERS_9_2_port, ZN => n1827);
   U1778 : INV_X1 port map( A => REGISTERS_13_2_port, ZN => n1891);
   U1779 : INV_X1 port map( A => REGISTERS_17_3_port, ZN => n1954);
   U1780 : INV_X1 port map( A => REGISTERS_21_3_port, ZN => n2018);
   U1781 : INV_X1 port map( A => REGISTERS_25_3_port, ZN => n2082);
   U1782 : INV_X1 port map( A => REGISTERS_31_3_port, ZN => n2146);
   U1783 : INV_X1 port map( A => REGISTERS_5_3_port, ZN => n504);
   U1784 : INV_X1 port map( A => REGISTERS_9_3_port, ZN => n1826);
   U1785 : INV_X1 port map( A => REGISTERS_13_3_port, ZN => n1890);
   U1786 : INV_X1 port map( A => REGISTERS_17_4_port, ZN => n1953);
   U1787 : INV_X1 port map( A => REGISTERS_21_4_port, ZN => n2017);
   U1788 : INV_X1 port map( A => REGISTERS_25_4_port, ZN => n2081);
   U1789 : INV_X1 port map( A => REGISTERS_31_4_port, ZN => n2145);
   U1790 : INV_X1 port map( A => REGISTERS_5_4_port, ZN => n503);
   U1791 : INV_X1 port map( A => REGISTERS_9_4_port, ZN => n1825);
   U1792 : INV_X1 port map( A => REGISTERS_13_4_port, ZN => n1889);
   U1793 : INV_X1 port map( A => REGISTERS_17_5_port, ZN => n1952);
   U1794 : INV_X1 port map( A => REGISTERS_21_5_port, ZN => n2016);
   U1795 : INV_X1 port map( A => REGISTERS_25_5_port, ZN => n2080);
   U1796 : INV_X1 port map( A => REGISTERS_31_5_port, ZN => n2144);
   U1797 : INV_X1 port map( A => REGISTERS_5_5_port, ZN => n502);
   U1798 : INV_X1 port map( A => REGISTERS_9_5_port, ZN => n1824);
   U1799 : INV_X1 port map( A => REGISTERS_13_5_port, ZN => n1888);
   U1800 : INV_X1 port map( A => REGISTERS_17_6_port, ZN => n1951);
   U1801 : INV_X1 port map( A => REGISTERS_21_6_port, ZN => n2015);
   U1802 : INV_X1 port map( A => REGISTERS_25_6_port, ZN => n2079);
   U1803 : INV_X1 port map( A => REGISTERS_31_6_port, ZN => n2143);
   U1804 : INV_X1 port map( A => REGISTERS_5_6_port, ZN => n501);
   U1805 : INV_X1 port map( A => REGISTERS_9_6_port, ZN => n1823);
   U1806 : INV_X1 port map( A => REGISTERS_13_6_port, ZN => n1887);
   U1807 : INV_X1 port map( A => REGISTERS_17_7_port, ZN => n1950);
   U1808 : INV_X1 port map( A => REGISTERS_21_7_port, ZN => n2014);
   U1809 : INV_X1 port map( A => REGISTERS_25_7_port, ZN => n2078);
   U1810 : INV_X1 port map( A => REGISTERS_31_7_port, ZN => n2142);
   U1811 : INV_X1 port map( A => REGISTERS_5_7_port, ZN => n500);
   U1812 : INV_X1 port map( A => REGISTERS_9_7_port, ZN => n1822);
   U1813 : INV_X1 port map( A => REGISTERS_13_7_port, ZN => n1886);
   U1814 : INV_X1 port map( A => REGISTERS_17_8_port, ZN => n1949);
   U1815 : INV_X1 port map( A => REGISTERS_21_8_port, ZN => n2013);
   U1816 : INV_X1 port map( A => REGISTERS_25_8_port, ZN => n2077);
   U1817 : INV_X1 port map( A => REGISTERS_31_8_port, ZN => n2141);
   U1818 : INV_X1 port map( A => REGISTERS_5_8_port, ZN => n499);
   U1819 : INV_X1 port map( A => REGISTERS_9_8_port, ZN => n1821);
   U1820 : INV_X1 port map( A => REGISTERS_13_8_port, ZN => n1885);
   U1821 : INV_X1 port map( A => REGISTERS_17_9_port, ZN => n1948);
   U1822 : INV_X1 port map( A => REGISTERS_21_9_port, ZN => n2012);
   U1823 : INV_X1 port map( A => REGISTERS_25_9_port, ZN => n2076);
   U1824 : INV_X1 port map( A => REGISTERS_31_9_port, ZN => n2140);
   U1825 : INV_X1 port map( A => REGISTERS_5_9_port, ZN => n498);
   U1826 : INV_X1 port map( A => REGISTERS_9_9_port, ZN => n1820);
   U1827 : INV_X1 port map( A => REGISTERS_13_9_port, ZN => n1884);
   U1828 : INV_X1 port map( A => REGISTERS_17_10_port, ZN => n1947);
   U1829 : INV_X1 port map( A => REGISTERS_21_10_port, ZN => n2011);
   U1830 : INV_X1 port map( A => REGISTERS_25_10_port, ZN => n2075);
   U1831 : INV_X1 port map( A => REGISTERS_31_10_port, ZN => n2139);
   U1832 : INV_X1 port map( A => REGISTERS_5_10_port, ZN => n497);
   U1833 : INV_X1 port map( A => REGISTERS_9_10_port, ZN => n1819);
   U1834 : INV_X1 port map( A => REGISTERS_13_10_port, ZN => n1883);
   U1835 : INV_X1 port map( A => REGISTERS_17_11_port, ZN => n1946);
   U1836 : INV_X1 port map( A => REGISTERS_21_11_port, ZN => n2010);
   U1837 : INV_X1 port map( A => REGISTERS_25_11_port, ZN => n2074);
   U1838 : INV_X1 port map( A => REGISTERS_31_11_port, ZN => n2138);
   U1839 : INV_X1 port map( A => REGISTERS_5_11_port, ZN => n496);
   U1840 : INV_X1 port map( A => REGISTERS_9_11_port, ZN => n1818);
   U1841 : INV_X1 port map( A => REGISTERS_13_11_port, ZN => n1882);
   U1842 : INV_X1 port map( A => REGISTERS_17_12_port, ZN => n1945);
   U1843 : INV_X1 port map( A => REGISTERS_21_12_port, ZN => n2009);
   U1844 : INV_X1 port map( A => REGISTERS_25_12_port, ZN => n2073);
   U1845 : INV_X1 port map( A => REGISTERS_31_12_port, ZN => n2137);
   U1846 : INV_X1 port map( A => REGISTERS_5_12_port, ZN => n495);
   U1847 : INV_X1 port map( A => REGISTERS_9_12_port, ZN => n1817);
   U1848 : INV_X1 port map( A => REGISTERS_13_12_port, ZN => n1881);
   U1849 : INV_X1 port map( A => REGISTERS_17_13_port, ZN => n1944);
   U1850 : INV_X1 port map( A => REGISTERS_21_13_port, ZN => n2008);
   U1851 : INV_X1 port map( A => REGISTERS_25_13_port, ZN => n2072);
   U1852 : INV_X1 port map( A => REGISTERS_31_13_port, ZN => n2136);
   U1853 : INV_X1 port map( A => REGISTERS_5_13_port, ZN => n494);
   U1854 : INV_X1 port map( A => REGISTERS_9_13_port, ZN => n1816);
   U1855 : INV_X1 port map( A => REGISTERS_13_13_port, ZN => n1880);
   U1856 : INV_X1 port map( A => REGISTERS_17_14_port, ZN => n1943);
   U1857 : INV_X1 port map( A => REGISTERS_21_14_port, ZN => n2007);
   U1858 : INV_X1 port map( A => REGISTERS_25_14_port, ZN => n2071);
   U1859 : INV_X1 port map( A => REGISTERS_31_14_port, ZN => n2135);
   U1860 : INV_X1 port map( A => REGISTERS_5_14_port, ZN => n493);
   U1861 : INV_X1 port map( A => REGISTERS_9_14_port, ZN => n1815);
   U1862 : INV_X1 port map( A => REGISTERS_13_14_port, ZN => n1879);
   U1863 : INV_X1 port map( A => REGISTERS_17_15_port, ZN => n1942);
   U1864 : INV_X1 port map( A => REGISTERS_21_15_port, ZN => n2006);
   U1865 : INV_X1 port map( A => REGISTERS_25_15_port, ZN => n2070);
   U1866 : INV_X1 port map( A => REGISTERS_31_15_port, ZN => n2134);
   U1867 : INV_X1 port map( A => REGISTERS_5_15_port, ZN => n492);
   U1868 : INV_X1 port map( A => REGISTERS_9_15_port, ZN => n1814);
   U1869 : INV_X1 port map( A => REGISTERS_13_15_port, ZN => n1878);
   U1870 : INV_X1 port map( A => REGISTERS_17_16_port, ZN => n1941);
   U1871 : INV_X1 port map( A => REGISTERS_21_16_port, ZN => n2005);
   U1872 : INV_X1 port map( A => REGISTERS_25_16_port, ZN => n2069);
   U1873 : INV_X1 port map( A => REGISTERS_31_16_port, ZN => n2133);
   U1874 : INV_X1 port map( A => REGISTERS_5_16_port, ZN => n491);
   U1875 : INV_X1 port map( A => REGISTERS_9_16_port, ZN => n1813);
   U1876 : INV_X1 port map( A => REGISTERS_13_16_port, ZN => n1877);
   U1877 : INV_X1 port map( A => REGISTERS_17_17_port, ZN => n1940);
   U1878 : INV_X1 port map( A => REGISTERS_21_17_port, ZN => n2004);
   U1879 : INV_X1 port map( A => REGISTERS_25_17_port, ZN => n2068);
   U1880 : INV_X1 port map( A => REGISTERS_31_17_port, ZN => n2132);
   U1881 : INV_X1 port map( A => REGISTERS_5_17_port, ZN => n490);
   U1882 : INV_X1 port map( A => REGISTERS_9_17_port, ZN => n1812);
   U1883 : INV_X1 port map( A => REGISTERS_13_17_port, ZN => n1876);
   U1884 : INV_X1 port map( A => REGISTERS_17_18_port, ZN => n1939);
   U1885 : INV_X1 port map( A => REGISTERS_21_18_port, ZN => n2003);
   U1886 : INV_X1 port map( A => REGISTERS_25_18_port, ZN => n2067);
   U1887 : INV_X1 port map( A => REGISTERS_31_18_port, ZN => n2131);
   U1888 : INV_X1 port map( A => REGISTERS_5_18_port, ZN => n489);
   U1889 : INV_X1 port map( A => REGISTERS_9_18_port, ZN => n1811);
   U1890 : INV_X1 port map( A => REGISTERS_13_18_port, ZN => n1875);
   U1891 : INV_X1 port map( A => REGISTERS_17_19_port, ZN => n1938);
   U1892 : INV_X1 port map( A => REGISTERS_21_19_port, ZN => n2002);
   U1893 : INV_X1 port map( A => REGISTERS_25_19_port, ZN => n2066);
   U1894 : INV_X1 port map( A => REGISTERS_31_19_port, ZN => n2130);
   U1895 : INV_X1 port map( A => REGISTERS_5_19_port, ZN => n488);
   U1896 : INV_X1 port map( A => REGISTERS_9_19_port, ZN => n1810);
   U1897 : INV_X1 port map( A => REGISTERS_13_19_port, ZN => n1874);
   U1898 : INV_X1 port map( A => REGISTERS_17_20_port, ZN => n1937);
   U1899 : INV_X1 port map( A => REGISTERS_21_20_port, ZN => n2001);
   U1900 : INV_X1 port map( A => REGISTERS_25_20_port, ZN => n2065);
   U1901 : INV_X1 port map( A => REGISTERS_31_20_port, ZN => n2129);
   U1902 : INV_X1 port map( A => REGISTERS_5_20_port, ZN => n487);
   U1903 : INV_X1 port map( A => REGISTERS_9_20_port, ZN => n1809);
   U1904 : INV_X1 port map( A => REGISTERS_13_20_port, ZN => n1873);
   U1917 : INV_X1 port map( A => REGISTERS_17_21_port, ZN => n1936);
   U1918 : INV_X1 port map( A => REGISTERS_21_21_port, ZN => n2000);
   U1919 : INV_X1 port map( A => REGISTERS_25_21_port, ZN => n2064);
   U1920 : INV_X1 port map( A => REGISTERS_31_21_port, ZN => n2128);
   U1921 : INV_X1 port map( A => REGISTERS_5_21_port, ZN => n486);
   U1922 : INV_X1 port map( A => REGISTERS_9_21_port, ZN => n1808);
   U1923 : INV_X1 port map( A => REGISTERS_13_21_port, ZN => n1872);
   U1924 : INV_X1 port map( A => REGISTERS_17_22_port, ZN => n1935);
   U1925 : INV_X1 port map( A => REGISTERS_21_22_port, ZN => n1999);
   U1926 : INV_X1 port map( A => REGISTERS_25_22_port, ZN => n2063);
   U1927 : INV_X1 port map( A => REGISTERS_31_22_port, ZN => n2127);
   U1928 : INV_X1 port map( A => REGISTERS_5_22_port, ZN => n485);
   U1929 : INV_X1 port map( A => REGISTERS_9_22_port, ZN => n1807);
   U1930 : INV_X1 port map( A => REGISTERS_13_22_port, ZN => n1871);
   U1931 : INV_X1 port map( A => REGISTERS_17_23_port, ZN => n1934);
   U1932 : INV_X1 port map( A => REGISTERS_21_23_port, ZN => n1998);
   U1933 : INV_X1 port map( A => REGISTERS_25_23_port, ZN => n2062);
   U1934 : INV_X1 port map( A => REGISTERS_31_23_port, ZN => n2126);
   U1935 : INV_X1 port map( A => REGISTERS_5_23_port, ZN => n484);
   U1936 : INV_X1 port map( A => REGISTERS_9_23_port, ZN => n1806);
   U1937 : INV_X1 port map( A => REGISTERS_13_23_port, ZN => n1870);
   U1938 : INV_X1 port map( A => REGISTERS_17_24_port, ZN => n1933);
   U1939 : INV_X1 port map( A => REGISTERS_21_24_port, ZN => n1997);
   U1940 : INV_X1 port map( A => REGISTERS_25_24_port, ZN => n2061);
   U1941 : INV_X1 port map( A => REGISTERS_31_24_port, ZN => n2125);
   U1942 : INV_X1 port map( A => REGISTERS_5_24_port, ZN => n483);
   U1943 : INV_X1 port map( A => REGISTERS_9_24_port, ZN => n1805);
   U1944 : INV_X1 port map( A => REGISTERS_13_24_port, ZN => n1869);
   U1945 : INV_X1 port map( A => REGISTERS_17_25_port, ZN => n1932);
   U1946 : INV_X1 port map( A => REGISTERS_21_25_port, ZN => n1996);
   U1947 : INV_X1 port map( A => REGISTERS_25_25_port, ZN => n2060);
   U1948 : INV_X1 port map( A => REGISTERS_31_25_port, ZN => n2124);
   U1949 : INV_X1 port map( A => REGISTERS_5_25_port, ZN => n482);
   U1950 : INV_X1 port map( A => REGISTERS_9_25_port, ZN => n1804);
   U1951 : INV_X1 port map( A => REGISTERS_13_25_port, ZN => n1868);
   U1952 : INV_X1 port map( A => REGISTERS_17_26_port, ZN => n1931);
   U1953 : INV_X1 port map( A => REGISTERS_21_26_port, ZN => n1995);
   U1954 : INV_X1 port map( A => REGISTERS_25_26_port, ZN => n2059);
   U1955 : INV_X1 port map( A => REGISTERS_31_26_port, ZN => n2123);
   U1956 : INV_X1 port map( A => REGISTERS_5_26_port, ZN => n481);
   U1957 : INV_X1 port map( A => REGISTERS_9_26_port, ZN => n1803);
   U1958 : INV_X1 port map( A => REGISTERS_13_26_port, ZN => n1867);
   U1959 : INV_X1 port map( A => REGISTERS_17_27_port, ZN => n1930);
   U1960 : INV_X1 port map( A => REGISTERS_21_27_port, ZN => n1994);
   U1961 : INV_X1 port map( A => REGISTERS_25_27_port, ZN => n2058);
   U1962 : INV_X1 port map( A => REGISTERS_31_27_port, ZN => n2122);
   U1963 : INV_X1 port map( A => REGISTERS_5_27_port, ZN => n480);
   U1964 : INV_X1 port map( A => REGISTERS_9_27_port, ZN => n1802);
   U1965 : INV_X1 port map( A => REGISTERS_13_27_port, ZN => n1866);
   U1966 : INV_X1 port map( A => REGISTERS_17_28_port, ZN => n1929);
   U1967 : INV_X1 port map( A => REGISTERS_21_28_port, ZN => n1993);
   U1968 : INV_X1 port map( A => REGISTERS_25_28_port, ZN => n2057);
   U1969 : INV_X1 port map( A => REGISTERS_31_28_port, ZN => n2121);
   U1970 : INV_X1 port map( A => REGISTERS_5_28_port, ZN => n479);
   U1971 : INV_X1 port map( A => REGISTERS_9_28_port, ZN => n1801);
   U1972 : INV_X1 port map( A => REGISTERS_13_28_port, ZN => n1865);
   U1973 : INV_X1 port map( A => REGISTERS_17_29_port, ZN => n1928);
   U1974 : INV_X1 port map( A => REGISTERS_21_29_port, ZN => n1992);
   U1975 : INV_X1 port map( A => REGISTERS_25_29_port, ZN => n2056);
   U1976 : INV_X1 port map( A => REGISTERS_31_29_port, ZN => n2120);
   U1977 : INV_X1 port map( A => REGISTERS_5_29_port, ZN => n478);
   U1978 : INV_X1 port map( A => REGISTERS_9_29_port, ZN => n1800);
   U1979 : INV_X1 port map( A => REGISTERS_13_29_port, ZN => n1864);
   U1980 : INV_X1 port map( A => REGISTERS_17_30_port, ZN => n1927);
   U1981 : INV_X1 port map( A => REGISTERS_21_30_port, ZN => n1991);
   U1982 : INV_X1 port map( A => REGISTERS_25_30_port, ZN => n2055);
   U1983 : INV_X1 port map( A => REGISTERS_31_30_port, ZN => n2119);
   U1984 : INV_X1 port map( A => REGISTERS_5_30_port, ZN => n477);
   U1985 : INV_X1 port map( A => REGISTERS_9_30_port, ZN => n1799);
   U1986 : INV_X1 port map( A => REGISTERS_13_30_port, ZN => n1863);
   U1987 : INV_X1 port map( A => REGISTERS_17_31_port, ZN => n1926);
   U1988 : INV_X1 port map( A => REGISTERS_21_31_port, ZN => n1990);
   U1989 : INV_X1 port map( A => REGISTERS_25_31_port, ZN => n2054);
   U1990 : INV_X1 port map( A => REGISTERS_31_31_port, ZN => n2118);
   U1991 : INV_X1 port map( A => REGISTERS_5_31_port, ZN => n476);
   U1992 : INV_X1 port map( A => REGISTERS_9_31_port, ZN => n1798);
   U1993 : INV_X1 port map( A => REGISTERS_13_31_port, ZN => n1862);
   U1994 : INV_X1 port map( A => REGISTERS_1_0_port, ZN => n443);
   U1995 : INV_X1 port map( A => REGISTERS_1_1_port, ZN => n442);
   U1996 : INV_X1 port map( A => REGISTERS_1_2_port, ZN => n441);
   U1997 : INV_X1 port map( A => REGISTERS_1_3_port, ZN => n440);
   U1998 : INV_X1 port map( A => REGISTERS_1_4_port, ZN => n439);
   U1999 : INV_X1 port map( A => REGISTERS_1_5_port, ZN => n438);
   U2000 : INV_X1 port map( A => REGISTERS_1_6_port, ZN => n437);
   U2001 : INV_X1 port map( A => REGISTERS_1_7_port, ZN => n436);
   U2002 : INV_X1 port map( A => REGISTERS_1_8_port, ZN => n435);
   U2003 : INV_X1 port map( A => REGISTERS_1_9_port, ZN => n434);
   U2004 : INV_X1 port map( A => REGISTERS_1_10_port, ZN => n433);
   U2005 : INV_X1 port map( A => REGISTERS_1_11_port, ZN => n432);
   U2006 : INV_X1 port map( A => REGISTERS_1_12_port, ZN => n431);
   U2007 : INV_X1 port map( A => REGISTERS_1_13_port, ZN => n430);
   U2008 : INV_X1 port map( A => REGISTERS_1_14_port, ZN => n429);
   U2009 : INV_X1 port map( A => REGISTERS_1_15_port, ZN => n428);
   U2010 : INV_X1 port map( A => REGISTERS_1_16_port, ZN => n427);
   U2011 : INV_X1 port map( A => REGISTERS_1_17_port, ZN => n426);
   U2012 : INV_X1 port map( A => REGISTERS_1_18_port, ZN => n425);
   U2013 : INV_X1 port map( A => REGISTERS_1_19_port, ZN => n424);
   U2014 : INV_X1 port map( A => REGISTERS_1_20_port, ZN => n423);
   U2015 : INV_X1 port map( A => REGISTERS_1_21_port, ZN => n422);
   U2016 : INV_X1 port map( A => REGISTERS_1_22_port, ZN => n421);
   U2017 : INV_X1 port map( A => REGISTERS_1_23_port, ZN => n420);
   U2018 : INV_X1 port map( A => REGISTERS_1_24_port, ZN => n419);
   U2019 : INV_X1 port map( A => REGISTERS_1_25_port, ZN => n418);
   U2020 : INV_X1 port map( A => REGISTERS_1_26_port, ZN => n417);
   U2021 : INV_X1 port map( A => REGISTERS_1_27_port, ZN => n416);
   U2022 : INV_X1 port map( A => REGISTERS_1_28_port, ZN => n415);
   U2023 : INV_X1 port map( A => REGISTERS_1_29_port, ZN => n414);
   U2024 : INV_X1 port map( A => REGISTERS_1_30_port, ZN => n413);
   U2025 : INV_X1 port map( A => REGISTERS_1_31_port, ZN => n412);
   U2026 : INV_X1 port map( A => REGISTERS_16_0_port, ZN => n1925);
   U2027 : INV_X1 port map( A => REGISTERS_20_0_port, ZN => n1989);
   U2028 : INV_X1 port map( A => REGISTERS_24_0_port, ZN => n2053);
   U2029 : INV_X1 port map( A => REGISTERS_30_0_port, ZN => n2117);
   U2030 : INV_X1 port map( A => REGISTERS_4_0_port, ZN => n475);
   U2031 : INV_X1 port map( A => REGISTERS_8_0_port, ZN => n1797);
   U2032 : INV_X1 port map( A => REGISTERS_12_0_port, ZN => n1861);
   U2033 : INV_X1 port map( A => REGISTERS_16_1_port, ZN => n1924);
   U2034 : INV_X1 port map( A => REGISTERS_20_1_port, ZN => n1988);
   U2035 : INV_X1 port map( A => REGISTERS_24_1_port, ZN => n2052);
   U2036 : INV_X1 port map( A => REGISTERS_30_1_port, ZN => n2116);
   U2037 : INV_X1 port map( A => REGISTERS_4_1_port, ZN => n474);
   U2038 : INV_X1 port map( A => REGISTERS_8_1_port, ZN => n1796);
   U2039 : INV_X1 port map( A => REGISTERS_12_1_port, ZN => n1860);
   U2040 : INV_X1 port map( A => REGISTERS_16_2_port, ZN => n1923);
   U2041 : INV_X1 port map( A => REGISTERS_20_2_port, ZN => n1987);
   U2042 : INV_X1 port map( A => REGISTERS_24_2_port, ZN => n2051);
   U2043 : INV_X1 port map( A => REGISTERS_30_2_port, ZN => n2115);
   U2044 : INV_X1 port map( A => REGISTERS_4_2_port, ZN => n473);
   U2045 : INV_X1 port map( A => REGISTERS_8_2_port, ZN => n1795);
   U2046 : INV_X1 port map( A => REGISTERS_12_2_port, ZN => n1859);
   U2047 : INV_X1 port map( A => REGISTERS_16_3_port, ZN => n1922);
   U2048 : INV_X1 port map( A => REGISTERS_20_3_port, ZN => n1986);
   U2049 : INV_X1 port map( A => REGISTERS_24_3_port, ZN => n2050);
   U2050 : INV_X1 port map( A => REGISTERS_30_3_port, ZN => n2114);
   U2051 : INV_X1 port map( A => REGISTERS_4_3_port, ZN => n472);
   U2052 : INV_X1 port map( A => REGISTERS_8_3_port, ZN => n1794);
   U2053 : INV_X1 port map( A => REGISTERS_12_3_port, ZN => n1858);
   U2054 : INV_X1 port map( A => REGISTERS_16_4_port, ZN => n1921);
   U2055 : INV_X1 port map( A => REGISTERS_20_4_port, ZN => n1985);
   U2056 : INV_X1 port map( A => REGISTERS_24_4_port, ZN => n2049);
   U2057 : INV_X1 port map( A => REGISTERS_30_4_port, ZN => n2113);
   U2058 : INV_X1 port map( A => REGISTERS_4_4_port, ZN => n471);
   U2059 : INV_X1 port map( A => REGISTERS_8_4_port, ZN => n1793);
   U2060 : INV_X1 port map( A => REGISTERS_12_4_port, ZN => n1857);
   U2061 : INV_X1 port map( A => REGISTERS_16_5_port, ZN => n1920);
   U2062 : INV_X1 port map( A => REGISTERS_20_5_port, ZN => n1984);
   U2063 : INV_X1 port map( A => REGISTERS_24_5_port, ZN => n2048);
   U2064 : INV_X1 port map( A => REGISTERS_30_5_port, ZN => n2112);
   U2065 : INV_X1 port map( A => REGISTERS_4_5_port, ZN => n470);
   U2066 : INV_X1 port map( A => REGISTERS_8_5_port, ZN => n1792);
   U2067 : INV_X1 port map( A => REGISTERS_12_5_port, ZN => n1856);
   U2068 : INV_X1 port map( A => REGISTERS_16_6_port, ZN => n1919);
   U2069 : INV_X1 port map( A => REGISTERS_20_6_port, ZN => n1983);
   U2070 : INV_X1 port map( A => REGISTERS_24_6_port, ZN => n2047);
   U2071 : INV_X1 port map( A => REGISTERS_30_6_port, ZN => n2111);
   U2072 : INV_X1 port map( A => REGISTERS_4_6_port, ZN => n469);
   U2073 : INV_X1 port map( A => REGISTERS_8_6_port, ZN => n1791);
   U2074 : INV_X1 port map( A => REGISTERS_12_6_port, ZN => n1855);
   U2075 : INV_X1 port map( A => REGISTERS_16_7_port, ZN => n1918);
   U2076 : INV_X1 port map( A => REGISTERS_20_7_port, ZN => n1982);
   U2077 : INV_X1 port map( A => REGISTERS_24_7_port, ZN => n2046);
   U2078 : INV_X1 port map( A => REGISTERS_30_7_port, ZN => n2110);
   U2079 : INV_X1 port map( A => REGISTERS_4_7_port, ZN => n468);
   U2080 : INV_X1 port map( A => REGISTERS_8_7_port, ZN => n1790);
   U2081 : INV_X1 port map( A => REGISTERS_12_7_port, ZN => n1854);
   U2082 : INV_X1 port map( A => REGISTERS_16_8_port, ZN => n1917);
   U2083 : INV_X1 port map( A => REGISTERS_20_8_port, ZN => n1981);
   U2084 : INV_X1 port map( A => REGISTERS_24_8_port, ZN => n2045);
   U2085 : INV_X1 port map( A => REGISTERS_30_8_port, ZN => n2109);
   U2086 : INV_X1 port map( A => REGISTERS_4_8_port, ZN => n467);
   U2087 : INV_X1 port map( A => REGISTERS_8_8_port, ZN => n1789);
   U2088 : INV_X1 port map( A => REGISTERS_12_8_port, ZN => n1853);
   U2089 : INV_X1 port map( A => REGISTERS_16_9_port, ZN => n1916);
   U2090 : INV_X1 port map( A => REGISTERS_20_9_port, ZN => n1980);
   U2091 : INV_X1 port map( A => REGISTERS_24_9_port, ZN => n2044);
   U2092 : INV_X1 port map( A => REGISTERS_30_9_port, ZN => n2108);
   U2093 : INV_X1 port map( A => REGISTERS_4_9_port, ZN => n466);
   U2094 : INV_X1 port map( A => REGISTERS_8_9_port, ZN => n1788);
   U2095 : INV_X1 port map( A => REGISTERS_12_9_port, ZN => n1852);
   U2096 : INV_X1 port map( A => REGISTERS_16_10_port, ZN => n1915);
   U2097 : INV_X1 port map( A => REGISTERS_20_10_port, ZN => n1979);
   U2098 : INV_X1 port map( A => REGISTERS_24_10_port, ZN => n2043);
   U2099 : INV_X1 port map( A => REGISTERS_30_10_port, ZN => n2107);
   U2100 : INV_X1 port map( A => REGISTERS_4_10_port, ZN => n465);
   U2101 : INV_X1 port map( A => REGISTERS_8_10_port, ZN => n1787);
   U2102 : INV_X1 port map( A => REGISTERS_12_10_port, ZN => n1851);
   U2103 : INV_X1 port map( A => REGISTERS_16_11_port, ZN => n1914);
   U2104 : INV_X1 port map( A => REGISTERS_20_11_port, ZN => n1978);
   U2105 : INV_X1 port map( A => REGISTERS_24_11_port, ZN => n2042);
   U2106 : INV_X1 port map( A => REGISTERS_30_11_port, ZN => n2106);
   U2107 : INV_X1 port map( A => REGISTERS_4_11_port, ZN => n464);
   U2108 : INV_X1 port map( A => REGISTERS_8_11_port, ZN => n1182);
   U2109 : INV_X1 port map( A => REGISTERS_12_11_port, ZN => n1850);
   U2110 : INV_X1 port map( A => REGISTERS_16_12_port, ZN => n1913);
   U2111 : INV_X1 port map( A => REGISTERS_20_12_port, ZN => n1977);
   U2112 : INV_X1 port map( A => REGISTERS_24_12_port, ZN => n2041);
   U2113 : INV_X1 port map( A => REGISTERS_30_12_port, ZN => n2105);
   U2114 : INV_X1 port map( A => REGISTERS_4_12_port, ZN => n463);
   U2115 : INV_X1 port map( A => REGISTERS_8_12_port, ZN => n558);
   U2116 : INV_X1 port map( A => REGISTERS_12_12_port, ZN => n1849);
   U2117 : INV_X1 port map( A => REGISTERS_16_13_port, ZN => n1912);
   U2118 : INV_X1 port map( A => REGISTERS_20_13_port, ZN => n1976);
   U2119 : INV_X1 port map( A => REGISTERS_24_13_port, ZN => n2040);
   U2120 : INV_X1 port map( A => REGISTERS_30_13_port, ZN => n2104);
   U2121 : INV_X1 port map( A => REGISTERS_4_13_port, ZN => n462);
   U2122 : INV_X1 port map( A => REGISTERS_8_13_port, ZN => n526);
   U2123 : INV_X1 port map( A => REGISTERS_12_13_port, ZN => n1848);
   U2124 : INV_X1 port map( A => REGISTERS_16_14_port, ZN => n1911);
   U2125 : INV_X1 port map( A => REGISTERS_20_14_port, ZN => n1975);
   U2126 : INV_X1 port map( A => REGISTERS_24_14_port, ZN => n2039);
   U2127 : INV_X1 port map( A => REGISTERS_30_14_port, ZN => n2103);
   U2128 : INV_X1 port map( A => REGISTERS_4_14_port, ZN => n461);
   U2129 : INV_X1 port map( A => REGISTERS_8_14_port, ZN => n525);
   U2130 : INV_X1 port map( A => REGISTERS_12_14_port, ZN => n1847);
   U2131 : INV_X1 port map( A => REGISTERS_16_15_port, ZN => n1910);
   U2132 : INV_X1 port map( A => REGISTERS_20_15_port, ZN => n1974);
   U2133 : INV_X1 port map( A => REGISTERS_24_15_port, ZN => n2038);
   U2134 : INV_X1 port map( A => REGISTERS_30_15_port, ZN => n2102);
   U2135 : INV_X1 port map( A => REGISTERS_4_15_port, ZN => n460);
   U2136 : INV_X1 port map( A => REGISTERS_8_15_port, ZN => n524);
   U2137 : INV_X1 port map( A => REGISTERS_12_15_port, ZN => n1846);
   U2138 : INV_X1 port map( A => REGISTERS_16_16_port, ZN => n1909);
   U2139 : INV_X1 port map( A => REGISTERS_20_16_port, ZN => n1973);
   U2140 : INV_X1 port map( A => REGISTERS_24_16_port, ZN => n2037);
   U2141 : INV_X1 port map( A => REGISTERS_30_16_port, ZN => n2101);
   U2142 : INV_X1 port map( A => REGISTERS_4_16_port, ZN => n459);
   U2143 : INV_X1 port map( A => REGISTERS_8_16_port, ZN => n523);
   U2144 : INV_X1 port map( A => REGISTERS_12_16_port, ZN => n1845);
   U2145 : INV_X1 port map( A => REGISTERS_16_17_port, ZN => n1908);
   U2146 : INV_X1 port map( A => REGISTERS_20_17_port, ZN => n1972);
   U2147 : INV_X1 port map( A => REGISTERS_24_17_port, ZN => n2036);
   U2148 : INV_X1 port map( A => REGISTERS_30_17_port, ZN => n2100);
   U2149 : INV_X1 port map( A => REGISTERS_4_17_port, ZN => n458);
   U2150 : INV_X1 port map( A => REGISTERS_8_17_port, ZN => n522);
   U2151 : INV_X1 port map( A => REGISTERS_12_17_port, ZN => n1844);
   U2152 : INV_X1 port map( A => REGISTERS_16_18_port, ZN => n1907);
   U2153 : INV_X1 port map( A => REGISTERS_20_18_port, ZN => n1971);
   U2154 : INV_X1 port map( A => REGISTERS_24_18_port, ZN => n2035);
   U2155 : INV_X1 port map( A => REGISTERS_30_18_port, ZN => n2099);
   U2156 : INV_X1 port map( A => REGISTERS_4_18_port, ZN => n457);
   U2157 : INV_X1 port map( A => REGISTERS_8_18_port, ZN => n521);
   U2158 : INV_X1 port map( A => REGISTERS_12_18_port, ZN => n1843);
   U2159 : INV_X1 port map( A => REGISTERS_16_19_port, ZN => n1906);
   U2160 : INV_X1 port map( A => REGISTERS_20_19_port, ZN => n1970);
   U2161 : INV_X1 port map( A => REGISTERS_24_19_port, ZN => n2034);
   U2162 : INV_X1 port map( A => REGISTERS_30_19_port, ZN => n2098);
   U2163 : INV_X1 port map( A => REGISTERS_4_19_port, ZN => n456);
   U2164 : INV_X1 port map( A => REGISTERS_8_19_port, ZN => n520);
   U2165 : INV_X1 port map( A => REGISTERS_12_19_port, ZN => n1842);
   U2166 : INV_X1 port map( A => REGISTERS_16_20_port, ZN => n1905);
   U2167 : INV_X1 port map( A => REGISTERS_20_20_port, ZN => n1969);
   U2168 : INV_X1 port map( A => REGISTERS_24_20_port, ZN => n2033);
   U2169 : INV_X1 port map( A => REGISTERS_30_20_port, ZN => n2097);
   U2170 : INV_X1 port map( A => REGISTERS_4_20_port, ZN => n455);
   U2171 : INV_X1 port map( A => REGISTERS_8_20_port, ZN => n519);
   U2172 : INV_X1 port map( A => REGISTERS_12_20_port, ZN => n1841);
   U2173 : INV_X1 port map( A => REGISTERS_16_21_port, ZN => n1904);
   U2174 : INV_X1 port map( A => REGISTERS_20_21_port, ZN => n1968);
   U2175 : INV_X1 port map( A => REGISTERS_24_21_port, ZN => n2032);
   U2176 : INV_X1 port map( A => REGISTERS_30_21_port, ZN => n2096);
   U2177 : INV_X1 port map( A => REGISTERS_4_21_port, ZN => n454);
   U2178 : INV_X1 port map( A => REGISTERS_8_21_port, ZN => n518);
   U2179 : INV_X1 port map( A => REGISTERS_12_21_port, ZN => n1840);
   U2180 : INV_X1 port map( A => REGISTERS_16_22_port, ZN => n1903);
   U2181 : INV_X1 port map( A => REGISTERS_20_22_port, ZN => n1967);
   U2182 : INV_X1 port map( A => REGISTERS_24_22_port, ZN => n2031);
   U2183 : INV_X1 port map( A => REGISTERS_30_22_port, ZN => n2095);
   U2184 : INV_X1 port map( A => REGISTERS_4_22_port, ZN => n453);
   U2185 : INV_X1 port map( A => REGISTERS_8_22_port, ZN => n517);
   U2186 : INV_X1 port map( A => REGISTERS_12_22_port, ZN => n1839);
   U2187 : INV_X1 port map( A => REGISTERS_16_23_port, ZN => n1902);
   U2188 : INV_X1 port map( A => REGISTERS_20_23_port, ZN => n1966);
   U2189 : INV_X1 port map( A => REGISTERS_24_23_port, ZN => n2030);
   U2190 : INV_X1 port map( A => REGISTERS_30_23_port, ZN => n2094);
   U2191 : INV_X1 port map( A => REGISTERS_4_23_port, ZN => n452);
   U2192 : INV_X1 port map( A => REGISTERS_8_23_port, ZN => n516);
   U2193 : INV_X1 port map( A => REGISTERS_12_23_port, ZN => n1838);
   U2194 : INV_X1 port map( A => REGISTERS_16_24_port, ZN => n1901);
   U2195 : INV_X1 port map( A => REGISTERS_20_24_port, ZN => n1965);
   U2196 : INV_X1 port map( A => REGISTERS_24_24_port, ZN => n2029);
   U2197 : INV_X1 port map( A => REGISTERS_30_24_port, ZN => n2093);
   U2198 : INV_X1 port map( A => REGISTERS_4_24_port, ZN => n451);
   U2199 : INV_X1 port map( A => REGISTERS_8_24_port, ZN => n515);
   U2200 : INV_X1 port map( A => REGISTERS_12_24_port, ZN => n1837);
   U2201 : INV_X1 port map( A => REGISTERS_16_25_port, ZN => n1900);
   U2202 : INV_X1 port map( A => REGISTERS_20_25_port, ZN => n1964);
   U2203 : INV_X1 port map( A => REGISTERS_24_25_port, ZN => n2028);
   U2204 : INV_X1 port map( A => REGISTERS_30_25_port, ZN => n2092);
   U2205 : INV_X1 port map( A => REGISTERS_4_25_port, ZN => n450);
   U2206 : INV_X1 port map( A => REGISTERS_8_25_port, ZN => n514);
   U2207 : INV_X1 port map( A => REGISTERS_12_25_port, ZN => n1836);
   U2208 : INV_X1 port map( A => REGISTERS_16_26_port, ZN => n1899);
   U2209 : INV_X1 port map( A => REGISTERS_20_26_port, ZN => n1963);
   U2210 : INV_X1 port map( A => REGISTERS_24_26_port, ZN => n2027);
   U2211 : INV_X1 port map( A => REGISTERS_30_26_port, ZN => n2091);
   U2212 : INV_X1 port map( A => REGISTERS_4_26_port, ZN => n449);
   U2213 : INV_X1 port map( A => REGISTERS_8_26_port, ZN => n513);
   U2214 : INV_X1 port map( A => REGISTERS_12_26_port, ZN => n1835);
   U2215 : INV_X1 port map( A => REGISTERS_16_27_port, ZN => n1898);
   U2216 : INV_X1 port map( A => REGISTERS_20_27_port, ZN => n1962);
   U2217 : INV_X1 port map( A => REGISTERS_24_27_port, ZN => n2026);
   U2218 : INV_X1 port map( A => REGISTERS_30_27_port, ZN => n2090);
   U2219 : INV_X1 port map( A => REGISTERS_4_27_port, ZN => n448);
   U2220 : INV_X1 port map( A => REGISTERS_8_27_port, ZN => n512);
   U2221 : INV_X1 port map( A => REGISTERS_12_27_port, ZN => n1834);
   U2222 : INV_X1 port map( A => REGISTERS_16_28_port, ZN => n1897);
   U2223 : INV_X1 port map( A => REGISTERS_20_28_port, ZN => n1961);
   U2224 : INV_X1 port map( A => REGISTERS_24_28_port, ZN => n2025);
   U2225 : INV_X1 port map( A => REGISTERS_30_28_port, ZN => n2089);
   U2226 : INV_X1 port map( A => REGISTERS_4_28_port, ZN => n447);
   U2227 : INV_X1 port map( A => REGISTERS_8_28_port, ZN => n511);
   U2228 : INV_X1 port map( A => REGISTERS_12_28_port, ZN => n1833);
   U2229 : INV_X1 port map( A => REGISTERS_16_29_port, ZN => n1896);
   U2230 : INV_X1 port map( A => REGISTERS_20_29_port, ZN => n1960);
   U2231 : INV_X1 port map( A => REGISTERS_24_29_port, ZN => n2024);
   U2232 : INV_X1 port map( A => REGISTERS_30_29_port, ZN => n2088);
   U2233 : INV_X1 port map( A => REGISTERS_4_29_port, ZN => n446);
   U2234 : INV_X1 port map( A => REGISTERS_8_29_port, ZN => n510);
   U2235 : INV_X1 port map( A => REGISTERS_12_29_port, ZN => n1832);
   U2236 : INV_X1 port map( A => REGISTERS_16_30_port, ZN => n1895);
   U2237 : INV_X1 port map( A => REGISTERS_20_30_port, ZN => n1959);
   U2238 : INV_X1 port map( A => REGISTERS_24_30_port, ZN => n2023);
   U2239 : INV_X1 port map( A => REGISTERS_30_30_port, ZN => n2087);
   U2240 : INV_X1 port map( A => REGISTERS_4_30_port, ZN => n445);
   U2241 : INV_X1 port map( A => REGISTERS_8_30_port, ZN => n509);
   U2242 : INV_X1 port map( A => REGISTERS_12_30_port, ZN => n1831);
   U2243 : INV_X1 port map( A => REGISTERS_16_31_port, ZN => n1894);
   U2244 : INV_X1 port map( A => REGISTERS_20_31_port, ZN => n1958);
   U2245 : INV_X1 port map( A => REGISTERS_24_31_port, ZN => n2022);
   U2246 : INV_X1 port map( A => REGISTERS_30_31_port, ZN => n2086);
   U2247 : INV_X1 port map( A => REGISTERS_4_31_port, ZN => n444);
   U2248 : INV_X1 port map( A => REGISTERS_8_31_port, ZN => n508);
   U2249 : INV_X1 port map( A => REGISTERS_12_31_port, ZN => n1830);
   U2250 : AND2_X1 port map( A1 => DATAIN(0), A2 => n406, ZN => N244);
   U2251 : AND2_X1 port map( A1 => DATAIN(1), A2 => n406, ZN => N245);
   U2252 : AND2_X1 port map( A1 => DATAIN(2), A2 => n405, ZN => N246);
   U2253 : AND2_X1 port map( A1 => DATAIN(3), A2 => n405, ZN => N247);
   U2254 : AND2_X1 port map( A1 => DATAIN(4), A2 => n405, ZN => N248);
   U2255 : AND2_X1 port map( A1 => DATAIN(5), A2 => n405, ZN => N249);
   U2256 : AND2_X1 port map( A1 => DATAIN(6), A2 => n405, ZN => N250);
   U2257 : AND2_X1 port map( A1 => DATAIN(7), A2 => n405, ZN => N251);
   U2258 : AND2_X1 port map( A1 => DATAIN(8), A2 => n405, ZN => N252);
   U2259 : AND2_X1 port map( A1 => DATAIN(9), A2 => n402, ZN => N253);
   U2260 : AND2_X1 port map( A1 => DATAIN(10), A2 => n404, ZN => N254);
   U2261 : AND2_X1 port map( A1 => DATAIN(11), A2 => n404, ZN => N255);
   U2262 : AND2_X1 port map( A1 => DATAIN(12), A2 => n404, ZN => N256);
   U2263 : AND2_X1 port map( A1 => DATAIN(13), A2 => n404, ZN => N257);
   U2264 : AND2_X1 port map( A1 => DATAIN(14), A2 => n404, ZN => N258);
   U2265 : AND2_X1 port map( A1 => DATAIN(15), A2 => n404, ZN => N259);
   U2266 : AND2_X1 port map( A1 => DATAIN(16), A2 => n404, ZN => N260);
   U2267 : AND2_X1 port map( A1 => DATAIN(17), A2 => n403, ZN => N261);
   U2268 : AND2_X1 port map( A1 => DATAIN(18), A2 => n403, ZN => N262);
   U2269 : AND2_X1 port map( A1 => DATAIN(19), A2 => n403, ZN => N263);
   U2270 : AND2_X1 port map( A1 => DATAIN(20), A2 => n403, ZN => N264);
   U2271 : AND2_X1 port map( A1 => DATAIN(21), A2 => n403, ZN => N265);
   U2272 : AND2_X1 port map( A1 => DATAIN(22), A2 => n403, ZN => N266);
   U2273 : AND2_X1 port map( A1 => DATAIN(23), A2 => n403, ZN => N267);
   U2274 : AND2_X1 port map( A1 => DATAIN(24), A2 => n402, ZN => N268);
   U2275 : AND2_X1 port map( A1 => DATAIN(25), A2 => n402, ZN => N269);
   U2276 : AND2_X1 port map( A1 => DATAIN(26), A2 => n402, ZN => N270);
   U2277 : AND2_X1 port map( A1 => DATAIN(27), A2 => n402, ZN => N271);
   U2278 : AND2_X1 port map( A1 => DATAIN(28), A2 => n402, ZN => N272);
   U2279 : AND2_X1 port map( A1 => DATAIN(29), A2 => n402, ZN => N273);
   U2280 : AND2_X1 port map( A1 => DATAIN(30), A2 => n401, ZN => N274);
   U2281 : AND2_X1 port map( A1 => DATAIN(31), A2 => n401, ZN => N275);
   U2282 : CLKBUF_X1 port map( A => N307, Z => n187);
   U2283 : CLKBUF_X1 port map( A => N307, Z => n188);
   U2284 : CLKBUF_X1 port map( A => N307, Z => n189);
   U2285 : CLKBUF_X1 port map( A => N307, Z => n190);
   U2286 : CLKBUF_X1 port map( A => N307, Z => n191);
   U2287 : CLKBUF_X1 port map( A => N307, Z => n192);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity IR_decoder is

   port( rst : in std_logic;  IR_OUT : in std_logic_vector (20 downto 0);  
         ADDS1, ADDS2, ADDD : out std_logic_vector (4 downto 0));

end IR_decoder;

architecture SYN_Behavioral of IR_decoder is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
      n27, n28, n29, n30, n31, n32, n33, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n34 : std_logic;

begin
   
   U50 : NAND3_X1 port map( A1 => n5, A2 => n4, A3 => n6, ZN => n28);
   U3 : AOI211_X1 port map( C1 => n13, C2 => n14, A => n9, B => n2, ZN => 
                           ADDS2(4));
   U4 : AND2_X1 port map( A1 => n15, A2 => n16, ZN => n13);
   U5 : NOR2_X1 port map( A1 => n17, A2 => n34, ZN => ADDS2(0));
   U6 : NOR2_X1 port map( A1 => n17, A2 => n11, ZN => ADDS2(2));
   U7 : NOR2_X1 port map( A1 => n17, A2 => n12, ZN => ADDS2(1));
   U8 : NOR2_X1 port map( A1 => n17, A2 => n10, ZN => ADDS2(3));
   U9 : OAI21_X1 port map( B1 => n3, B2 => n18, A => n1, ZN => n17);
   U10 : NAND2_X1 port map( A1 => n16, A2 => n15, ZN => n18);
   U11 : INV_X1 port map( A => n14, ZN => n3);
   U12 : NOR2_X1 port map( A1 => n16, A2 => n2, ZN => n23);
   U13 : NAND2_X1 port map( A1 => n1, A2 => n19, ZN => n22);
   U14 : INV_X1 port map( A => rst, ZN => n2);
   U15 : NAND4_X1 port map( A1 => IR_OUT(20), A2 => IR_OUT(18), A3 => n30, A4 
                           => n31, ZN => n15);
   U16 : NOR2_X1 port map( A1 => IR_OUT(19), A2 => IR_OUT(17), ZN => n30);
   U17 : NOR3_X1 port map( A1 => n28, A2 => n7, A3 => n8, ZN => n19);
   U18 : INV_X1 port map( A => IR_OUT(16), ZN => n7);
   U19 : NAND2_X1 port map( A1 => IR_OUT(16), A2 => n8, ZN => n31);
   U20 : NAND2_X1 port map( A1 => IR_OUT(19), A2 => n19, ZN => n14);
   U21 : INV_X1 port map( A => IR_OUT(17), ZN => n6);
   U22 : INV_X1 port map( A => IR_OUT(18), ZN => n5);
   U23 : OR4_X1 port map( A1 => n28, A2 => IR_OUT(15), A3 => IR_OUT(16), A4 => 
                           IR_OUT(19), ZN => n16);
   U24 : INV_X1 port map( A => IR_OUT(20), ZN => n4);
   U25 : AND2_X1 port map( A1 => IR_OUT(10), A2 => n1, ZN => ADDS1(0));
   U26 : AND2_X1 port map( A1 => IR_OUT(14), A2 => n1, ZN => ADDS1(4));
   U27 : AND2_X1 port map( A1 => IR_OUT(12), A2 => n1, ZN => ADDS1(2));
   U28 : AND2_X1 port map( A1 => IR_OUT(11), A2 => n1, ZN => ADDS1(1));
   U29 : INV_X1 port map( A => IR_OUT(15), ZN => n8);
   U30 : AND2_X1 port map( A1 => IR_OUT(13), A2 => n1, ZN => ADDS1(3));
   U31 : INV_X1 port map( A => IR_OUT(5), ZN => n34);
   U32 : INV_X1 port map( A => IR_OUT(6), ZN => n12);
   U33 : INV_X1 port map( A => IR_OUT(7), ZN => n11);
   U34 : INV_X1 port map( A => IR_OUT(8), ZN => n10);
   U35 : INV_X1 port map( A => IR_OUT(9), ZN => n9);
   U36 : NAND4_X1 port map( A1 => n1, A2 => n16, A3 => n29, A4 => n15, ZN => 
                           n20);
   U37 : OAI211_X1 port map( C1 => n32, C2 => n33, A => n5, B => n4, ZN => n29)
                           ;
   U38 : NOR2_X1 port map( A1 => IR_OUT(17), A2 => n31, ZN => n33);
   U39 : NOR3_X1 port map( A1 => n6, A2 => IR_OUT(19), A3 => IR_OUT(16), ZN => 
                           n32);
   U40 : OAI211_X1 port map( C1 => n34, C2 => n20, A => n27, B => n22, ZN => 
                           ADDD(0));
   U41 : NAND2_X1 port map( A1 => IR_OUT(0), A2 => n23, ZN => n27);
   U42 : OAI211_X1 port map( C1 => n12, C2 => n20, A => n26, B => n22, ZN => 
                           ADDD(1));
   U43 : NAND2_X1 port map( A1 => IR_OUT(1), A2 => n23, ZN => n26);
   U44 : OAI211_X1 port map( C1 => n11, C2 => n20, A => n25, B => n22, ZN => 
                           ADDD(2));
   U45 : NAND2_X1 port map( A1 => IR_OUT(2), A2 => n23, ZN => n25);
   U46 : OAI211_X1 port map( C1 => n10, C2 => n20, A => n24, B => n22, ZN => 
                           ADDD(3));
   U47 : NAND2_X1 port map( A1 => IR_OUT(3), A2 => n23, ZN => n24);
   U48 : OAI211_X1 port map( C1 => n9, C2 => n20, A => n21, B => n22, ZN => 
                           ADDD(4));
   U49 : NAND2_X1 port map( A1 => IR_OUT(4), A2 => n23, ZN => n21);
   U51 : INV_X1 port map( A => n2, ZN => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity IF_ID is

   port( CLK, RST, DISCARD : in std_logic;  NPC_IN, NPC_L_IN, IR_IN : in 
         std_logic_vector (31 downto 0);  PR_IN : in std_logic;  NPC_OUT, 
         NPC_L_OUT, IR_OUT : out std_logic_vector (31 downto 0);  PR_OUT : out 
         std_logic);

end IF_ID;

architecture SYN_Behavioral of IF_ID is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_IF_ID
      port( CLK, EN : in std_logic;  ENCLK : out std_logic;  TE : in std_logic
            );
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net1013, net1014, n99, n101, n103, n105, n107, n109, n111, n113, n115
      , n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, n137, n139,
      n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, n161, n163, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n100, n102, n104, n106, 
      n108, n110, n112, n114, n116, n118, n120, n122, n124, n126, n128, n130, 
      n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, 
      n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, 
      n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, 
      n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, 
      n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, 
      n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, 
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, 
      n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717 : std_logic;

begin
   
   net1014 <= '0';
   PR_OUT_reg : DFFR_X1 port map( D => PR_IN, CK => net1013, RN => n47, Q => 
                           PR_OUT, QN => n_1621);
   IR_OUT_reg_31_inst : DFFR_X1 port map( D => IR_IN(31), CK => CLK, RN => n35,
                           Q => IR_OUT(31), QN => n_1622);
   IR_OUT_reg_30_inst : DFFS_X1 port map( D => IR_IN(30), CK => CLK, SN => n36,
                           Q => IR_OUT(30), QN => n_1623);
   IR_OUT_reg_29_inst : DFFR_X1 port map( D => IR_IN(29), CK => CLK, RN => n34,
                           Q => IR_OUT(29), QN => n_1624);
   IR_OUT_reg_28_inst : DFFS_X1 port map( D => IR_IN(28), CK => CLK, SN => n36,
                           Q => IR_OUT(28), QN => n_1625);
   IR_OUT_reg_27_inst : DFFR_X1 port map( D => IR_IN(27), CK => CLK, RN => n34,
                           Q => IR_OUT(27), QN => n_1626);
   IR_OUT_reg_26_inst : DFFS_X1 port map( D => IR_IN(26), CK => CLK, SN => n36,
                           Q => IR_OUT(26), QN => n_1627);
   IR_OUT_reg_25_inst : DFFR_X1 port map( D => IR_IN(25), CK => CLK, RN => n34,
                           Q => IR_OUT(25), QN => n_1628);
   IR_OUT_reg_24_inst : DFFR_X1 port map( D => IR_IN(24), CK => CLK, RN => n34,
                           Q => IR_OUT(24), QN => n_1629);
   IR_OUT_reg_23_inst : DFFR_X1 port map( D => IR_IN(23), CK => CLK, RN => n34,
                           Q => IR_OUT(23), QN => n_1630);
   IR_OUT_reg_22_inst : DFFR_X1 port map( D => IR_IN(22), CK => CLK, RN => n34,
                           Q => IR_OUT(22), QN => n_1631);
   IR_OUT_reg_21_inst : DFFR_X1 port map( D => IR_IN(21), CK => CLK, RN => n34,
                           Q => IR_OUT(21), QN => n_1632);
   IR_OUT_reg_20_inst : DFFR_X1 port map( D => IR_IN(20), CK => CLK, RN => n34,
                           Q => IR_OUT(20), QN => n_1633);
   IR_OUT_reg_19_inst : DFFR_X1 port map( D => IR_IN(19), CK => CLK, RN => n34,
                           Q => IR_OUT(19), QN => n_1634);
   IR_OUT_reg_18_inst : DFFR_X1 port map( D => IR_IN(18), CK => CLK, RN => n34,
                           Q => IR_OUT(18), QN => n_1635);
   IR_OUT_reg_17_inst : DFFR_X1 port map( D => IR_IN(17), CK => CLK, RN => n34,
                           Q => IR_OUT(17), QN => n_1636);
   IR_OUT_reg_16_inst : DFFR_X1 port map( D => IR_IN(16), CK => CLK, RN => n35,
                           Q => IR_OUT(16), QN => n_1637);
   IR_OUT_reg_15_inst : DFFR_X1 port map( D => IR_IN(15), CK => CLK, RN => n35,
                           Q => IR_OUT(15), QN => n_1638);
   IR_OUT_reg_14_inst : DFFR_X1 port map( D => IR_IN(14), CK => CLK, RN => n35,
                           Q => IR_OUT(14), QN => n_1639);
   IR_OUT_reg_13_inst : DFFR_X1 port map( D => IR_IN(13), CK => CLK, RN => n35,
                           Q => IR_OUT(13), QN => n_1640);
   IR_OUT_reg_12_inst : DFFR_X1 port map( D => IR_IN(12), CK => CLK, RN => n35,
                           Q => IR_OUT(12), QN => n_1641);
   IR_OUT_reg_11_inst : DFFR_X1 port map( D => IR_IN(11), CK => CLK, RN => n35,
                           Q => IR_OUT(11), QN => n_1642);
   IR_OUT_reg_10_inst : DFFR_X1 port map( D => IR_IN(10), CK => CLK, RN => n35,
                           Q => IR_OUT(10), QN => n_1643);
   IR_OUT_reg_9_inst : DFFR_X1 port map( D => IR_IN(9), CK => CLK, RN => n35, Q
                           => IR_OUT(9), QN => n_1644);
   IR_OUT_reg_8_inst : DFFR_X1 port map( D => IR_IN(8), CK => CLK, RN => n35, Q
                           => IR_OUT(8), QN => n_1645);
   IR_OUT_reg_7_inst : DFFR_X1 port map( D => IR_IN(7), CK => CLK, RN => n35, Q
                           => IR_OUT(7), QN => n_1646);
   IR_OUT_reg_6_inst : DFFR_X1 port map( D => IR_IN(6), CK => CLK, RN => n35, Q
                           => IR_OUT(6), QN => n_1647);
   IR_OUT_reg_5_inst : DFFR_X1 port map( D => IR_IN(5), CK => CLK, RN => n36, Q
                           => IR_OUT(5), QN => n_1648);
   IR_OUT_reg_4_inst : DFFR_X1 port map( D => IR_IN(4), CK => CLK, RN => n36, Q
                           => IR_OUT(4), QN => n_1649);
   IR_OUT_reg_3_inst : DFFR_X1 port map( D => IR_IN(3), CK => CLK, RN => n36, Q
                           => IR_OUT(3), QN => n_1650);
   IR_OUT_reg_2_inst : DFFR_X1 port map( D => IR_IN(2), CK => CLK, RN => n36, Q
                           => IR_OUT(2), QN => n_1651);
   IR_OUT_reg_1_inst : DFFR_X1 port map( D => IR_IN(1), CK => CLK, RN => n36, Q
                           => IR_OUT(1), QN => n_1652);
   IR_OUT_reg_0_inst : DFFR_X1 port map( D => IR_IN(0), CK => CLK, RN => n34, Q
                           => IR_OUT(0), QN => n_1653);
   NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => NPC_L_IN(31), CK => net1013, 
                           RN => n47, Q => NPC_L_OUT(31), QN => n_1654);
   NPC_L_OUT_reg_30_inst : DFFR_X1 port map( D => NPC_L_IN(30), CK => net1013, 
                           RN => n47, Q => NPC_L_OUT(30), QN => n_1655);
   NPC_L_OUT_reg_29_inst : DFFR_X1 port map( D => NPC_L_IN(29), CK => net1013, 
                           RN => n47, Q => NPC_L_OUT(29), QN => n_1656);
   NPC_L_OUT_reg_28_inst : DFFR_X1 port map( D => NPC_L_IN(28), CK => net1013, 
                           RN => n47, Q => NPC_L_OUT(28), QN => n_1657);
   NPC_L_OUT_reg_27_inst : DFFR_X1 port map( D => NPC_L_IN(27), CK => net1013, 
                           RN => n47, Q => NPC_L_OUT(27), QN => n_1658);
   NPC_L_OUT_reg_26_inst : DFFR_X1 port map( D => NPC_L_IN(26), CK => net1013, 
                           RN => n47, Q => NPC_L_OUT(26), QN => n_1659);
   NPC_L_OUT_reg_25_inst : DFFR_X1 port map( D => NPC_L_IN(25), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(25), QN => n_1660);
   NPC_L_OUT_reg_24_inst : DFFR_X1 port map( D => NPC_L_IN(24), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(24), QN => n_1661);
   NPC_L_OUT_reg_23_inst : DFFR_X1 port map( D => NPC_L_IN(23), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(23), QN => n_1662);
   NPC_L_OUT_reg_22_inst : DFFR_X1 port map( D => NPC_L_IN(22), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(22), QN => n_1663);
   NPC_L_OUT_reg_21_inst : DFFR_X1 port map( D => NPC_L_IN(21), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(21), QN => n_1664);
   NPC_L_OUT_reg_20_inst : DFFR_X1 port map( D => NPC_L_IN(20), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(20), QN => n_1665);
   NPC_L_OUT_reg_19_inst : DFFR_X1 port map( D => NPC_L_IN(19), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(19), QN => n_1666);
   NPC_L_OUT_reg_18_inst : DFFR_X1 port map( D => NPC_L_IN(18), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(18), QN => n_1667);
   NPC_L_OUT_reg_17_inst : DFFR_X1 port map( D => NPC_L_IN(17), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(17), QN => n_1668);
   NPC_L_OUT_reg_16_inst : DFFR_X1 port map( D => NPC_L_IN(16), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(16), QN => n_1669);
   NPC_L_OUT_reg_15_inst : DFFR_X1 port map( D => NPC_L_IN(15), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(15), QN => n_1670);
   NPC_L_OUT_reg_14_inst : DFFR_X1 port map( D => NPC_L_IN(14), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(14), QN => n_1671);
   NPC_L_OUT_reg_13_inst : DFFR_X1 port map( D => NPC_L_IN(13), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(13), QN => n_1672);
   NPC_L_OUT_reg_12_inst : DFFR_X1 port map( D => NPC_L_IN(12), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(12), QN => n_1673);
   NPC_L_OUT_reg_11_inst : DFFR_X1 port map( D => NPC_L_IN(11), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(11), QN => n_1674);
   NPC_L_OUT_reg_10_inst : DFFR_X1 port map( D => NPC_L_IN(10), CK => net1013, 
                           RN => n48, Q => NPC_L_OUT(10), QN => n_1675);
   NPC_L_OUT_reg_9_inst : DFFR_X1 port map( D => NPC_L_IN(9), CK => net1013, RN
                           => n48, Q => NPC_L_OUT(9), QN => n_1676);
   NPC_L_OUT_reg_8_inst : DFFR_X1 port map( D => NPC_L_IN(8), CK => net1013, RN
                           => n48, Q => NPC_L_OUT(8), QN => n_1677);
   NPC_L_OUT_reg_7_inst : DFFR_X1 port map( D => NPC_L_IN(7), CK => net1013, RN
                           => n48, Q => NPC_L_OUT(7), QN => n_1678);
   NPC_L_OUT_reg_6_inst : DFFR_X1 port map( D => NPC_L_IN(6), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(6), QN => n_1679);
   NPC_L_OUT_reg_5_inst : DFFR_X1 port map( D => NPC_L_IN(5), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(5), QN => n_1680);
   NPC_L_OUT_reg_4_inst : DFFR_X1 port map( D => NPC_L_IN(4), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(4), QN => n_1681);
   NPC_L_OUT_reg_3_inst : DFFR_X1 port map( D => NPC_L_IN(3), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(3), QN => n_1682);
   NPC_L_OUT_reg_2_inst : DFFR_X1 port map( D => NPC_L_IN(2), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(2), QN => n_1683);
   NPC_L_OUT_reg_1_inst : DFFR_X1 port map( D => NPC_L_IN(1), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(1), QN => n_1684);
   NPC_L_OUT_reg_0_inst : DFFR_X1 port map( D => NPC_L_IN(0), CK => net1013, RN
                           => n49, Q => NPC_L_OUT(0), QN => n_1685);
   clk_gate_PR_OUT_reg : SNPS_CLOCK_GATE_HIGH_IF_ID port map( CLK => CLK, EN =>
                           n39, ENCLK => net1013, TE => net1014);
   NPC_OUT_reg_31_inst : DFFRS_X1 port map( D => NPC_IN(31), CK => CLK, RN => 
                           n73, SN => n25, Q => NPC_OUT(31), QN => n_1686);
   NPC_OUT_reg_30_inst : DFFRS_X1 port map( D => NPC_IN(30), CK => CLK, RN => 
                           n72, SN => n24, Q => NPC_OUT(30), QN => n_1687);
   NPC_OUT_reg_29_inst : DFFRS_X1 port map( D => NPC_IN(29), CK => CLK, RN => 
                           n71, SN => n23, Q => NPC_OUT(29), QN => n_1688);
   NPC_OUT_reg_28_inst : DFFRS_X1 port map( D => NPC_IN(28), CK => CLK, RN => 
                           n70, SN => n22, Q => NPC_OUT(28), QN => n_1689);
   NPC_OUT_reg_27_inst : DFFRS_X1 port map( D => NPC_IN(27), CK => CLK, RN => 
                           n69, SN => n21, Q => NPC_OUT(27), QN => n_1690);
   NPC_OUT_reg_26_inst : DFFRS_X1 port map( D => NPC_IN(26), CK => CLK, RN => 
                           n68, SN => n20, Q => NPC_OUT(26), QN => n_1691);
   NPC_OUT_reg_25_inst : DFFRS_X1 port map( D => NPC_IN(25), CK => CLK, RN => 
                           n67, SN => n19, Q => NPC_OUT(25), QN => n_1692);
   NPC_OUT_reg_24_inst : DFFRS_X1 port map( D => NPC_IN(24), CK => CLK, RN => 
                           n66, SN => n18, Q => NPC_OUT(24), QN => n_1693);
   NPC_OUT_reg_23_inst : DFFRS_X1 port map( D => NPC_IN(23), CK => CLK, RN => 
                           n65, SN => n17, Q => NPC_OUT(23), QN => n_1694);
   NPC_OUT_reg_22_inst : DFFRS_X1 port map( D => NPC_IN(22), CK => CLK, RN => 
                           n64, SN => n16, Q => NPC_OUT(22), QN => n_1695);
   NPC_OUT_reg_21_inst : DFFRS_X1 port map( D => NPC_IN(21), CK => CLK, RN => 
                           n63, SN => n15, Q => NPC_OUT(21), QN => n_1696);
   NPC_OUT_reg_20_inst : DFFRS_X1 port map( D => NPC_IN(20), CK => CLK, RN => 
                           n62, SN => n14, Q => NPC_OUT(20), QN => n_1697);
   NPC_OUT_reg_19_inst : DFFRS_X1 port map( D => NPC_IN(19), CK => CLK, RN => 
                           n61, SN => n13, Q => NPC_OUT(19), QN => n_1698);
   NPC_OUT_reg_18_inst : DFFRS_X1 port map( D => NPC_IN(18), CK => CLK, RN => 
                           n60, SN => n12, Q => NPC_OUT(18), QN => n_1699);
   NPC_OUT_reg_17_inst : DFFRS_X1 port map( D => NPC_IN(17), CK => CLK, RN => 
                           n59, SN => n11, Q => NPC_OUT(17), QN => n_1700);
   NPC_OUT_reg_16_inst : DFFRS_X1 port map( D => NPC_IN(16), CK => CLK, RN => 
                           n58, SN => n33, Q => NPC_OUT(16), QN => n_1701);
   NPC_OUT_reg_15_inst : DFFRS_X1 port map( D => NPC_IN(15), CK => CLK, RN => 
                           n57, SN => n32, Q => NPC_OUT(15), QN => n_1702);
   NPC_OUT_reg_14_inst : DFFRS_X1 port map( D => NPC_IN(14), CK => CLK, RN => 
                           n56, SN => n31, Q => NPC_OUT(14), QN => n_1703);
   NPC_OUT_reg_13_inst : DFFRS_X1 port map( D => NPC_IN(13), CK => CLK, RN => 
                           n55, SN => n30, Q => NPC_OUT(13), QN => n_1704);
   NPC_OUT_reg_12_inst : DFFRS_X1 port map( D => NPC_IN(12), CK => CLK, RN => 
                           n54, SN => n29, Q => NPC_OUT(12), QN => n_1705);
   NPC_OUT_reg_11_inst : DFFRS_X1 port map( D => NPC_IN(11), CK => CLK, RN => 
                           n53, SN => n28, Q => NPC_OUT(11), QN => n_1706);
   NPC_OUT_reg_10_inst : DFFRS_X1 port map( D => NPC_IN(10), CK => CLK, RN => 
                           n52, SN => n27, Q => NPC_OUT(10), QN => n_1707);
   NPC_OUT_reg_9_inst : DFFRS_X1 port map( D => NPC_IN(9), CK => CLK, RN => n51
                           , SN => n26, Q => NPC_OUT(9), QN => n_1708);
   NPC_OUT_reg_8_inst : DFFRS_X1 port map( D => NPC_IN(8), CK => CLK, RN => n50
                           , SN => n10, Q => NPC_OUT(8), QN => n_1709);
   NPC_OUT_reg_7_inst : DFFRS_X1 port map( D => NPC_IN(7), CK => CLK, RN => n81
                           , SN => n9, Q => NPC_OUT(7), QN => n_1710);
   NPC_OUT_reg_6_inst : DFFRS_X1 port map( D => NPC_IN(6), CK => CLK, RN => n80
                           , SN => n8, Q => NPC_OUT(6), QN => n_1711);
   NPC_OUT_reg_5_inst : DFFRS_X1 port map( D => NPC_IN(5), CK => CLK, RN => n79
                           , SN => n7, Q => NPC_OUT(5), QN => n_1712);
   NPC_OUT_reg_4_inst : DFFRS_X1 port map( D => NPC_IN(4), CK => CLK, RN => n78
                           , SN => n6, Q => NPC_OUT(4), QN => n_1713);
   NPC_OUT_reg_3_inst : DFFRS_X1 port map( D => NPC_IN(3), CK => CLK, RN => n77
                           , SN => n5, Q => NPC_OUT(3), QN => n_1714);
   NPC_OUT_reg_2_inst : DFFRS_X1 port map( D => NPC_IN(2), CK => CLK, RN => n76
                           , SN => n4, Q => NPC_OUT(2), QN => n_1715);
   NPC_OUT_reg_1_inst : DFFRS_X1 port map( D => NPC_IN(1), CK => CLK, RN => n75
                           , SN => n3, Q => NPC_OUT(1), QN => n_1716);
   NPC_OUT_reg_0_inst : DFFRS_X1 port map( D => NPC_IN(0), CK => CLK, RN => n74
                           , SN => n2, Q => NPC_OUT(0), QN => n_1717);
   U3 : INV_X1 port map( A => NPC_IN(0), ZN => n130);
   U4 : INV_X1 port map( A => NPC_IN(1), ZN => n128);
   U5 : INV_X1 port map( A => NPC_IN(2), ZN => n126);
   U6 : INV_X1 port map( A => NPC_IN(3), ZN => n124);
   U7 : INV_X1 port map( A => NPC_IN(4), ZN => n122);
   U8 : INV_X1 port map( A => NPC_IN(5), ZN => n120);
   U9 : INV_X1 port map( A => NPC_IN(6), ZN => n118);
   U10 : INV_X1 port map( A => NPC_IN(7), ZN => n116);
   U11 : INV_X1 port map( A => NPC_IN(8), ZN => n114);
   U12 : INV_X1 port map( A => NPC_IN(9), ZN => n112);
   U13 : INV_X1 port map( A => NPC_IN(10), ZN => n110);
   U14 : INV_X1 port map( A => NPC_IN(11), ZN => n108);
   U15 : INV_X1 port map( A => NPC_IN(12), ZN => n106);
   U16 : INV_X1 port map( A => NPC_IN(13), ZN => n104);
   U17 : INV_X1 port map( A => NPC_IN(14), ZN => n102);
   U18 : INV_X1 port map( A => NPC_IN(15), ZN => n100);
   U19 : INV_X1 port map( A => NPC_IN(16), ZN => n98);
   U20 : INV_X1 port map( A => NPC_IN(17), ZN => n97);
   U21 : INV_X1 port map( A => NPC_IN(18), ZN => n96);
   U22 : INV_X1 port map( A => NPC_IN(19), ZN => n95);
   U23 : INV_X1 port map( A => NPC_IN(20), ZN => n94);
   U24 : INV_X1 port map( A => NPC_IN(21), ZN => n93);
   U25 : INV_X1 port map( A => NPC_IN(22), ZN => n92);
   U26 : INV_X1 port map( A => NPC_IN(23), ZN => n91);
   U27 : INV_X1 port map( A => NPC_IN(24), ZN => n90);
   U28 : INV_X1 port map( A => NPC_IN(25), ZN => n89);
   U29 : INV_X1 port map( A => NPC_IN(26), ZN => n88);
   U30 : INV_X1 port map( A => NPC_IN(27), ZN => n87);
   U31 : INV_X1 port map( A => NPC_IN(28), ZN => n86);
   U32 : INV_X1 port map( A => NPC_IN(29), ZN => n85);
   U33 : INV_X1 port map( A => NPC_IN(30), ZN => n84);
   U34 : INV_X1 port map( A => NPC_IN(31), ZN => n83);
   U35 : BUF_X1 port map( A => n1, Z => n34);
   U36 : BUF_X1 port map( A => n1, Z => n35);
   U37 : BUF_X1 port map( A => n1, Z => n36);
   U38 : BUF_X1 port map( A => n82, Z => n39);
   U39 : BUF_X1 port map( A => n82, Z => n37);
   U40 : BUF_X1 port map( A => n82, Z => n38);
   U41 : BUF_X1 port map( A => n99, Z => n41);
   U42 : BUF_X1 port map( A => n99, Z => n40);
   U43 : BUF_X1 port map( A => n99, Z => n42);
   U44 : AND2_X1 port map( A1 => n47, A2 => n37, ZN => n1);
   U45 : INV_X1 port map( A => DISCARD, ZN => n82);
   U46 : BUF_X1 port map( A => n44, Z => n48);
   U47 : BUF_X1 port map( A => n43, Z => n45);
   U48 : BUF_X1 port map( A => n43, Z => n46);
   U49 : BUF_X1 port map( A => n43, Z => n47);
   U50 : NAND2_X1 port map( A1 => DISCARD, A2 => n45, ZN => n99);
   U51 : BUF_X1 port map( A => n44, Z => n49);
   U52 : BUF_X1 port map( A => RST, Z => n43);
   U53 : BUF_X1 port map( A => RST, Z => n44);
   U54 : INV_X1 port map( A => n101, ZN => n74);
   U55 : OAI21_X1 port map( B1 => NPC_IN(0), B2 => n39, A => n46, ZN => n101);
   U56 : INV_X1 port map( A => n103, ZN => n75);
   U57 : OAI21_X1 port map( B1 => NPC_IN(1), B2 => n39, A => n46, ZN => n103);
   U58 : INV_X1 port map( A => n105, ZN => n76);
   U59 : OAI21_X1 port map( B1 => NPC_IN(2), B2 => n39, A => n47, ZN => n105);
   U60 : INV_X1 port map( A => n107, ZN => n77);
   U61 : OAI21_X1 port map( B1 => NPC_IN(3), B2 => n39, A => n47, ZN => n107);
   U62 : INV_X1 port map( A => n109, ZN => n78);
   U63 : OAI21_X1 port map( B1 => NPC_IN(4), B2 => n39, A => n47, ZN => n109);
   U64 : INV_X1 port map( A => n111, ZN => n79);
   U65 : OAI21_X1 port map( B1 => NPC_IN(5), B2 => n39, A => n47, ZN => n111);
   U66 : INV_X1 port map( A => n113, ZN => n80);
   U67 : OAI21_X1 port map( B1 => NPC_IN(6), B2 => n39, A => n47, ZN => n113);
   U68 : INV_X1 port map( A => n115, ZN => n81);
   U69 : OAI21_X1 port map( B1 => NPC_IN(7), B2 => n39, A => n47, ZN => n115);
   U70 : INV_X1 port map( A => n163, ZN => n73);
   U71 : OAI21_X1 port map( B1 => NPC_IN(31), B2 => n39, A => n46, ZN => n163);
   U72 : INV_X1 port map( A => n119, ZN => n51);
   U73 : OAI21_X1 port map( B1 => NPC_IN(9), B2 => n37, A => n45, ZN => n119);
   U74 : INV_X1 port map( A => n121, ZN => n52);
   U75 : OAI21_X1 port map( B1 => NPC_IN(10), B2 => n37, A => n45, ZN => n121);
   U76 : INV_X1 port map( A => n123, ZN => n53);
   U77 : OAI21_X1 port map( B1 => NPC_IN(11), B2 => n37, A => n45, ZN => n123);
   U78 : INV_X1 port map( A => n125, ZN => n54);
   U79 : OAI21_X1 port map( B1 => NPC_IN(12), B2 => n37, A => n45, ZN => n125);
   U80 : INV_X1 port map( A => n127, ZN => n55);
   U81 : OAI21_X1 port map( B1 => NPC_IN(13), B2 => n37, A => n45, ZN => n127);
   U82 : INV_X1 port map( A => n129, ZN => n56);
   U83 : OAI21_X1 port map( B1 => NPC_IN(14), B2 => n37, A => n45, ZN => n129);
   U84 : INV_X1 port map( A => n131, ZN => n57);
   U85 : OAI21_X1 port map( B1 => NPC_IN(15), B2 => n37, A => n45, ZN => n131);
   U86 : INV_X1 port map( A => n133, ZN => n58);
   U87 : OAI21_X1 port map( B1 => NPC_IN(16), B2 => n37, A => n45, ZN => n133);
   U88 : INV_X1 port map( A => n135, ZN => n59);
   U89 : OAI21_X1 port map( B1 => NPC_IN(17), B2 => n37, A => n45, ZN => n135);
   U90 : INV_X1 port map( A => n137, ZN => n60);
   U91 : OAI21_X1 port map( B1 => NPC_IN(18), B2 => n37, A => n45, ZN => n137);
   U92 : INV_X1 port map( A => n139, ZN => n61);
   U93 : OAI21_X1 port map( B1 => NPC_IN(19), B2 => n37, A => n45, ZN => n139);
   U94 : INV_X1 port map( A => n117, ZN => n50);
   U95 : OAI21_X1 port map( B1 => NPC_IN(8), B2 => n38, A => n47, ZN => n117);
   U96 : INV_X1 port map( A => n141, ZN => n62);
   U97 : OAI21_X1 port map( B1 => NPC_IN(20), B2 => n38, A => n45, ZN => n141);
   U98 : INV_X1 port map( A => n143, ZN => n63);
   U99 : OAI21_X1 port map( B1 => NPC_IN(21), B2 => n38, A => n46, ZN => n143);
   U100 : INV_X1 port map( A => n145, ZN => n64);
   U101 : OAI21_X1 port map( B1 => NPC_IN(22), B2 => n38, A => n46, ZN => n145)
                           ;
   U102 : INV_X1 port map( A => n147, ZN => n65);
   U103 : OAI21_X1 port map( B1 => NPC_IN(23), B2 => n38, A => n46, ZN => n147)
                           ;
   U104 : INV_X1 port map( A => n149, ZN => n66);
   U105 : OAI21_X1 port map( B1 => NPC_IN(24), B2 => n38, A => n46, ZN => n149)
                           ;
   U106 : INV_X1 port map( A => n151, ZN => n67);
   U107 : OAI21_X1 port map( B1 => NPC_IN(25), B2 => n38, A => n46, ZN => n151)
                           ;
   U108 : INV_X1 port map( A => n153, ZN => n68);
   U109 : OAI21_X1 port map( B1 => NPC_IN(26), B2 => n38, A => n46, ZN => n153)
                           ;
   U110 : INV_X1 port map( A => n155, ZN => n69);
   U111 : OAI21_X1 port map( B1 => NPC_IN(27), B2 => n38, A => n46, ZN => n155)
                           ;
   U112 : INV_X1 port map( A => n157, ZN => n70);
   U113 : OAI21_X1 port map( B1 => NPC_IN(28), B2 => n38, A => n46, ZN => n157)
                           ;
   U114 : INV_X1 port map( A => n159, ZN => n71);
   U115 : OAI21_X1 port map( B1 => NPC_IN(29), B2 => n38, A => n46, ZN => n159)
                           ;
   U116 : INV_X1 port map( A => n161, ZN => n72);
   U117 : OAI21_X1 port map( B1 => NPC_IN(30), B2 => n38, A => n46, ZN => n161)
                           ;
   U118 : OR2_X1 port map( A1 => n40, A2 => n130, ZN => n2);
   U119 : OR2_X1 port map( A1 => n40, A2 => n128, ZN => n3);
   U120 : OR2_X1 port map( A1 => n40, A2 => n126, ZN => n4);
   U121 : OR2_X1 port map( A1 => n40, A2 => n124, ZN => n5);
   U122 : OR2_X1 port map( A1 => n40, A2 => n122, ZN => n6);
   U123 : OR2_X1 port map( A1 => n40, A2 => n120, ZN => n7);
   U124 : OR2_X1 port map( A1 => n40, A2 => n118, ZN => n8);
   U125 : OR2_X1 port map( A1 => n40, A2 => n116, ZN => n9);
   U126 : OR2_X1 port map( A1 => n40, A2 => n114, ZN => n10);
   U127 : OR2_X1 port map( A1 => n41, A2 => n97, ZN => n11);
   U128 : OR2_X1 port map( A1 => n41, A2 => n96, ZN => n12);
   U129 : OR2_X1 port map( A1 => n41, A2 => n95, ZN => n13);
   U130 : OR2_X1 port map( A1 => n41, A2 => n94, ZN => n14);
   U131 : OR2_X1 port map( A1 => n41, A2 => n93, ZN => n15);
   U132 : OR2_X1 port map( A1 => n41, A2 => n92, ZN => n16);
   U133 : OR2_X1 port map( A1 => n41, A2 => n91, ZN => n17);
   U134 : OR2_X1 port map( A1 => n41, A2 => n90, ZN => n18);
   U135 : OR2_X1 port map( A1 => n41, A2 => n89, ZN => n19);
   U136 : OR2_X1 port map( A1 => n41, A2 => n88, ZN => n20);
   U137 : OR2_X1 port map( A1 => n41, A2 => n87, ZN => n21);
   U138 : OR2_X1 port map( A1 => n41, A2 => n86, ZN => n22);
   U139 : OR2_X1 port map( A1 => n40, A2 => n85, ZN => n23);
   U140 : OR2_X1 port map( A1 => n40, A2 => n84, ZN => n24);
   U141 : OR2_X1 port map( A1 => n40, A2 => n83, ZN => n25);
   U142 : OR2_X1 port map( A1 => n42, A2 => n112, ZN => n26);
   U143 : OR2_X1 port map( A1 => n42, A2 => n110, ZN => n27);
   U144 : OR2_X1 port map( A1 => n42, A2 => n108, ZN => n28);
   U145 : OR2_X1 port map( A1 => n42, A2 => n106, ZN => n29);
   U146 : OR2_X1 port map( A1 => n42, A2 => n104, ZN => n30);
   U147 : OR2_X1 port map( A1 => n42, A2 => n102, ZN => n31);
   U148 : OR2_X1 port map( A1 => n42, A2 => n100, ZN => n32);
   U149 : OR2_X1 port map( A1 => n42, A2 => n98, ZN => n33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity NPC_adder is

   port( inPC : in std_logic_vector (31 downto 0);  outPC : out 
         std_logic_vector (31 downto 0));

end NPC_adder;

architecture SYN_Behavioral of NPC_adder is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NPC_adder_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, N0, N1, N2, N3, N4, N5, N6, N7, N8, N9,
      N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24
      , N25, N26, N27, N28, N29, N30, N31, N32, n1_port, n2_port, n3_port, 
      n4_port, n5_port, n6_port, n7_port, n8_port, n9_port, n10_port, n11_port,
      n12_port, n13_port, n14_port, n15_port, n16_port, n17_port, n_1718 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   outPC_reg_31_inst : DLH_X1 port map( G => n4_port, D => N32, Q => outPC(31))
                           ;
   outPC_reg_30_inst : DLH_X1 port map( G => n4_port, D => N31, Q => outPC(30))
                           ;
   outPC_reg_29_inst : DLH_X1 port map( G => n4_port, D => N30, Q => outPC(29))
                           ;
   outPC_reg_28_inst : DLH_X1 port map( G => n4_port, D => N29, Q => outPC(28))
                           ;
   outPC_reg_27_inst : DLH_X1 port map( G => n4_port, D => N28, Q => outPC(27))
                           ;
   outPC_reg_26_inst : DLH_X1 port map( G => n4_port, D => N27, Q => outPC(26))
                           ;
   outPC_reg_25_inst : DLH_X1 port map( G => n4_port, D => N26, Q => outPC(25))
                           ;
   outPC_reg_24_inst : DLH_X1 port map( G => n4_port, D => N25, Q => outPC(24))
                           ;
   outPC_reg_23_inst : DLH_X1 port map( G => n4_port, D => N24, Q => outPC(23))
                           ;
   outPC_reg_22_inst : DLH_X1 port map( G => n4_port, D => N23, Q => outPC(22))
                           ;
   outPC_reg_21_inst : DLH_X1 port map( G => n3_port, D => N22, Q => outPC(21))
                           ;
   outPC_reg_20_inst : DLH_X1 port map( G => n3_port, D => N21, Q => outPC(20))
                           ;
   outPC_reg_19_inst : DLH_X1 port map( G => n3_port, D => N20, Q => outPC(19))
                           ;
   outPC_reg_18_inst : DLH_X1 port map( G => n3_port, D => N19, Q => outPC(18))
                           ;
   outPC_reg_17_inst : DLH_X1 port map( G => n3_port, D => N18, Q => outPC(17))
                           ;
   outPC_reg_16_inst : DLH_X1 port map( G => n3_port, D => N17, Q => outPC(16))
                           ;
   outPC_reg_15_inst : DLH_X1 port map( G => n3_port, D => N16, Q => outPC(15))
                           ;
   outPC_reg_14_inst : DLH_X1 port map( G => n3_port, D => N15, Q => outPC(14))
                           ;
   outPC_reg_13_inst : DLH_X1 port map( G => n3_port, D => N14, Q => outPC(13))
                           ;
   outPC_reg_12_inst : DLH_X1 port map( G => n3_port, D => N13, Q => outPC(12))
                           ;
   outPC_reg_11_inst : DLH_X1 port map( G => n3_port, D => N12, Q => outPC(11))
                           ;
   outPC_reg_10_inst : DLH_X1 port map( G => n2_port, D => N11, Q => outPC(10))
                           ;
   outPC_reg_9_inst : DLH_X1 port map( G => n2_port, D => N10, Q => outPC(9));
   outPC_reg_8_inst : DLH_X1 port map( G => n2_port, D => N9, Q => outPC(8));
   outPC_reg_7_inst : DLH_X1 port map( G => n2_port, D => N8, Q => outPC(7));
   outPC_reg_6_inst : DLH_X1 port map( G => n2_port, D => N7, Q => outPC(6));
   outPC_reg_5_inst : DLH_X1 port map( G => n2_port, D => N6, Q => outPC(5));
   outPC_reg_4_inst : DLH_X1 port map( G => n2_port, D => N5, Q => outPC(4));
   outPC_reg_3_inst : DLH_X1 port map( G => n2_port, D => N4, Q => outPC(3));
   outPC_reg_2_inst : DLH_X1 port map( G => n2_port, D => N3, Q => outPC(2));
   outPC_reg_1_inst : DLH_X1 port map( G => n2_port, D => N2, Q => outPC(1));
   outPC_reg_0_inst : DLH_X1 port map( G => n2_port, D => N1, Q => outPC(0));
   n1_port <= '0';
   add_40 : NPC_adder_DW01_add_0 port map( A(31) => inPC(31), A(30) => inPC(30)
                           , A(29) => inPC(29), A(28) => inPC(28), A(27) => 
                           inPC(27), A(26) => inPC(26), A(25) => inPC(25), 
                           A(24) => inPC(24), A(23) => inPC(23), A(22) => 
                           inPC(22), A(21) => inPC(21), A(20) => inPC(20), 
                           A(19) => inPC(19), A(18) => inPC(18), A(17) => 
                           inPC(17), A(16) => inPC(16), A(15) => inPC(15), 
                           A(14) => inPC(14), A(13) => inPC(13), A(12) => 
                           inPC(12), A(11) => inPC(11), A(10) => inPC(10), A(9)
                           => inPC(9), A(8) => inPC(8), A(7) => inPC(7), A(6) 
                           => inPC(6), A(5) => inPC(5), A(4) => inPC(4), A(3) 
                           => inPC(3), A(2) => inPC(2), A(1) => inPC(1), A(0) 
                           => inPC(0), B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic1_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, CI => n1_port, SUM(31) => N32, 
                           SUM(30) => N31, SUM(29) => N30, SUM(28) => N29, 
                           SUM(27) => N28, SUM(26) => N27, SUM(25) => N26, 
                           SUM(24) => N25, SUM(23) => N24, SUM(22) => N23, 
                           SUM(21) => N22, SUM(20) => N21, SUM(19) => N20, 
                           SUM(18) => N19, SUM(17) => N18, SUM(16) => N17, 
                           SUM(15) => N16, SUM(14) => N15, SUM(13) => N14, 
                           SUM(12) => N13, SUM(11) => N12, SUM(10) => N11, 
                           SUM(9) => N10, SUM(8) => N9, SUM(7) => N8, SUM(6) =>
                           N7, SUM(5) => N6, SUM(4) => N5, SUM(3) => N4, SUM(2)
                           => N3, SUM(1) => N2, SUM(0) => N1, CO => n_1718);
   U4 : BUF_X1 port map( A => N0, Z => n2_port);
   U5 : BUF_X1 port map( A => N0, Z => n3_port);
   U6 : BUF_X1 port map( A => N0, Z => n4_port);
   U7 : INV_X1 port map( A => inPC(31), ZN => n17_port);
   U8 : NOR2_X1 port map( A1 => inPC(21), A2 => inPC(20), ZN => n8_port);
   U9 : NOR3_X1 port map( A1 => inPC(22), A2 => inPC(24), A3 => inPC(23), ZN =>
                           n7_port);
   U10 : NOR3_X1 port map( A1 => inPC(25), A2 => inPC(27), A3 => inPC(26), ZN 
                           => n6_port);
   U11 : NOR3_X1 port map( A1 => inPC(28), A2 => inPC(30), A3 => inPC(29), ZN 
                           => n5_port);
   U12 : NAND4_X1 port map( A1 => n8_port, A2 => n7_port, A3 => n6_port, A4 => 
                           n5_port, ZN => n16_port);
   U13 : AND4_X1 port map( A1 => inPC(9), A2 => inPC(8), A3 => inPC(7), A4 => 
                           inPC(6), ZN => n10_port);
   U14 : AND4_X1 port map( A1 => inPC(5), A2 => inPC(4), A3 => inPC(3), A4 => 
                           inPC(2), ZN => n9_port);
   U15 : AOI21_X1 port map( B1 => n10_port, B2 => n9_port, A => inPC(10), ZN =>
                           n14_port);
   U16 : NOR3_X1 port map( A1 => inPC(11), A2 => inPC(13), A3 => inPC(12), ZN 
                           => n13_port);
   U17 : NOR3_X1 port map( A1 => inPC(14), A2 => inPC(16), A3 => inPC(15), ZN 
                           => n12_port);
   U18 : NOR3_X1 port map( A1 => inPC(17), A2 => inPC(19), A3 => inPC(18), ZN 
                           => n11_port);
   U19 : NAND4_X1 port map( A1 => n14_port, A2 => n13_port, A3 => n12_port, A4 
                           => n11_port, ZN => n15_port);
   U20 : OAI21_X1 port map( B1 => n16_port, B2 => n15_port, A => n17_port, ZN 
                           => N0);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor is

   port( RST : in std_logic;  PC_IN, PC_FAIL, IR_IN : in std_logic_vector (31 
         downto 0);  IR_FAIL : in std_logic_vector (15 downto 0);  WRONG_PRE, 
         RIGHT_PRE : in std_logic;  NPC_OUT, LINK_ADD : out std_logic_vector 
         (31 downto 0);  SEL, TAKEN : out std_logic);

end branch_predictor;

architecture SYN_Behavioral of branch_predictor is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component branch_predictor_DW01_add_3
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component branch_predictor_DW01_add_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component branch_predictor_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component branch_predictor_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, CACHE_mem_0_1_port, CACHE_mem_0_0_port,
      CACHE_mem_1_1_port, CACHE_mem_1_0_port, CACHE_mem_2_1_port, 
      CACHE_mem_2_0_port, CACHE_mem_3_1_port, CACHE_mem_3_0_port, 
      CACHE_mem_4_1_port, CACHE_mem_4_0_port, CACHE_mem_5_1_port, 
      CACHE_mem_5_0_port, CACHE_mem_6_1_port, CACHE_mem_6_0_port, 
      CACHE_mem_7_1_port, CACHE_mem_7_0_port, CACHE_mem_8_1_port, 
      CACHE_mem_8_0_port, CACHE_mem_9_1_port, CACHE_mem_9_0_port, 
      CACHE_mem_10_1_port, CACHE_mem_10_0_port, CACHE_mem_11_1_port, 
      CACHE_mem_11_0_port, CACHE_mem_12_1_port, CACHE_mem_12_0_port, 
      CACHE_mem_13_1_port, CACHE_mem_13_0_port, CACHE_mem_14_1_port, 
      CACHE_mem_14_0_port, CACHE_mem_15_1_port, CACHE_mem_15_0_port, 
      CACHE_mem_16_1_port, CACHE_mem_16_0_port, CACHE_mem_17_1_port, 
      CACHE_mem_17_0_port, CACHE_mem_18_1_port, CACHE_mem_18_0_port, 
      CACHE_mem_19_1_port, CACHE_mem_19_0_port, CACHE_mem_20_1_port, 
      CACHE_mem_20_0_port, CACHE_mem_21_1_port, CACHE_mem_21_0_port, 
      CACHE_mem_22_1_port, CACHE_mem_22_0_port, CACHE_mem_23_1_port, 
      CACHE_mem_23_0_port, CACHE_mem_24_1_port, CACHE_mem_24_0_port, 
      CACHE_mem_25_1_port, CACHE_mem_25_0_port, CACHE_mem_26_1_port, 
      CACHE_mem_26_0_port, CACHE_mem_27_1_port, CACHE_mem_27_0_port, 
      CACHE_mem_28_1_port, CACHE_mem_28_0_port, CACHE_mem_29_1_port, 
      CACHE_mem_29_0_port, CACHE_mem_30_1_port, CACHE_mem_30_0_port, 
      CACHE_mem_31_1_port, CACHE_mem_31_0_port, N46, N47, N48, N49, N50, N51, 
      N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66
      , N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N81, N82, N83, 
      N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98
      , N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
      N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, 
      N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, 
      N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N216, N219, 
      N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, 
      N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, 
      N244, N245, N246, N247, N248, N249, N250, N323, N356, N357, N358, N359, 
      N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, 
      N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, 
      N384, N385, N386, N387, N388, N479, N480, N612, N613, N614, N615, N616, 
      N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, 
      N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, 
      N641, N642, N643, N644, N645, n1, n2, n3, n4, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, 
      n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, 
      n69_port, n70_port, n71_port, n72_port, n73_port, n74_port, n75_port, 
      n76_port, n77_port, n78, n79, n80, n81_port, n82_port, n83_port, n84_port
      , n85_port, n86_port, n87_port, n88_port, n89_port, n90_port, n91_port, 
      n92_port, n93_port, n94_port, n95_port, n96_port, n97_port, n98_port, 
      n99_port, n100_port, n101_port, n102_port, n103_port, n104_port, 
      n105_port, n106_port, n107_port, n108_port, n109_port, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46_port, n47_port, n48_port, 
      n49_port, n50_port, n51_port, n52_port, n110_port, n111_port, n112_port, 
      n113_port, n114_port, n115_port, n116_port, n117_port, n118_port, 
      n119_port, n120_port, n121_port, n122_port, n123_port, n124_port, 
      n125_port, n126_port, n127_port, n128_port, n129_port, n130_port, 
      n131_port, n132_port, n133_port, n134_port, n135_port, n136_port, 
      n137_port, n138_port, n139_port, n140_port, n141_port, n142_port, 
      n143_port, n144_port, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216_port, n217, n218, n219_port, n220_port, n221_port,
      n222_port, n223_port, n224_port, n225_port, n226_port, n227_port, 
      n228_port, n229_port, n230_port, n231_port, n232_port, n233_port, 
      n234_port, n235_port, n236_port, n237_port, n238_port, n239_port, n_1720,
      n_1721, n_1722, n_1723 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   NPC_OUT_reg_31_inst : DLH_X1 port map( G => n188, D => n199, Q => 
                           NPC_OUT(31));
   NPC_OUT_reg_30_inst : DLH_X1 port map( G => n188, D => n200, Q => 
                           NPC_OUT(30));
   NPC_OUT_reg_29_inst : DLH_X1 port map( G => n188, D => n201, Q => 
                           NPC_OUT(29));
   NPC_OUT_reg_28_inst : DLH_X1 port map( G => n188, D => n202, Q => 
                           NPC_OUT(28));
   NPC_OUT_reg_27_inst : DLH_X1 port map( G => n188, D => n203, Q => 
                           NPC_OUT(27));
   NPC_OUT_reg_26_inst : DLH_X1 port map( G => n188, D => n204, Q => 
                           NPC_OUT(26));
   NPC_OUT_reg_25_inst : DLH_X1 port map( G => n188, D => n205, Q => 
                           NPC_OUT(25));
   NPC_OUT_reg_24_inst : DLH_X1 port map( G => n188, D => n206, Q => 
                           NPC_OUT(24));
   NPC_OUT_reg_23_inst : DLH_X1 port map( G => n188, D => n207, Q => 
                           NPC_OUT(23));
   NPC_OUT_reg_22_inst : DLH_X1 port map( G => n188, D => n208, Q => 
                           NPC_OUT(22));
   NPC_OUT_reg_21_inst : DLH_X1 port map( G => n188, D => n209, Q => 
                           NPC_OUT(21));
   NPC_OUT_reg_20_inst : DLH_X1 port map( G => n189, D => n210, Q => 
                           NPC_OUT(20));
   NPC_OUT_reg_19_inst : DLH_X1 port map( G => n189, D => n211, Q => 
                           NPC_OUT(19));
   NPC_OUT_reg_18_inst : DLH_X1 port map( G => n189, D => n212, Q => 
                           NPC_OUT(18));
   NPC_OUT_reg_17_inst : DLH_X1 port map( G => n189, D => n213, Q => 
                           NPC_OUT(17));
   NPC_OUT_reg_16_inst : DLH_X1 port map( G => n189, D => n214, Q => 
                           NPC_OUT(16));
   NPC_OUT_reg_15_inst : DLH_X1 port map( G => n189, D => n215, Q => 
                           NPC_OUT(15));
   NPC_OUT_reg_14_inst : DLH_X1 port map( G => n189, D => n216_port, Q => 
                           NPC_OUT(14));
   NPC_OUT_reg_13_inst : DLH_X1 port map( G => n189, D => n217, Q => 
                           NPC_OUT(13));
   NPC_OUT_reg_12_inst : DLH_X1 port map( G => n189, D => n218, Q => 
                           NPC_OUT(12));
   NPC_OUT_reg_11_inst : DLH_X1 port map( G => n189, D => n219_port, Q => 
                           NPC_OUT(11));
   NPC_OUT_reg_10_inst : DLH_X1 port map( G => n189, D => n220_port, Q => 
                           NPC_OUT(10));
   NPC_OUT_reg_9_inst : DLH_X1 port map( G => n190, D => n221_port, Q => 
                           NPC_OUT(9));
   NPC_OUT_reg_8_inst : DLH_X1 port map( G => n190, D => n222_port, Q => 
                           NPC_OUT(8));
   NPC_OUT_reg_7_inst : DLH_X1 port map( G => n190, D => n223_port, Q => 
                           NPC_OUT(7));
   NPC_OUT_reg_6_inst : DLH_X1 port map( G => n190, D => n224_port, Q => 
                           NPC_OUT(6));
   NPC_OUT_reg_5_inst : DLH_X1 port map( G => n190, D => n225_port, Q => 
                           NPC_OUT(5));
   NPC_OUT_reg_4_inst : DLH_X1 port map( G => n190, D => n226_port, Q => 
                           NPC_OUT(4));
   NPC_OUT_reg_3_inst : DLH_X1 port map( G => n190, D => n227_port, Q => 
                           NPC_OUT(3));
   NPC_OUT_reg_2_inst : DLH_X1 port map( G => n190, D => n228_port, Q => 
                           NPC_OUT(2));
   NPC_OUT_reg_1_inst : DLH_X1 port map( G => n190, D => n229_port, Q => 
                           NPC_OUT(1));
   NPC_OUT_reg_0_inst : DLH_X1 port map( G => n190, D => n230_port, Q => 
                           NPC_OUT(0));
   LINK_ADD_reg_31_inst : DLH_X1 port map( G => n186, D => N388, Q => 
                           LINK_ADD(31));
   LINK_ADD_reg_30_inst : DLH_X1 port map( G => n186, D => N387, Q => 
                           LINK_ADD(30));
   LINK_ADD_reg_29_inst : DLH_X1 port map( G => n186, D => N386, Q => 
                           LINK_ADD(29));
   LINK_ADD_reg_28_inst : DLH_X1 port map( G => n186, D => N385, Q => 
                           LINK_ADD(28));
   LINK_ADD_reg_27_inst : DLH_X1 port map( G => n186, D => N384, Q => 
                           LINK_ADD(27));
   LINK_ADD_reg_26_inst : DLH_X1 port map( G => n186, D => N383, Q => 
                           LINK_ADD(26));
   LINK_ADD_reg_25_inst : DLH_X1 port map( G => n186, D => N382, Q => 
                           LINK_ADD(25));
   LINK_ADD_reg_24_inst : DLH_X1 port map( G => n186, D => N381, Q => 
                           LINK_ADD(24));
   LINK_ADD_reg_23_inst : DLH_X1 port map( G => n186, D => N380, Q => 
                           LINK_ADD(23));
   LINK_ADD_reg_22_inst : DLH_X1 port map( G => n186, D => N379, Q => 
                           LINK_ADD(22));
   LINK_ADD_reg_21_inst : DLH_X1 port map( G => n186, D => N378, Q => 
                           LINK_ADD(21));
   LINK_ADD_reg_20_inst : DLH_X1 port map( G => n186, D => N377, Q => 
                           LINK_ADD(20));
   LINK_ADD_reg_19_inst : DLH_X1 port map( G => n186, D => N376, Q => 
                           LINK_ADD(19));
   LINK_ADD_reg_18_inst : DLH_X1 port map( G => n186, D => N375, Q => 
                           LINK_ADD(18));
   LINK_ADD_reg_17_inst : DLH_X1 port map( G => n186, D => N374, Q => 
                           LINK_ADD(17));
   LINK_ADD_reg_16_inst : DLH_X1 port map( G => n186, D => N373, Q => 
                           LINK_ADD(16));
   LINK_ADD_reg_15_inst : DLH_X1 port map( G => n186, D => N372, Q => 
                           LINK_ADD(15));
   LINK_ADD_reg_14_inst : DLH_X1 port map( G => n186, D => N371, Q => 
                           LINK_ADD(14));
   LINK_ADD_reg_13_inst : DLH_X1 port map( G => n186, D => N370, Q => 
                           LINK_ADD(13));
   LINK_ADD_reg_12_inst : DLH_X1 port map( G => n186, D => N369, Q => 
                           LINK_ADD(12));
   LINK_ADD_reg_11_inst : DLH_X1 port map( G => n186, D => N368, Q => 
                           LINK_ADD(11));
   LINK_ADD_reg_10_inst : DLH_X1 port map( G => n186, D => N367, Q => 
                           LINK_ADD(10));
   LINK_ADD_reg_9_inst : DLH_X1 port map( G => n186, D => N366, Q => 
                           LINK_ADD(9));
   LINK_ADD_reg_8_inst : DLH_X1 port map( G => n186, D => N365, Q => 
                           LINK_ADD(8));
   LINK_ADD_reg_7_inst : DLH_X1 port map( G => n187, D => N364, Q => 
                           LINK_ADD(7));
   LINK_ADD_reg_6_inst : DLH_X1 port map( G => n187, D => N363, Q => 
                           LINK_ADD(6));
   LINK_ADD_reg_5_inst : DLH_X1 port map( G => n187, D => N362, Q => 
                           LINK_ADD(5));
   LINK_ADD_reg_4_inst : DLH_X1 port map( G => n187, D => N361, Q => 
                           LINK_ADD(4));
   LINK_ADD_reg_3_inst : DLH_X1 port map( G => n187, D => N360, Q => 
                           LINK_ADD(3));
   LINK_ADD_reg_2_inst : DLH_X1 port map( G => n187, D => N359, Q => 
                           LINK_ADD(2));
   LINK_ADD_reg_1_inst : DLH_X1 port map( G => n187, D => N358, Q => 
                           LINK_ADD(1));
   LINK_ADD_reg_0_inst : DLH_X1 port map( G => n187, D => N357, Q => 
                           LINK_ADD(0));
   CACHE_mem_reg_0_1_inst : DLH_X1 port map( G => N643, D => n180, Q => 
                           CACHE_mem_0_1_port);
   CACHE_mem_reg_0_0_inst : DLH_X1 port map( G => N643, D => n183, Q => 
                           CACHE_mem_0_0_port);
   CACHE_mem_reg_1_1_inst : DLH_X1 port map( G => N642, D => n180, Q => 
                           CACHE_mem_1_1_port);
   CACHE_mem_reg_1_0_inst : DLH_X1 port map( G => N642, D => n183, Q => 
                           CACHE_mem_1_0_port);
   CACHE_mem_reg_2_1_inst : DLH_X1 port map( G => N641, D => n180, Q => 
                           CACHE_mem_2_1_port);
   CACHE_mem_reg_2_0_inst : DLH_X1 port map( G => N641, D => n183, Q => 
                           CACHE_mem_2_0_port);
   CACHE_mem_reg_3_1_inst : DLH_X1 port map( G => N640, D => n180, Q => 
                           CACHE_mem_3_1_port);
   CACHE_mem_reg_3_0_inst : DLH_X1 port map( G => N640, D => n183, Q => 
                           CACHE_mem_3_0_port);
   CACHE_mem_reg_4_1_inst : DLH_X1 port map( G => N639, D => n180, Q => 
                           CACHE_mem_4_1_port);
   CACHE_mem_reg_4_0_inst : DLH_X1 port map( G => N639, D => n183, Q => 
                           CACHE_mem_4_0_port);
   CACHE_mem_reg_5_1_inst : DLH_X1 port map( G => N638, D => n180, Q => 
                           CACHE_mem_5_1_port);
   CACHE_mem_reg_5_0_inst : DLH_X1 port map( G => N638, D => n183, Q => 
                           CACHE_mem_5_0_port);
   CACHE_mem_reg_6_1_inst : DLH_X1 port map( G => N637, D => n180, Q => 
                           CACHE_mem_6_1_port);
   CACHE_mem_reg_6_0_inst : DLH_X1 port map( G => N637, D => n183, Q => 
                           CACHE_mem_6_0_port);
   CACHE_mem_reg_7_1_inst : DLH_X1 port map( G => N636, D => n180, Q => 
                           CACHE_mem_7_1_port);
   CACHE_mem_reg_7_0_inst : DLH_X1 port map( G => N636, D => n183, Q => 
                           CACHE_mem_7_0_port);
   CACHE_mem_reg_8_1_inst : DLH_X1 port map( G => N635, D => n180, Q => 
                           CACHE_mem_8_1_port);
   CACHE_mem_reg_8_0_inst : DLH_X1 port map( G => N635, D => n183, Q => 
                           CACHE_mem_8_0_port);
   CACHE_mem_reg_9_1_inst : DLH_X1 port map( G => N634, D => n180, Q => 
                           CACHE_mem_9_1_port);
   CACHE_mem_reg_9_0_inst : DLH_X1 port map( G => N634, D => n183, Q => 
                           CACHE_mem_9_0_port);
   CACHE_mem_reg_10_1_inst : DLH_X1 port map( G => N633, D => n180, Q => 
                           CACHE_mem_10_1_port);
   CACHE_mem_reg_10_0_inst : DLH_X1 port map( G => N633, D => n183, Q => 
                           CACHE_mem_10_0_port);
   CACHE_mem_reg_11_1_inst : DLH_X1 port map( G => N632, D => n181, Q => 
                           CACHE_mem_11_1_port);
   CACHE_mem_reg_11_0_inst : DLH_X1 port map( G => N632, D => n184, Q => 
                           CACHE_mem_11_0_port);
   CACHE_mem_reg_12_1_inst : DLH_X1 port map( G => N631, D => n181, Q => 
                           CACHE_mem_12_1_port);
   CACHE_mem_reg_12_0_inst : DLH_X1 port map( G => N631, D => n184, Q => 
                           CACHE_mem_12_0_port);
   CACHE_mem_reg_13_1_inst : DLH_X1 port map( G => N630, D => n181, Q => 
                           CACHE_mem_13_1_port);
   CACHE_mem_reg_13_0_inst : DLH_X1 port map( G => N630, D => n184, Q => 
                           CACHE_mem_13_0_port);
   CACHE_mem_reg_14_1_inst : DLH_X1 port map( G => N629, D => n181, Q => 
                           CACHE_mem_14_1_port);
   CACHE_mem_reg_14_0_inst : DLH_X1 port map( G => N629, D => n184, Q => 
                           CACHE_mem_14_0_port);
   CACHE_mem_reg_15_1_inst : DLH_X1 port map( G => N628, D => n181, Q => 
                           CACHE_mem_15_1_port);
   CACHE_mem_reg_15_0_inst : DLH_X1 port map( G => N628, D => n184, Q => 
                           CACHE_mem_15_0_port);
   CACHE_mem_reg_16_1_inst : DLH_X1 port map( G => N627, D => n181, Q => 
                           CACHE_mem_16_1_port);
   CACHE_mem_reg_16_0_inst : DLH_X1 port map( G => N627, D => n184, Q => 
                           CACHE_mem_16_0_port);
   CACHE_mem_reg_17_1_inst : DLH_X1 port map( G => N626, D => n181, Q => 
                           CACHE_mem_17_1_port);
   CACHE_mem_reg_17_0_inst : DLH_X1 port map( G => N626, D => n184, Q => 
                           CACHE_mem_17_0_port);
   CACHE_mem_reg_18_1_inst : DLH_X1 port map( G => N625, D => n181, Q => 
                           CACHE_mem_18_1_port);
   CACHE_mem_reg_18_0_inst : DLH_X1 port map( G => N625, D => n184, Q => 
                           CACHE_mem_18_0_port);
   CACHE_mem_reg_19_1_inst : DLH_X1 port map( G => N624, D => n181, Q => 
                           CACHE_mem_19_1_port);
   CACHE_mem_reg_19_0_inst : DLH_X1 port map( G => N624, D => n184, Q => 
                           CACHE_mem_19_0_port);
   CACHE_mem_reg_20_1_inst : DLH_X1 port map( G => N623, D => n181, Q => 
                           CACHE_mem_20_1_port);
   CACHE_mem_reg_20_0_inst : DLH_X1 port map( G => N623, D => n184, Q => 
                           CACHE_mem_20_0_port);
   CACHE_mem_reg_21_1_inst : DLH_X1 port map( G => N622, D => n181, Q => 
                           CACHE_mem_21_1_port);
   CACHE_mem_reg_21_0_inst : DLH_X1 port map( G => N622, D => n184, Q => 
                           CACHE_mem_21_0_port);
   CACHE_mem_reg_22_1_inst : DLH_X1 port map( G => N621, D => n182, Q => 
                           CACHE_mem_22_1_port);
   CACHE_mem_reg_22_0_inst : DLH_X1 port map( G => N621, D => n185, Q => 
                           CACHE_mem_22_0_port);
   CACHE_mem_reg_23_1_inst : DLH_X1 port map( G => N620, D => n182, Q => 
                           CACHE_mem_23_1_port);
   CACHE_mem_reg_23_0_inst : DLH_X1 port map( G => N620, D => n185, Q => 
                           CACHE_mem_23_0_port);
   CACHE_mem_reg_24_1_inst : DLH_X1 port map( G => N619, D => n182, Q => 
                           CACHE_mem_24_1_port);
   CACHE_mem_reg_24_0_inst : DLH_X1 port map( G => N619, D => n185, Q => 
                           CACHE_mem_24_0_port);
   CACHE_mem_reg_25_1_inst : DLH_X1 port map( G => N618, D => n182, Q => 
                           CACHE_mem_25_1_port);
   CACHE_mem_reg_25_0_inst : DLH_X1 port map( G => N618, D => n185, Q => 
                           CACHE_mem_25_0_port);
   CACHE_mem_reg_26_1_inst : DLH_X1 port map( G => N617, D => n182, Q => 
                           CACHE_mem_26_1_port);
   CACHE_mem_reg_26_0_inst : DLH_X1 port map( G => N617, D => n185, Q => 
                           CACHE_mem_26_0_port);
   CACHE_mem_reg_27_1_inst : DLH_X1 port map( G => N616, D => n182, Q => 
                           CACHE_mem_27_1_port);
   CACHE_mem_reg_27_0_inst : DLH_X1 port map( G => N616, D => n185, Q => 
                           CACHE_mem_27_0_port);
   CACHE_mem_reg_28_1_inst : DLH_X1 port map( G => N615, D => n182, Q => 
                           CACHE_mem_28_1_port);
   CACHE_mem_reg_28_0_inst : DLH_X1 port map( G => N615, D => n185, Q => 
                           CACHE_mem_28_0_port);
   CACHE_mem_reg_29_1_inst : DLH_X1 port map( G => N614, D => n182, Q => 
                           CACHE_mem_29_1_port);
   CACHE_mem_reg_29_0_inst : DLH_X1 port map( G => N614, D => n185, Q => 
                           CACHE_mem_29_0_port);
   CACHE_mem_reg_30_1_inst : DLH_X1 port map( G => N613, D => n182, Q => 
                           CACHE_mem_30_1_port);
   CACHE_mem_reg_30_0_inst : DLH_X1 port map( G => N613, D => n185, Q => 
                           CACHE_mem_30_0_port);
   CACHE_mem_reg_31_1_inst : DLH_X1 port map( G => N612, D => n182, Q => 
                           CACHE_mem_31_1_port);
   CACHE_mem_reg_31_0_inst : DLH_X1 port map( G => N612, D => n185, Q => 
                           CACHE_mem_31_0_port);
   U166 : NAND3_X1 port map( A1 => n233_port, A2 => n191, A3 => n69_port, ZN =>
                           n60_port);
   U167 : NAND3_X1 port map( A1 => n69_port, A2 => n191, A3 => PC_FAIL(5), ZN 
                           => n70_port);
   U168 : NAND3_X1 port map( A1 => n69_port, A2 => n233_port, A3 => PC_FAIL(6),
                           ZN => n71_port);
   U169 : NAND3_X1 port map( A1 => n235_port, A2 => n234_port, A3 => n236_port,
                           ZN => n61_port);
   U170 : NAND3_X1 port map( A1 => n235_port, A2 => n234_port, A3 => PC_FAIL(2)
                           , ZN => n62_port);
   U171 : NAND3_X1 port map( A1 => n236_port, A2 => n234_port, A3 => PC_FAIL(3)
                           , ZN => n63_port);
   U172 : NAND3_X1 port map( A1 => PC_FAIL(2), A2 => n234_port, A3 => 
                           PC_FAIL(3), ZN => n64_port);
   U173 : NAND3_X1 port map( A1 => n236_port, A2 => n235_port, A3 => PC_FAIL(4)
                           , ZN => n65_port);
   U174 : NAND3_X1 port map( A1 => PC_FAIL(2), A2 => n235_port, A3 => 
                           PC_FAIL(4), ZN => n66_port);
   U175 : NAND3_X1 port map( A1 => PC_FAIL(3), A2 => n236_port, A3 => 
                           PC_FAIL(4), ZN => n67_port);
   U176 : NAND3_X1 port map( A1 => PC_FAIL(5), A2 => n69_port, A3 => PC_FAIL(6)
                           , ZN => n72_port);
   U177 : NAND3_X1 port map( A1 => PC_FAIL(3), A2 => PC_FAIL(2), A3 => 
                           PC_FAIL(4), ZN => n68_port);
   U178 : NAND3_X1 port map( A1 => n109_port, A2 => n239_port, A3 => IR_IN(27),
                           ZN => n108_port);
   add_65 : branch_predictor_DW01_add_0 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => 
                           IR_IN(15), B(30) => IR_IN(15), B(29) => IR_IN(15), 
                           B(28) => IR_IN(15), B(27) => IR_IN(15), B(26) => 
                           IR_IN(15), B(25) => IR_IN(15), B(24) => IR_IN(15), 
                           B(23) => IR_IN(15), B(22) => IR_IN(15), B(21) => 
                           IR_IN(15), B(20) => IR_IN(15), B(19) => IR_IN(15), 
                           B(18) => IR_IN(15), B(17) => IR_IN(15), B(16) => 
                           IR_IN(15), B(15) => IR_IN(15), B(14) => IR_IN(14), 
                           B(13) => IR_IN(13), B(12) => IR_IN(12), B(11) => 
                           IR_IN(11), B(10) => IR_IN(10), B(9) => IR_IN(9), 
                           B(8) => IR_IN(8), B(7) => IR_IN(7), B(6) => IR_IN(6)
                           , B(5) => IR_IN(5), B(4) => IR_IN(4), B(3) => 
                           IR_IN(3), B(2) => IR_IN(2), B(1) => IR_IN(1), B(0) 
                           => IR_IN(0), CI => n1, SUM(31) => N250, SUM(30) => 
                           N249, SUM(29) => N248, SUM(28) => N247, SUM(27) => 
                           N246, SUM(26) => N245, SUM(25) => N244, SUM(24) => 
                           N243, SUM(23) => N242, SUM(22) => N241, SUM(21) => 
                           N240, SUM(20) => N239, SUM(19) => N238, SUM(18) => 
                           N237, SUM(17) => N236, SUM(16) => N235, SUM(15) => 
                           N234, SUM(14) => N233, SUM(13) => N232, SUM(12) => 
                           N231, SUM(11) => N230, SUM(10) => N229, SUM(9) => 
                           N228, SUM(8) => N227, SUM(7) => N226, SUM(6) => N225
                           , SUM(5) => N224, SUM(4) => N223, SUM(3) => N222, 
                           SUM(2) => N221, SUM(1) => N220, SUM(0) => N219, CO 
                           => n_1720);
   add_60 : branch_predictor_DW01_add_1 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => 
                           X_Logic0_port, B(30) => X_Logic0_port, B(29) => 
                           X_Logic0_port, B(28) => X_Logic0_port, B(27) => 
                           X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic1_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, CI => n2, 
                           SUM(31) => N144, SUM(30) => N143, SUM(29) => N142, 
                           SUM(28) => N141, SUM(27) => N140, SUM(26) => N139, 
                           SUM(25) => N138, SUM(24) => N137, SUM(23) => N136, 
                           SUM(22) => N135, SUM(21) => N134, SUM(20) => N133, 
                           SUM(19) => N132, SUM(18) => N131, SUM(17) => N130, 
                           SUM(16) => N129, SUM(15) => N128, SUM(14) => N127, 
                           SUM(13) => N126, SUM(12) => N125, SUM(11) => N124, 
                           SUM(10) => N123, SUM(9) => N122, SUM(8) => N121, 
                           SUM(7) => N120, SUM(6) => N119, SUM(5) => N118, 
                           SUM(4) => N117, SUM(3) => N116, SUM(2) => N115, 
                           SUM(1) => N114, SUM(0) => N113, CO => n_1721);
   add_59 : branch_predictor_DW01_add_2 port map( A(31) => PC_IN(31), A(30) => 
                           PC_IN(30), A(29) => PC_IN(29), A(28) => PC_IN(28), 
                           A(27) => PC_IN(27), A(26) => PC_IN(26), A(25) => 
                           PC_IN(25), A(24) => PC_IN(24), A(23) => PC_IN(23), 
                           A(22) => PC_IN(22), A(21) => PC_IN(21), A(20) => 
                           PC_IN(20), A(19) => PC_IN(19), A(18) => PC_IN(18), 
                           A(17) => PC_IN(17), A(16) => PC_IN(16), A(15) => 
                           PC_IN(15), A(14) => PC_IN(14), A(13) => PC_IN(13), 
                           A(12) => PC_IN(12), A(11) => PC_IN(11), A(10) => 
                           PC_IN(10), A(9) => PC_IN(9), A(8) => PC_IN(8), A(7) 
                           => PC_IN(7), A(6) => PC_IN(6), A(5) => PC_IN(5), 
                           A(4) => PC_IN(4), A(3) => PC_IN(3), A(2) => PC_IN(2)
                           , A(1) => PC_IN(1), A(0) => PC_IN(0), B(31) => 
                           IR_IN(25), B(30) => IR_IN(25), B(29) => IR_IN(25), 
                           B(28) => IR_IN(25), B(27) => IR_IN(25), B(26) => 
                           IR_IN(25), B(25) => IR_IN(25), B(24) => IR_IN(24), 
                           B(23) => IR_IN(23), B(22) => IR_IN(22), B(21) => 
                           IR_IN(21), B(20) => IR_IN(20), B(19) => IR_IN(19), 
                           B(18) => IR_IN(18), B(17) => IR_IN(17), B(16) => 
                           IR_IN(16), B(15) => IR_IN(15), B(14) => IR_IN(14), 
                           B(13) => IR_IN(13), B(12) => IR_IN(12), B(11) => 
                           IR_IN(11), B(10) => IR_IN(10), B(9) => IR_IN(9), 
                           B(8) => IR_IN(8), B(7) => IR_IN(7), B(6) => IR_IN(6)
                           , B(5) => IR_IN(5), B(4) => IR_IN(4), B(3) => 
                           IR_IN(3), B(2) => IR_IN(2), B(1) => IR_IN(1), B(0) 
                           => IR_IN(0), CI => n3, SUM(31) => N112, SUM(30) => 
                           N111, SUM(29) => N110, SUM(28) => N109, SUM(27) => 
                           N108, SUM(26) => N107, SUM(25) => N106, SUM(24) => 
                           N105, SUM(23) => N104, SUM(22) => N103, SUM(21) => 
                           N102, SUM(20) => N101, SUM(19) => N100, SUM(18) => 
                           N99, SUM(17) => N98, SUM(16) => N97, SUM(15) => N96,
                           SUM(14) => N95, SUM(13) => N94, SUM(12) => N93, 
                           SUM(11) => N92, SUM(10) => N91, SUM(9) => N90, 
                           SUM(8) => N89, SUM(7) => N88, SUM(6) => N87, SUM(5) 
                           => N86, SUM(4) => N85, SUM(3) => N84, SUM(2) => N83,
                           SUM(1) => N82, SUM(0) => N81, CO => n_1722);
   add_53_aco : branch_predictor_DW01_add_3 port map( A(31) => PC_FAIL(31), 
                           A(30) => PC_FAIL(30), A(29) => PC_FAIL(29), A(28) =>
                           PC_FAIL(28), A(27) => PC_FAIL(27), A(26) => 
                           PC_FAIL(26), A(25) => PC_FAIL(25), A(24) => 
                           PC_FAIL(24), A(23) => PC_FAIL(23), A(22) => 
                           PC_FAIL(22), A(21) => PC_FAIL(21), A(20) => 
                           PC_FAIL(20), A(19) => PC_FAIL(19), A(18) => 
                           PC_FAIL(18), A(17) => PC_FAIL(17), A(16) => 
                           PC_FAIL(16), A(15) => PC_FAIL(15), A(14) => 
                           PC_FAIL(14), A(13) => PC_FAIL(13), A(12) => 
                           PC_FAIL(12), A(11) => PC_FAIL(11), A(10) => 
                           PC_FAIL(10), A(9) => PC_FAIL(9), A(8) => PC_FAIL(8),
                           A(7) => PC_FAIL(7), A(6) => PC_FAIL(6), A(5) => 
                           PC_FAIL(5), A(4) => PC_FAIL(4), A(3) => PC_FAIL(3), 
                           A(2) => PC_FAIL(2), A(1) => PC_FAIL(1), A(0) => 
                           PC_FAIL(0), B(31) => n5, B(30) => n5, B(29) => n5, 
                           B(28) => n5, B(27) => n5, B(26) => n5, B(25) => n5, 
                           B(24) => n5, B(23) => n5, B(22) => n5, B(21) => n5, 
                           B(20) => n5, B(19) => n5, B(18) => n5, B(17) => n5, 
                           B(16) => n5, B(15) => n5, B(14) => n19, B(13) => n18
                           , B(12) => n17, B(11) => n16, B(10) => n15, B(9) => 
                           n14, B(8) => n13, B(7) => n12, B(6) => n11, B(5) => 
                           n7, B(4) => n10, B(3) => n9, B(2) => n8, B(1) => n6,
                           B(0) => n20, CI => n4, SUM(31) => N77, SUM(30) => 
                           N76, SUM(29) => N75, SUM(28) => N74, SUM(27) => N73,
                           SUM(26) => N72, SUM(25) => N71, SUM(24) => N70, 
                           SUM(23) => N69, SUM(22) => N68, SUM(21) => N67, 
                           SUM(20) => N66, SUM(19) => N65, SUM(18) => N64, 
                           SUM(17) => N63, SUM(16) => N62, SUM(15) => N61, 
                           SUM(14) => N60, SUM(13) => N59, SUM(12) => N58, 
                           SUM(11) => N57, SUM(10) => N56, SUM(9) => N55, 
                           SUM(8) => N54, SUM(7) => N53, SUM(6) => N52, SUM(5) 
                           => N51, SUM(4) => N50, SUM(3) => N49, SUM(2) => N48,
                           SUM(1) => N47, SUM(0) => N46, CO => n_1723);
   U3 : AND2_X1 port map( A1 => N116, A2 => n192, ZN => N360);
   U4 : AND2_X1 port map( A1 => N117, A2 => n193, ZN => N361);
   U5 : AND2_X1 port map( A1 => N118, A2 => n192, ZN => N362);
   U6 : AND2_X1 port map( A1 => N119, A2 => n195, ZN => N363);
   U7 : AND2_X1 port map( A1 => N120, A2 => n195, ZN => N364);
   U8 : AND2_X1 port map( A1 => N121, A2 => n195, ZN => N365);
   U9 : AND2_X1 port map( A1 => N122, A2 => n195, ZN => N366);
   U14 : AND2_X1 port map( A1 => N123, A2 => n195, ZN => N367);
   U15 : AND2_X1 port map( A1 => N124, A2 => n195, ZN => N368);
   U16 : AND2_X1 port map( A1 => N125, A2 => n195, ZN => N369);
   U17 : AND2_X1 port map( A1 => N126, A2 => n195, ZN => N370);
   U18 : AND2_X1 port map( A1 => N127, A2 => n194, ZN => N371);
   U19 : AND2_X1 port map( A1 => N128, A2 => n195, ZN => N372);
   U20 : AND2_X1 port map( A1 => N129, A2 => n195, ZN => N373);
   U21 : AND2_X1 port map( A1 => N130, A2 => n195, ZN => N374);
   U22 : AND2_X1 port map( A1 => N131, A2 => n195, ZN => N375);
   U23 : AND2_X1 port map( A1 => N132, A2 => n195, ZN => N376);
   U24 : AND2_X1 port map( A1 => N133, A2 => n195, ZN => N377);
   U25 : AND2_X1 port map( A1 => N134, A2 => n195, ZN => N378);
   U26 : AND2_X1 port map( A1 => N135, A2 => n195, ZN => N379);
   U27 : AND2_X1 port map( A1 => N136, A2 => n195, ZN => N380);
   U28 : AND2_X1 port map( A1 => N137, A2 => n195, ZN => N381);
   U29 : AND2_X1 port map( A1 => N138, A2 => n195, ZN => N382);
   U30 : AND2_X1 port map( A1 => N139, A2 => n195, ZN => N383);
   U31 : AND2_X1 port map( A1 => N140, A2 => n194, ZN => N384);
   U32 : AND2_X1 port map( A1 => N141, A2 => n194, ZN => N385);
   U33 : AND2_X1 port map( A1 => N142, A2 => n194, ZN => N386);
   U34 : AND2_X1 port map( A1 => N143, A2 => n194, ZN => N387);
   U35 : AND2_X1 port map( A1 => N144, A2 => n194, ZN => N388);
   U36 : AND2_X2 port map( A1 => IR_FAIL(15), A2 => N479, ZN => n5);
   U37 : AND2_X1 port map( A1 => IR_FAIL(1), A2 => N479, ZN => n6);
   U38 : BUF_X1 port map( A => n231_port, Z => n173);
   U39 : BUF_X1 port map( A => n231_port, Z => n171);
   U40 : BUF_X1 port map( A => n231_port, Z => n172);
   U41 : BUF_X1 port map( A => n75_port, Z => n174);
   U42 : BUF_X1 port map( A => n75_port, Z => n175);
   U43 : BUF_X1 port map( A => n75_port, Z => n176);
   U44 : INV_X1 port map( A => n56_port, ZN => n231_port);
   U45 : BUF_X1 port map( A => n53_port, Z => n179);
   U46 : NOR2_X1 port map( A1 => n197, A2 => WRONG_PRE, ZN => n107_port);
   U47 : INV_X1 port map( A => n198, ZN => n192);
   U48 : INV_X1 port map( A => n198, ZN => n193);
   U49 : INV_X1 port map( A => n197, ZN => n195);
   U50 : INV_X1 port map( A => n198, ZN => n194);
   U51 : BUF_X1 port map( A => n53_port, Z => n177);
   U52 : BUF_X1 port map( A => n53_port, Z => n178);
   U53 : OAI21_X1 port map( B1 => n60_port, B2 => n61_port, A => n193, ZN => 
                           N643);
   U54 : BUF_X1 port map( A => N356, Z => n186);
   U55 : NAND2_X1 port map( A1 => WRONG_PRE, A2 => n192, ZN => n56_port);
   U56 : BUF_X1 port map( A => PC_FAIL(6), Z => n140_port);
   U57 : BUF_X1 port map( A => PC_FAIL(6), Z => n139_port);
   U58 : OAI21_X1 port map( B1 => n61_port, B2 => n71_port, A => n193, ZN => 
                           N627);
   U59 : BUF_X1 port map( A => PC_FAIL(6), Z => n138_port);
   U60 : BUF_X1 port map( A => N323, Z => n189);
   U61 : BUF_X1 port map( A => N323, Z => n188);
   U62 : BUF_X1 port map( A => N644, Z => n184);
   U63 : BUF_X1 port map( A => N644, Z => n183);
   U64 : BUF_X1 port map( A => N645, Z => n181);
   U65 : BUF_X1 port map( A => N645, Z => n180);
   U66 : BUF_X1 port map( A => N323, Z => n190);
   U67 : AND2_X1 port map( A1 => n238_port, A2 => n107_port, ZN => n75_port);
   U68 : BUF_X1 port map( A => N644, Z => n185);
   U69 : BUF_X1 port map( A => N645, Z => n182);
   U70 : BUF_X1 port map( A => N356, Z => n187);
   U71 : AND2_X1 port map( A1 => n107_port, A2 => n108_port, ZN => n53_port);
   U72 : AND2_X1 port map( A1 => n179, A2 => n54_port, ZN => TAKEN);
   U73 : OAI21_X1 port map( B1 => n60_port, B2 => n68_port, A => n192, ZN => 
                           N636);
   U74 : OAI21_X1 port map( B1 => n60_port, B2 => n67_port, A => n192, ZN => 
                           N637);
   U75 : OAI21_X1 port map( B1 => n60_port, B2 => n66_port, A => n192, ZN => 
                           N638);
   U76 : OAI21_X1 port map( B1 => n60_port, B2 => n65_port, A => n192, ZN => 
                           N639);
   U77 : OAI21_X1 port map( B1 => n60_port, B2 => n64_port, A => n192, ZN => 
                           N640);
   U78 : OAI21_X1 port map( B1 => n60_port, B2 => n63_port, A => n192, ZN => 
                           N641);
   U79 : OAI21_X1 port map( B1 => n60_port, B2 => n62_port, A => n192, ZN => 
                           N642);
   U80 : OAI21_X1 port map( B1 => n68_port, B2 => n72_port, A => n194, ZN => 
                           N612);
   U81 : OAI21_X1 port map( B1 => n67_port, B2 => n72_port, A => n194, ZN => 
                           N613);
   U82 : OAI21_X1 port map( B1 => n66_port, B2 => n72_port, A => n194, ZN => 
                           N614);
   U83 : OAI21_X1 port map( B1 => n65_port, B2 => n72_port, A => n194, ZN => 
                           N615);
   U84 : OAI21_X1 port map( B1 => n64_port, B2 => n72_port, A => n194, ZN => 
                           N616);
   U85 : OAI21_X1 port map( B1 => n63_port, B2 => n72_port, A => n194, ZN => 
                           N617);
   U86 : OAI21_X1 port map( B1 => n62_port, B2 => n72_port, A => n194, ZN => 
                           N618);
   U87 : OAI21_X1 port map( B1 => n61_port, B2 => n72_port, A => n194, ZN => 
                           N619);
   U88 : OAI21_X1 port map( B1 => n68_port, B2 => n70_port, A => n193, ZN => 
                           N628);
   U89 : OAI21_X1 port map( B1 => n67_port, B2 => n70_port, A => n193, ZN => 
                           N629);
   U90 : OAI21_X1 port map( B1 => n66_port, B2 => n70_port, A => n193, ZN => 
                           N630);
   U91 : OAI21_X1 port map( B1 => n65_port, B2 => n70_port, A => n192, ZN => 
                           N631);
   U92 : OAI21_X1 port map( B1 => n64_port, B2 => n70_port, A => n193, ZN => 
                           N632);
   U93 : OAI21_X1 port map( B1 => n63_port, B2 => n70_port, A => n192, ZN => 
                           N633);
   U94 : OAI21_X1 port map( B1 => n62_port, B2 => n70_port, A => n192, ZN => 
                           N634);
   U95 : OAI21_X1 port map( B1 => n61_port, B2 => n70_port, A => n192, ZN => 
                           N635);
   U96 : OAI21_X1 port map( B1 => n68_port, B2 => n71_port, A => n193, ZN => 
                           N620);
   U97 : OAI21_X1 port map( B1 => n67_port, B2 => n71_port, A => n193, ZN => 
                           N621);
   U98 : OAI21_X1 port map( B1 => n66_port, B2 => n71_port, A => n193, ZN => 
                           N622);
   U99 : OAI21_X1 port map( B1 => n65_port, B2 => n71_port, A => n193, ZN => 
                           N623);
   U100 : OAI21_X1 port map( B1 => n64_port, B2 => n71_port, A => n193, ZN => 
                           N624);
   U101 : OAI21_X1 port map( B1 => n63_port, B2 => n71_port, A => n193, ZN => 
                           N625);
   U102 : OAI21_X1 port map( B1 => n62_port, B2 => n71_port, A => n193, ZN => 
                           N626);
   U103 : OAI21_X1 port map( B1 => WRONG_PRE, B2 => n108_port, A => n192, ZN =>
                           N356);
   U104 : INV_X1 port map( A => N479, ZN => n232_port);
   U105 : NOR2_X1 port map( A1 => N480, A2 => n56_port, ZN => N644);
   U106 : NOR2_X1 port map( A1 => n57_port, A2 => n196, ZN => N645);
   U107 : AOI22_X1 port map( A1 => n173, A2 => n58_port, B1 => n59_port, B2 => 
                           n56_port, ZN => n57_port);
   U108 : OAI21_X1 port map( B1 => N480, B2 => n232_port, A => n59_port, ZN => 
                           n58_port);
   U109 : NAND2_X1 port map( A1 => N480, A2 => n232_port, ZN => n59_port);
   U110 : NAND2_X1 port map( A1 => n56_port, A2 => n73_port, ZN => n69_port);
   U111 : NAND2_X1 port map( A1 => RIGHT_PRE, A2 => N480, ZN => n73_port);
   U112 : OAI21_X1 port map( B1 => n55_port, B2 => n196, A => n56_port, ZN => 
                           SEL);
   U113 : NOR2_X1 port map( A1 => n238_port, A2 => n54_port, ZN => n55_port);
   U114 : INV_X1 port map( A => n108_port, ZN => n238_port);
   U115 : OR3_X1 port map( A1 => n186, A2 => WRONG_PRE, A3 => n54_port, ZN => 
                           N323);
   U116 : INV_X1 port map( A => n82_port, ZN => n206);
   U117 : AOI222_X1 port map( A1 => N70, A2 => n173, B1 => N105, B2 => n176, C1
                           => N243, C2 => n179, ZN => n82_port);
   U118 : INV_X1 port map( A => n81_port, ZN => n205);
   U119 : AOI222_X1 port map( A1 => N71, A2 => n173, B1 => N106, B2 => n176, C1
                           => N244, C2 => n179, ZN => n81_port);
   U120 : INV_X1 port map( A => n80, ZN => n204);
   U121 : AOI222_X1 port map( A1 => N72, A2 => n173, B1 => N107, B2 => n176, C1
                           => N245, C2 => n179, ZN => n80);
   U122 : INV_X1 port map( A => n79, ZN => n203);
   U123 : AOI222_X1 port map( A1 => N73, A2 => n173, B1 => N108, B2 => n176, C1
                           => N246, C2 => n179, ZN => n79);
   U124 : INV_X1 port map( A => n78, ZN => n202);
   U125 : AOI222_X1 port map( A1 => N74, A2 => n173, B1 => N109, B2 => n176, C1
                           => N247, C2 => n179, ZN => n78);
   U126 : INV_X1 port map( A => n77_port, ZN => n201);
   U127 : AOI222_X1 port map( A1 => N75, A2 => n173, B1 => N110, B2 => n176, C1
                           => N248, C2 => n179, ZN => n77_port);
   U128 : INV_X1 port map( A => n76_port, ZN => n200);
   U129 : AOI222_X1 port map( A1 => N76, A2 => n173, B1 => N111, B2 => n176, C1
                           => N249, C2 => n179, ZN => n76_port);
   U130 : INV_X1 port map( A => n106_port, ZN => n230_port);
   U131 : AOI222_X1 port map( A1 => N46, A2 => n171, B1 => N81, B2 => n174, C1 
                           => N219, C2 => n177, ZN => n106_port);
   U132 : INV_X1 port map( A => n105_port, ZN => n229_port);
   U133 : AOI222_X1 port map( A1 => N47, A2 => n171, B1 => N82, B2 => n174, C1 
                           => N220, C2 => n177, ZN => n105_port);
   U134 : INV_X1 port map( A => n104_port, ZN => n228_port);
   U135 : AOI222_X1 port map( A1 => N48, A2 => n171, B1 => N83, B2 => n174, C1 
                           => N221, C2 => n177, ZN => n104_port);
   U136 : INV_X1 port map( A => n103_port, ZN => n227_port);
   U137 : AOI222_X1 port map( A1 => N49, A2 => n171, B1 => N84, B2 => n174, C1 
                           => N222, C2 => n177, ZN => n103_port);
   U138 : INV_X1 port map( A => n102_port, ZN => n226_port);
   U139 : AOI222_X1 port map( A1 => N50, A2 => n171, B1 => N85, B2 => n174, C1 
                           => N223, C2 => n177, ZN => n102_port);
   U140 : INV_X1 port map( A => n101_port, ZN => n225_port);
   U141 : AOI222_X1 port map( A1 => N51, A2 => n171, B1 => N86, B2 => n174, C1 
                           => N224, C2 => n177, ZN => n101_port);
   U142 : INV_X1 port map( A => n100_port, ZN => n224_port);
   U143 : AOI222_X1 port map( A1 => N52, A2 => n171, B1 => N87, B2 => n174, C1 
                           => N225, C2 => n177, ZN => n100_port);
   U144 : INV_X1 port map( A => n99_port, ZN => n223_port);
   U145 : AOI222_X1 port map( A1 => N53, A2 => n171, B1 => N88, B2 => n174, C1 
                           => N226, C2 => n177, ZN => n99_port);
   U146 : INV_X1 port map( A => n98_port, ZN => n222_port);
   U147 : AOI222_X1 port map( A1 => N54, A2 => n171, B1 => N89, B2 => n174, C1 
                           => N227, C2 => n177, ZN => n98_port);
   U148 : INV_X1 port map( A => n97_port, ZN => n221_port);
   U149 : AOI222_X1 port map( A1 => N55, A2 => n171, B1 => N90, B2 => n174, C1 
                           => N228, C2 => n177, ZN => n97_port);
   U150 : INV_X1 port map( A => n96_port, ZN => n220_port);
   U151 : AOI222_X1 port map( A1 => N56, A2 => n171, B1 => N91, B2 => n174, C1 
                           => N229, C2 => n177, ZN => n96_port);
   U152 : INV_X1 port map( A => n95_port, ZN => n219_port);
   U153 : AOI222_X1 port map( A1 => N57, A2 => n171, B1 => N92, B2 => n174, C1 
                           => N230, C2 => n177, ZN => n95_port);
   U154 : INV_X1 port map( A => n94_port, ZN => n218);
   U155 : AOI222_X1 port map( A1 => N58, A2 => n172, B1 => N93, B2 => n175, C1 
                           => N231, C2 => n178, ZN => n94_port);
   U156 : INV_X1 port map( A => n93_port, ZN => n217);
   U157 : AOI222_X1 port map( A1 => N59, A2 => n172, B1 => N94, B2 => n175, C1 
                           => N232, C2 => n178, ZN => n93_port);
   U158 : INV_X1 port map( A => n92_port, ZN => n216_port);
   U159 : AOI222_X1 port map( A1 => N60, A2 => n172, B1 => N95, B2 => n175, C1 
                           => N233, C2 => n178, ZN => n92_port);
   U160 : INV_X1 port map( A => n91_port, ZN => n215);
   U161 : AOI222_X1 port map( A1 => N61, A2 => n172, B1 => N96, B2 => n175, C1 
                           => N234, C2 => n178, ZN => n91_port);
   U162 : INV_X1 port map( A => n90_port, ZN => n214);
   U163 : AOI222_X1 port map( A1 => N62, A2 => n172, B1 => N97, B2 => n175, C1 
                           => N235, C2 => n178, ZN => n90_port);
   U164 : INV_X1 port map( A => n89_port, ZN => n213);
   U165 : AOI222_X1 port map( A1 => N63, A2 => n172, B1 => N98, B2 => n175, C1 
                           => N236, C2 => n178, ZN => n89_port);
   U179 : INV_X1 port map( A => n88_port, ZN => n212);
   U180 : AOI222_X1 port map( A1 => N64, A2 => n172, B1 => N99, B2 => n175, C1 
                           => N237, C2 => n178, ZN => n88_port);
   U181 : INV_X1 port map( A => n87_port, ZN => n211);
   U182 : AOI222_X1 port map( A1 => N65, A2 => n172, B1 => N100, B2 => n175, C1
                           => N238, C2 => n178, ZN => n87_port);
   U183 : INV_X1 port map( A => n86_port, ZN => n210);
   U184 : AOI222_X1 port map( A1 => N66, A2 => n172, B1 => N101, B2 => n175, C1
                           => N239, C2 => n178, ZN => n86_port);
   U185 : INV_X1 port map( A => n85_port, ZN => n209);
   U186 : AOI222_X1 port map( A1 => N67, A2 => n172, B1 => N102, B2 => n175, C1
                           => N240, C2 => n178, ZN => n85_port);
   U187 : INV_X1 port map( A => n84_port, ZN => n208);
   U188 : AOI222_X1 port map( A1 => N68, A2 => n172, B1 => N103, B2 => n175, C1
                           => N241, C2 => n178, ZN => n84_port);
   U189 : INV_X1 port map( A => n83_port, ZN => n207);
   U190 : AOI222_X1 port map( A1 => N69, A2 => n172, B1 => N104, B2 => n175, C1
                           => N242, C2 => n178, ZN => n83_port);
   U191 : NOR4_X1 port map( A1 => n237_port, A2 => n239_port, A3 => N216, A4 =>
                           IR_IN(27), ZN => n54_port);
   U192 : INV_X1 port map( A => n109_port, ZN => n237_port);
   U193 : NOR3_X1 port map( A1 => IR_IN(31), A2 => IR_IN(30), A3 => IR_IN(29), 
                           ZN => n109_port);
   U194 : INV_X1 port map( A => PC_FAIL(5), ZN => n233_port);
   U195 : INV_X1 port map( A => PC_FAIL(4), ZN => n234_port);
   U196 : INV_X1 port map( A => PC_FAIL(2), ZN => n236_port);
   U197 : AND2_X1 port map( A1 => IR_FAIL(5), A2 => N479, ZN => n7);
   U198 : AND2_X1 port map( A1 => IR_FAIL(2), A2 => N479, ZN => n8);
   U199 : AND2_X1 port map( A1 => IR_FAIL(3), A2 => N479, ZN => n9);
   U200 : AND2_X1 port map( A1 => IR_FAIL(4), A2 => N479, ZN => n10);
   U201 : AND2_X1 port map( A1 => IR_FAIL(6), A2 => N479, ZN => n11);
   U202 : AND2_X1 port map( A1 => IR_FAIL(7), A2 => N479, ZN => n12);
   U203 : AND2_X1 port map( A1 => IR_FAIL(8), A2 => N479, ZN => n13);
   U204 : AND2_X1 port map( A1 => N479, A2 => IR_FAIL(9), ZN => n14);
   U205 : AND2_X1 port map( A1 => IR_FAIL(10), A2 => N479, ZN => n15);
   U206 : AND2_X1 port map( A1 => IR_FAIL(11), A2 => N479, ZN => n16);
   U207 : AND2_X1 port map( A1 => IR_FAIL(12), A2 => N479, ZN => n17);
   U208 : AND2_X1 port map( A1 => IR_FAIL(13), A2 => N479, ZN => n18);
   U209 : AND2_X1 port map( A1 => IR_FAIL(14), A2 => N479, ZN => n19);
   U210 : INV_X1 port map( A => PC_FAIL(3), ZN => n235_port);
   U211 : AND2_X1 port map( A1 => IR_FAIL(0), A2 => N479, ZN => n20);
   U212 : INV_X1 port map( A => n74_port, ZN => n199);
   U213 : AOI222_X1 port map( A1 => N77, A2 => n173, B1 => N112, B2 => n176, C1
                           => N250, C2 => n179, ZN => n74_port);
   U214 : INV_X1 port map( A => IR_IN(28), ZN => n239_port);
   U215 : AND2_X1 port map( A1 => N114, A2 => n193, ZN => N358);
   U216 : AND2_X1 port map( A1 => N115, A2 => n193, ZN => N359);
   U217 : MUX2_X1 port map( A => CACHE_mem_15_0_port, B => CACHE_mem_31_0_port,
                           S => n138_port, Z => n21);
   U218 : MUX2_X1 port map( A => CACHE_mem_7_0_port, B => CACHE_mem_23_0_port, 
                           S => n138_port, Z => n22);
   U219 : MUX2_X1 port map( A => n22, B => n21, S => PC_FAIL(5), Z => n23);
   U220 : MUX2_X1 port map( A => CACHE_mem_11_0_port, B => CACHE_mem_27_0_port,
                           S => n138_port, Z => n24);
   U221 : MUX2_X1 port map( A => CACHE_mem_3_0_port, B => CACHE_mem_19_0_port, 
                           S => n138_port, Z => n25);
   U222 : MUX2_X1 port map( A => n25, B => n24, S => PC_FAIL(5), Z => n26);
   U223 : MUX2_X1 port map( A => n26, B => n23, S => PC_FAIL(4), Z => n27);
   U224 : MUX2_X1 port map( A => CACHE_mem_14_0_port, B => CACHE_mem_30_0_port,
                           S => n138_port, Z => n28);
   U225 : MUX2_X1 port map( A => CACHE_mem_6_0_port, B => CACHE_mem_22_0_port, 
                           S => n138_port, Z => n29);
   U226 : MUX2_X1 port map( A => n29, B => n28, S => PC_FAIL(5), Z => n30);
   U227 : MUX2_X1 port map( A => CACHE_mem_10_0_port, B => CACHE_mem_26_0_port,
                           S => n138_port, Z => n31);
   U228 : MUX2_X1 port map( A => CACHE_mem_2_0_port, B => CACHE_mem_18_0_port, 
                           S => n138_port, Z => n32);
   U229 : MUX2_X1 port map( A => n32, B => n31, S => PC_FAIL(5), Z => n33);
   U230 : MUX2_X1 port map( A => n33, B => n30, S => PC_FAIL(4), Z => n34);
   U231 : MUX2_X1 port map( A => n34, B => n27, S => PC_FAIL(2), Z => n35);
   U232 : MUX2_X1 port map( A => CACHE_mem_13_0_port, B => CACHE_mem_29_0_port,
                           S => n139_port, Z => n36);
   U233 : MUX2_X1 port map( A => CACHE_mem_5_0_port, B => CACHE_mem_21_0_port, 
                           S => n139_port, Z => n37);
   U234 : MUX2_X1 port map( A => n37, B => n36, S => PC_FAIL(5), Z => n38);
   U235 : MUX2_X1 port map( A => CACHE_mem_9_0_port, B => CACHE_mem_25_0_port, 
                           S => n139_port, Z => n39);
   U236 : MUX2_X1 port map( A => CACHE_mem_1_0_port, B => CACHE_mem_17_0_port, 
                           S => n139_port, Z => n40);
   U237 : MUX2_X1 port map( A => n40, B => n39, S => PC_FAIL(5), Z => n41);
   U238 : MUX2_X1 port map( A => n41, B => n38, S => PC_FAIL(4), Z => n42);
   U239 : MUX2_X1 port map( A => CACHE_mem_12_0_port, B => CACHE_mem_28_0_port,
                           S => n139_port, Z => n43);
   U240 : MUX2_X1 port map( A => CACHE_mem_4_0_port, B => CACHE_mem_20_0_port, 
                           S => n139_port, Z => n44);
   U241 : MUX2_X1 port map( A => n44, B => n43, S => PC_FAIL(5), Z => n45);
   U242 : MUX2_X1 port map( A => CACHE_mem_8_0_port, B => CACHE_mem_24_0_port, 
                           S => n139_port, Z => n46_port);
   U243 : MUX2_X1 port map( A => CACHE_mem_0_0_port, B => CACHE_mem_16_0_port, 
                           S => n139_port, Z => n47_port);
   U244 : MUX2_X1 port map( A => n47_port, B => n46_port, S => PC_FAIL(5), Z =>
                           n48_port);
   U245 : MUX2_X1 port map( A => n48_port, B => n45, S => PC_FAIL(4), Z => 
                           n49_port);
   U246 : MUX2_X1 port map( A => n49_port, B => n42, S => PC_FAIL(2), Z => 
                           n50_port);
   U247 : MUX2_X1 port map( A => n50_port, B => n35, S => PC_FAIL(3), Z => N480
                           );
   U248 : MUX2_X1 port map( A => CACHE_mem_15_1_port, B => CACHE_mem_31_1_port,
                           S => n139_port, Z => n51_port);
   U249 : MUX2_X1 port map( A => CACHE_mem_7_1_port, B => CACHE_mem_23_1_port, 
                           S => n139_port, Z => n52_port);
   U250 : MUX2_X1 port map( A => n52_port, B => n51_port, S => PC_FAIL(5), Z =>
                           n110_port);
   U251 : MUX2_X1 port map( A => CACHE_mem_11_1_port, B => CACHE_mem_27_1_port,
                           S => n139_port, Z => n111_port);
   U252 : MUX2_X1 port map( A => CACHE_mem_3_1_port, B => CACHE_mem_19_1_port, 
                           S => n139_port, Z => n112_port);
   U253 : MUX2_X1 port map( A => n112_port, B => n111_port, S => PC_FAIL(5), Z 
                           => n113_port);
   U254 : MUX2_X1 port map( A => n113_port, B => n110_port, S => PC_FAIL(4), Z 
                           => n114_port);
   U255 : MUX2_X1 port map( A => CACHE_mem_14_1_port, B => CACHE_mem_30_1_port,
                           S => n140_port, Z => n115_port);
   U256 : MUX2_X1 port map( A => CACHE_mem_6_1_port, B => CACHE_mem_22_1_port, 
                           S => n140_port, Z => n116_port);
   U257 : MUX2_X1 port map( A => n116_port, B => n115_port, S => PC_FAIL(5), Z 
                           => n117_port);
   U258 : MUX2_X1 port map( A => CACHE_mem_10_1_port, B => CACHE_mem_26_1_port,
                           S => n140_port, Z => n118_port);
   U259 : MUX2_X1 port map( A => CACHE_mem_2_1_port, B => CACHE_mem_18_1_port, 
                           S => n140_port, Z => n119_port);
   U260 : MUX2_X1 port map( A => n119_port, B => n118_port, S => PC_FAIL(5), Z 
                           => n120_port);
   U261 : MUX2_X1 port map( A => n120_port, B => n117_port, S => PC_FAIL(4), Z 
                           => n121_port);
   U262 : MUX2_X1 port map( A => n121_port, B => n114_port, S => PC_FAIL(2), Z 
                           => n122_port);
   U263 : MUX2_X1 port map( A => CACHE_mem_13_1_port, B => CACHE_mem_29_1_port,
                           S => n140_port, Z => n123_port);
   U264 : MUX2_X1 port map( A => CACHE_mem_5_1_port, B => CACHE_mem_21_1_port, 
                           S => n140_port, Z => n124_port);
   U265 : MUX2_X1 port map( A => n124_port, B => n123_port, S => PC_FAIL(5), Z 
                           => n125_port);
   U266 : MUX2_X1 port map( A => CACHE_mem_9_1_port, B => CACHE_mem_25_1_port, 
                           S => n140_port, Z => n126_port);
   U267 : MUX2_X1 port map( A => CACHE_mem_1_1_port, B => CACHE_mem_17_1_port, 
                           S => n140_port, Z => n127_port);
   U268 : MUX2_X1 port map( A => n127_port, B => n126_port, S => PC_FAIL(5), Z 
                           => n128_port);
   U269 : MUX2_X1 port map( A => n128_port, B => n125_port, S => PC_FAIL(4), Z 
                           => n129_port);
   U270 : MUX2_X1 port map( A => CACHE_mem_12_1_port, B => CACHE_mem_28_1_port,
                           S => n140_port, Z => n130_port);
   U271 : MUX2_X1 port map( A => CACHE_mem_4_1_port, B => CACHE_mem_20_1_port, 
                           S => n140_port, Z => n131_port);
   U272 : MUX2_X1 port map( A => n131_port, B => n130_port, S => PC_FAIL(5), Z 
                           => n132_port);
   U273 : MUX2_X1 port map( A => CACHE_mem_8_1_port, B => CACHE_mem_24_1_port, 
                           S => n140_port, Z => n133_port);
   U274 : MUX2_X1 port map( A => CACHE_mem_0_1_port, B => CACHE_mem_16_1_port, 
                           S => n140_port, Z => n134_port);
   U275 : MUX2_X1 port map( A => n134_port, B => n133_port, S => PC_FAIL(5), Z 
                           => n135_port);
   U276 : MUX2_X1 port map( A => n135_port, B => n132_port, S => PC_FAIL(4), Z 
                           => n136_port);
   U277 : MUX2_X1 port map( A => n136_port, B => n129_port, S => PC_FAIL(2), Z 
                           => n137_port);
   U278 : MUX2_X1 port map( A => n137_port, B => n122_port, S => PC_FAIL(3), Z 
                           => N479);
   U279 : MUX2_X1 port map( A => CACHE_mem_15_1_port, B => CACHE_mem_31_1_port,
                           S => PC_IN(6), Z => n141_port);
   U280 : MUX2_X1 port map( A => CACHE_mem_7_1_port, B => CACHE_mem_23_1_port, 
                           S => PC_IN(6), Z => n142_port);
   U281 : MUX2_X1 port map( A => n142_port, B => n141_port, S => PC_IN(5), Z =>
                           n143_port);
   U282 : MUX2_X1 port map( A => CACHE_mem_11_1_port, B => CACHE_mem_27_1_port,
                           S => PC_IN(6), Z => n144_port);
   U283 : MUX2_X1 port map( A => CACHE_mem_3_1_port, B => CACHE_mem_19_1_port, 
                           S => PC_IN(6), Z => n145);
   U284 : MUX2_X1 port map( A => n145, B => n144_port, S => PC_IN(5), Z => n146
                           );
   U285 : MUX2_X1 port map( A => n146, B => n143_port, S => PC_IN(4), Z => n147
                           );
   U286 : MUX2_X1 port map( A => CACHE_mem_14_1_port, B => CACHE_mem_30_1_port,
                           S => PC_IN(6), Z => n148);
   U287 : MUX2_X1 port map( A => CACHE_mem_6_1_port, B => CACHE_mem_22_1_port, 
                           S => PC_IN(6), Z => n149);
   U288 : MUX2_X1 port map( A => n149, B => n148, S => PC_IN(5), Z => n150);
   U289 : MUX2_X1 port map( A => CACHE_mem_10_1_port, B => CACHE_mem_26_1_port,
                           S => PC_IN(6), Z => n151);
   U290 : MUX2_X1 port map( A => CACHE_mem_2_1_port, B => CACHE_mem_18_1_port, 
                           S => PC_IN(6), Z => n152);
   U291 : MUX2_X1 port map( A => n152, B => n151, S => PC_IN(5), Z => n153);
   U292 : MUX2_X1 port map( A => n153, B => n150, S => PC_IN(4), Z => n154);
   U293 : MUX2_X1 port map( A => n154, B => n147, S => PC_IN(2), Z => n155);
   U294 : MUX2_X1 port map( A => CACHE_mem_13_1_port, B => CACHE_mem_29_1_port,
                           S => PC_IN(6), Z => n156);
   U295 : MUX2_X1 port map( A => CACHE_mem_5_1_port, B => CACHE_mem_21_1_port, 
                           S => PC_IN(6), Z => n157);
   U296 : MUX2_X1 port map( A => n157, B => n156, S => PC_IN(5), Z => n158);
   U297 : MUX2_X1 port map( A => CACHE_mem_9_1_port, B => CACHE_mem_25_1_port, 
                           S => PC_IN(6), Z => n159);
   U298 : MUX2_X1 port map( A => CACHE_mem_1_1_port, B => CACHE_mem_17_1_port, 
                           S => PC_IN(6), Z => n160);
   U299 : MUX2_X1 port map( A => n160, B => n159, S => PC_IN(5), Z => n161);
   U300 : MUX2_X1 port map( A => n161, B => n158, S => PC_IN(4), Z => n162);
   U301 : MUX2_X1 port map( A => CACHE_mem_12_1_port, B => CACHE_mem_28_1_port,
                           S => PC_IN(6), Z => n163);
   U302 : MUX2_X1 port map( A => CACHE_mem_4_1_port, B => CACHE_mem_20_1_port, 
                           S => PC_IN(6), Z => n164);
   U303 : MUX2_X1 port map( A => n164, B => n163, S => PC_IN(5), Z => n165);
   U304 : MUX2_X1 port map( A => CACHE_mem_8_1_port, B => CACHE_mem_24_1_port, 
                           S => PC_IN(6), Z => n166);
   U305 : MUX2_X1 port map( A => CACHE_mem_0_1_port, B => CACHE_mem_16_1_port, 
                           S => PC_IN(6), Z => n167);
   U306 : MUX2_X1 port map( A => n167, B => n166, S => PC_IN(5), Z => n168);
   U307 : MUX2_X1 port map( A => n168, B => n165, S => PC_IN(4), Z => n169);
   U308 : MUX2_X1 port map( A => n169, B => n162, S => PC_IN(2), Z => n170);
   U309 : MUX2_X1 port map( A => n170, B => n155, S => PC_IN(3), Z => N216);
   U310 : AND2_X1 port map( A1 => N113, A2 => n194, ZN => N357);
   U311 : INV_X1 port map( A => PC_FAIL(6), ZN => n191);
   U312 : INV_X1 port map( A => RST, ZN => n196);
   U313 : INV_X1 port map( A => RST, ZN => n197);
   U314 : INV_X1 port map( A => RST, ZN => n198);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity register_e_N32 is

   port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  O : 
         out std_logic_vector (31 downto 0));

end register_e_N32;

architecture SYN_Behavioral of register_e_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, n1, n2_port, n3_port, n_1724, n_1725, n_1726, n_1727, n_1728,
      n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, 
      n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, 
      n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755 : 
      std_logic;

begin
   
   O_reg_10_inst : DFF_X1 port map( D => N12, CK => clk, Q => O(10), QN => 
                           n_1724);
   O_reg_9_inst : DFF_X1 port map( D => N11, CK => clk, Q => O(9), QN => n_1725
                           );
   O_reg_4_inst : DFF_X1 port map( D => N6, CK => clk, Q => O(4), QN => n_1726)
                           ;
   O_reg_8_inst : DFF_X1 port map( D => N10, CK => clk, Q => O(8), QN => n_1727
                           );
   O_reg_15_inst : DFF_X1 port map( D => N17, CK => clk, Q => O(15), QN => 
                           n_1728);
   O_reg_14_inst : DFF_X1 port map( D => N16, CK => clk, Q => O(14), QN => 
                           n_1729);
   O_reg_13_inst : DFF_X1 port map( D => N15, CK => clk, Q => O(13), QN => 
                           n_1730);
   O_reg_3_inst : DFF_X1 port map( D => N5, CK => clk, Q => O(3), QN => n_1731)
                           ;
   O_reg_12_inst : DFF_X1 port map( D => N14, CK => clk, Q => O(12), QN => 
                           n_1732);
   O_reg_28_inst : DFF_X1 port map( D => N30, CK => clk, Q => O(28), QN => 
                           n_1733);
   O_reg_7_inst : DFF_X1 port map( D => N9, CK => clk, Q => O(7), QN => n_1734)
                           ;
   O_reg_1_inst : DFF_X1 port map( D => N3, CK => clk, Q => O(1), QN => n_1735)
                           ;
   O_reg_6_inst : DFF_X1 port map( D => N8, CK => clk, Q => O(6), QN => n_1736)
                           ;
   O_reg_5_inst : DFF_X1 port map( D => N7, CK => clk, Q => O(5), QN => n_1737)
                           ;
   O_reg_22_inst : DFF_X1 port map( D => N24, CK => clk, Q => O(22), QN => 
                           n_1738);
   O_reg_21_inst : DFF_X1 port map( D => N23, CK => clk, Q => O(21), QN => 
                           n_1739);
   O_reg_20_inst : DFF_X1 port map( D => N22, CK => clk, Q => O(20), QN => 
                           n_1740);
   O_reg_11_inst : DFF_X1 port map( D => N13, CK => clk, Q => O(11), QN => 
                           n_1741);
   O_reg_16_inst : DFF_X1 port map( D => N18, CK => clk, Q => O(16), QN => 
                           n_1742);
   O_reg_0_inst : DFF_X1 port map( D => N2, CK => clk, Q => O(0), QN => n_1743)
                           ;
   O_reg_2_inst : DFF_X1 port map( D => N4, CK => clk, Q => O(2), QN => n_1744)
                           ;
   O_reg_19_inst : DFF_X1 port map( D => N21, CK => clk, Q => O(19), QN => 
                           n_1745);
   O_reg_18_inst : DFF_X1 port map( D => N20, CK => clk, Q => O(18), QN => 
                           n_1746);
   O_reg_17_inst : DFF_X1 port map( D => N19, CK => clk, Q => O(17), QN => 
                           n_1747);
   O_reg_30_inst : DFF_X1 port map( D => N32, CK => clk, Q => O(30), QN => 
                           n_1748);
   O_reg_29_inst : DFF_X1 port map( D => N31, CK => clk, Q => O(29), QN => 
                           n_1749);
   O_reg_23_inst : DFF_X1 port map( D => N25, CK => clk, Q => O(23), QN => 
                           n_1750);
   O_reg_26_inst : DFF_X1 port map( D => N28, CK => clk, Q => O(26), QN => 
                           n_1751);
   O_reg_25_inst : DFF_X1 port map( D => N27, CK => clk, Q => O(25), QN => 
                           n_1752);
   O_reg_24_inst : DFF_X1 port map( D => N26, CK => clk, Q => O(24), QN => 
                           n_1753);
   O_reg_31_inst : DFF_X1 port map( D => N33, CK => clk, Q => O(31), QN => 
                           n_1754);
   O_reg_27_inst : DFF_X1 port map( D => N29, CK => clk, Q => O(27), QN => 
                           n_1755);
   U3 : BUF_X1 port map( A => rst, Z => n1);
   U4 : BUF_X1 port map( A => rst, Z => n2_port);
   U5 : BUF_X1 port map( A => rst, Z => n3_port);
   U6 : AND2_X1 port map( A1 => D(9), A2 => n1, ZN => N11);
   U7 : AND2_X1 port map( A1 => D(8), A2 => n1, ZN => N10);
   U8 : AND2_X1 port map( A1 => D(10), A2 => n1, ZN => N12);
   U9 : AND2_X1 port map( A1 => D(11), A2 => n1, ZN => N13);
   U10 : AND2_X1 port map( A1 => n1, A2 => D(7), ZN => N9);
   U11 : AND2_X1 port map( A1 => D(6), A2 => n1, ZN => N8);
   U12 : AND2_X1 port map( A1 => D(4), A2 => n1, ZN => N6);
   U13 : AND2_X1 port map( A1 => D(5), A2 => n1, ZN => N7);
   U14 : AND2_X1 port map( A1 => D(1), A2 => n1, ZN => N3);
   U15 : AND2_X1 port map( A1 => D(2), A2 => n1, ZN => N4);
   U16 : AND2_X1 port map( A1 => D(3), A2 => n1, ZN => N5);
   U17 : AND2_X1 port map( A1 => D(0), A2 => n2_port, ZN => N2);
   U18 : AND2_X1 port map( A1 => D(12), A2 => n1, ZN => N14);
   U19 : AND2_X1 port map( A1 => D(13), A2 => n3_port, ZN => N15);
   U20 : AND2_X1 port map( A1 => D(14), A2 => n3_port, ZN => N16);
   U21 : AND2_X1 port map( A1 => D(15), A2 => n3_port, ZN => N17);
   U22 : AND2_X1 port map( A1 => D(16), A2 => n3_port, ZN => N18);
   U23 : AND2_X1 port map( A1 => D(17), A2 => n2_port, ZN => N19);
   U24 : AND2_X1 port map( A1 => D(18), A2 => n2_port, ZN => N20);
   U25 : AND2_X1 port map( A1 => D(19), A2 => n2_port, ZN => N21);
   U26 : AND2_X1 port map( A1 => D(20), A2 => n2_port, ZN => N22);
   U27 : AND2_X1 port map( A1 => D(21), A2 => n2_port, ZN => N23);
   U28 : AND2_X1 port map( A1 => D(22), A2 => n2_port, ZN => N24);
   U29 : AND2_X1 port map( A1 => D(23), A2 => n2_port, ZN => N25);
   U30 : AND2_X1 port map( A1 => D(24), A2 => n2_port, ZN => N26);
   U31 : AND2_X1 port map( A1 => D(25), A2 => n2_port, ZN => N27);
   U32 : AND2_X1 port map( A1 => D(26), A2 => n2_port, ZN => N28);
   U33 : AND2_X1 port map( A1 => D(27), A2 => n2_port, ZN => N29);
   U34 : AND2_X1 port map( A1 => D(28), A2 => n2_port, ZN => N30);
   U35 : AND2_X1 port map( A1 => D(29), A2 => n2_port, ZN => N31);
   U36 : AND2_X1 port map( A1 => D(30), A2 => n2_port, ZN => N32);
   U37 : AND2_X1 port map( A1 => D(31), A2 => n2_port, ZN => N33);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity MUX21_GENERIC_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_N32_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n43, n54, n63, n64, n1, n2, n3, n4
      , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n41
      , n42, n44, n45, n46, n47, n48, n49 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n49);
   U2 : INV_X1 port map( A => n49, ZN => n32);
   U3 : INV_X1 port map( A => n49, ZN => n29);
   U4 : INV_X1 port map( A => n49, ZN => n7);
   U5 : INV_X1 port map( A => n49, ZN => n10);
   U6 : INV_X1 port map( A => n49, ZN => n26);
   U7 : INV_X1 port map( A => n49, ZN => n23);
   U8 : INV_X1 port map( A => n49, ZN => n20);
   U9 : NAND2_X1 port map( A1 => B(31), A2 => n49, ZN => n15);
   U10 : INV_X1 port map( A => n47, ZN => n4);
   U11 : INV_X1 port map( A => SEL, ZN => n47);
   U12 : INV_X1 port map( A => SEL, ZN => n46);
   U13 : NAND2_X1 port map( A1 => A(0), A2 => n1, ZN => n2);
   U14 : NAND2_X1 port map( A1 => B(0), A2 => n49, ZN => n3);
   U15 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Y(0));
   U16 : INV_X1 port map( A => n49, ZN => n1);
   U17 : NAND2_X1 port map( A1 => A(22), A2 => n4, ZN => n5);
   U18 : NAND2_X1 port map( A1 => B(22), A2 => n47, ZN => n6);
   U19 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Y(22));
   U20 : NAND2_X1 port map( A1 => A(26), A2 => n7, ZN => n8);
   U21 : NAND2_X1 port map( A1 => B(26), A2 => n49, ZN => n9);
   U22 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => Y(26));
   U23 : NAND2_X1 port map( A1 => A(23), A2 => n10, ZN => n11);
   U24 : NAND2_X1 port map( A1 => B(23), A2 => n49, ZN => n12);
   U25 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Y(23));
   U26 : NAND2_X1 port map( A1 => A(31), A2 => n13, ZN => n14);
   U27 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(31));
   U28 : INV_X1 port map( A => n49, ZN => n13);
   U29 : NAND2_X1 port map( A1 => A(30), A2 => n4, ZN => n16);
   U30 : NAND2_X1 port map( A1 => B(30), A2 => n46, ZN => n17);
   U31 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(30));
   U32 : NAND2_X1 port map( A1 => A(29), A2 => n42, ZN => n18);
   U33 : NAND2_X1 port map( A1 => B(29), A2 => n47, ZN => n19);
   U34 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(29));
   U35 : NAND2_X1 port map( A1 => A(28), A2 => n20, ZN => n21);
   U36 : NAND2_X1 port map( A1 => B(28), A2 => n49, ZN => n22);
   U37 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => Y(28));
   U38 : NAND2_X1 port map( A1 => A(21), A2 => n23, ZN => n24);
   U39 : NAND2_X1 port map( A1 => B(21), A2 => n49, ZN => n25);
   U40 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(21));
   U41 : NAND2_X1 port map( A1 => A(20), A2 => n26, ZN => n27);
   U42 : NAND2_X1 port map( A1 => B(20), A2 => n49, ZN => n28);
   U43 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => Y(20));
   U44 : NAND2_X1 port map( A1 => A(25), A2 => n29, ZN => n30);
   U45 : NAND2_X1 port map( A1 => B(25), A2 => n49, ZN => n31);
   U46 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(25));
   U47 : NAND2_X1 port map( A1 => A(24), A2 => n32, ZN => n33);
   U48 : NAND2_X1 port map( A1 => B(24), A2 => n49, ZN => n41);
   U49 : NAND2_X1 port map( A1 => n33, A2 => n41, ZN => Y(24));
   U50 : MUX2_X1 port map( A => A(27), B => B(27), S => n49, Z => Y(27));
   U51 : INV_X1 port map( A => n49, ZN => n44);
   U52 : INV_X1 port map( A => n48, ZN => n42);
   U53 : INV_X1 port map( A => n34, ZN => Y(9));
   U54 : AOI22_X1 port map( A1 => n42, A2 => A(9), B1 => B(9), B2 => n48, ZN =>
                           n34);
   U55 : INV_X1 port map( A => n35, ZN => Y(8));
   U56 : AOI22_X1 port map( A1 => A(8), A2 => n42, B1 => B(8), B2 => n47, ZN =>
                           n35);
   U57 : INV_X1 port map( A => n64, ZN => Y(10));
   U58 : AOI22_X1 port map( A1 => A(10), A2 => n42, B1 => B(10), B2 => n46, ZN 
                           => n64);
   U59 : INV_X1 port map( A => n63, ZN => Y(11));
   U60 : AOI22_X1 port map( A1 => A(11), A2 => n42, B1 => B(11), B2 => n48, ZN 
                           => n63);
   U61 : INV_X1 port map( A => n36, ZN => Y(7));
   U62 : AOI22_X1 port map( A1 => A(7), A2 => n42, B1 => B(7), B2 => n47, ZN =>
                           n36);
   U63 : INV_X1 port map( A => n37, ZN => Y(6));
   U64 : AOI22_X1 port map( A1 => A(6), A2 => n42, B1 => B(6), B2 => n47, ZN =>
                           n37);
   U65 : INV_X1 port map( A => n39, ZN => Y(4));
   U66 : AOI22_X1 port map( A1 => A(4), A2 => n42, B1 => B(4), B2 => n46, ZN =>
                           n39);
   U67 : INV_X1 port map( A => n38, ZN => Y(5));
   U68 : AOI22_X1 port map( A1 => A(5), A2 => n42, B1 => B(5), B2 => n46, ZN =>
                           n38);
   U69 : INV_X1 port map( A => n54, ZN => Y(1));
   U70 : AOI22_X1 port map( A1 => A(1), A2 => n42, B1 => B(1), B2 => n48, ZN =>
                           n54);
   U71 : INV_X1 port map( A => n43, ZN => Y(2));
   U72 : AOI22_X1 port map( A1 => A(2), A2 => n42, B1 => B(2), B2 => n47, ZN =>
                           n43);
   U73 : INV_X1 port map( A => n40, ZN => Y(3));
   U74 : AOI22_X1 port map( A1 => A(3), A2 => n42, B1 => B(3), B2 => n46, ZN =>
                           n40);
   U75 : INV_X1 port map( A => n49, ZN => n45);
   U76 : INV_X1 port map( A => SEL, ZN => n48);
   U77 : MUX2_X1 port map( A => B(12), B => A(12), S => n42, Z => Y(12));
   U78 : MUX2_X1 port map( A => B(13), B => A(13), S => n45, Z => Y(13));
   U79 : MUX2_X1 port map( A => B(14), B => A(14), S => n45, Z => Y(14));
   U80 : MUX2_X1 port map( A => B(15), B => A(15), S => n44, Z => Y(15));
   U81 : MUX2_X1 port map( A => B(16), B => A(16), S => n44, Z => Y(16));
   U82 : MUX2_X1 port map( A => B(17), B => A(17), S => n44, Z => Y(17));
   U83 : MUX2_X1 port map( A => B(18), B => A(18), S => n44, Z => Y(18));
   U84 : MUX2_X1 port map( A => B(19), B => A(19), S => n44, Z => Y(19));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity DPATH is

   port( Clk, Rst, MUXA_SEL, MUXB_SEL, BR_EN : in std_logic;  ALU_OPCODE : in 
         std_logic_vector (0 to 4);  WB_MUX_SEL : in std_logic_vector (1 downto
         0);  RF_WE : in std_logic;  DRAM_OUT, IRAM_OUT : in std_logic_vector 
         (31 downto 0);  IR1, DRAM_IN : out std_logic_vector (31 downto 0);  
         DRAM_ADD : out std_logic_vector (11 downto 0);  IR_ADD : out 
         std_logic_vector (7 downto 0));

end DPATH;

architecture SYN_STRUCTURAL of DPATH is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux_3to1_N32_1
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MEM_WB
      port( CLK, RST : in std_logic;  NPC_L_IN, ALU_IN, LMD_IN : in 
            std_logic_vector (31 downto 0);  RD_IN : in std_logic_vector (4 
            downto 0);  OPCODE_IN : in std_logic_vector (5 downto 0);  
            NPC_L_OUT, ALU_OUT, LMD_OUT : out std_logic_vector (31 downto 0);  
            RD_OUT : out std_logic_vector (4 downto 0);  OPCODE_OUT : out 
            std_logic_vector (5 downto 0));
   end component;
   
   component EX_MEM
      port( CLK, RST : in std_logic;  NPC_IN, NPC_L_IN, ALU_IN, B_IN : in 
            std_logic_vector (31 downto 0);  RD_IN : in std_logic_vector (4 
            downto 0);  OPCODE_IN : in std_logic_vector (5 downto 0);  NPC_OUT,
            NPC_L_OUT, ALU_OUT, B_OUT : out std_logic_vector (31 downto 0);  
            RD_OUT : out std_logic_vector (4 downto 0);  OPCODE_OUT : out 
            std_logic_vector (5 downto 0));
   end component;
   
   component branch_cond_N32
      port( A : in std_logic_vector (31 downto 0);  EN : in std_logic;  OP : in
            std_logic_vector (0 to 4);  PRE : in std_logic;  DISCARD, WRONG, 
            RIGHT, SEL : out std_logic);
   end component;
   
   component mux_3to1_N32_2
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_UNIT_BRANCH
      port( Rst : in std_logic;  Rs1, Rd_M, Rd_W : in std_logic_vector (4 
            downto 0);  ICODE, ICODE_M, ICODE_W : in std_logic_vector (5 downto
            0);  SEL : out std_logic_vector (1 downto 0));
   end component;
   
   component ALU_N32
      port( INA, INB : in std_logic_vector (31 downto 0);  OP : in 
            std_logic_vector (0 to 4);  alu_out : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux_3to1_N32_3
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux_3to1_N32_0
      port( A, B, C : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component FWD_UNIT
      port( Rst : in std_logic;  Rs1, Rs2, Rd_M, Rd_W : in std_logic_vector (4 
            downto 0);  ICODE, ICODE_M, ICODE_W : in std_logic_vector (5 downto
            0);  SEL_A, SEL_B : out std_logic_vector (1 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component ID_EX
      port( CLK, RST : in std_logic;  NPC_IN, NPC_L_IN, A_IN, B_IN, IMM_IN : in
            std_logic_vector (31 downto 0);  RS1_IN, RS2_IN, RD_IN : in 
            std_logic_vector (4 downto 0);  OPCODE_IN : in std_logic_vector (5 
            downto 0);  IR_IN : in std_logic_vector (15 downto 0);  PR_IN : in 
            std_logic;  NPC_OUT, NPC_L_OUT, A_OUT, B_OUT, IMM_OUT : out 
            std_logic_vector (31 downto 0);  RS1_OUT, RS2_OUT, RD_OUT : out 
            std_logic_vector (4 downto 0);  OPCODE_OUT : out std_logic_vector 
            (5 downto 0);  IR_OUT : out std_logic_vector (15 downto 0);  PR_OUT
            : out std_logic);
   end component;
   
   component sign_extender
      port( d_in : in std_logic_vector (31 downto 0);  rst : in std_logic;  
            d_ext : out std_logic_vector (31 downto 0));
   end component;
   
   component register_file_N32_addBit5
      port( RESET, RE, WE : in std_logic;  ADD_WR, ADD_RDA, ADD_RDB : in 
            std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
            downto 0);  OUTA, OUTB : out std_logic_vector (31 downto 0));
   end component;
   
   component IR_decoder
      port( rst : in std_logic;  IR_OUT : in std_logic_vector (20 downto 0);  
            ADDS1, ADDS2, ADDD : out std_logic_vector (4 downto 0));
   end component;
   
   component IF_ID
      port( CLK, RST, DISCARD : in std_logic;  NPC_IN, NPC_L_IN, IR_IN : in 
            std_logic_vector (31 downto 0);  PR_IN : in std_logic;  NPC_OUT, 
            NPC_L_OUT, IR_OUT : out std_logic_vector (31 downto 0);  PR_OUT : 
            out std_logic);
   end component;
   
   component NPC_adder
      port( inPC : in std_logic_vector (31 downto 0);  outPC : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component branch_predictor
      port( RST : in std_logic;  PC_IN, PC_FAIL, IR_IN : in std_logic_vector 
            (31 downto 0);  IR_FAIL : in std_logic_vector (15 downto 0);  
            WRONG_PRE, RIGHT_PRE : in std_logic;  NPC_OUT, LINK_ADD : out 
            std_logic_vector (31 downto 0);  SEL, TAKEN : out std_logic);
   end component;
   
   component register_e_N32
      port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  O
            : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, IR1_31_port, IR1_30_port, IR1_29_port, IR1_28_port, 
      IR1_27_port, IR1_26_port, IR1_25_port, IR1_24_port, IR1_23_port, 
      IR1_22_port, IR1_21_port, IR1_20_port, IR1_19_port, IR1_18_port, 
      IR1_17_port, IR1_16_port, IR1_15_port, IR1_14_port, IR1_13_port, 
      IR1_12_port, IR1_11_port, IR1_10_port, IR1_9_port, IR1_8_port, IR1_7_port
      , IR1_6_port, IR1_5_port, IR1_4_port, IR1_3_port, IR1_2_port, IR1_1_port,
      IR1_0_port, DRAM_ADD_11_port, DRAM_ADD_10_port, DRAM_ADD_9_port, 
      DRAM_ADD_8_port, DRAM_ADD_7_port, DRAM_ADD_6_port, DRAM_ADD_5_port, 
      DRAM_ADD_4_port, DRAM_ADD_3_port, DRAM_ADD_2_port, DRAM_ADD_1_port, 
      DRAM_ADD_0_port, IR_ADD_7_port, IR_ADD_6_port, IR_ADD_5_port, 
      IR_ADD_4_port, IR_ADD_3_port, IR_ADD_2_port, IR_ADD_1_port, IR_ADD_0_port
      , alu_out_31_port, alu_out_30_port, alu_out_29_port, alu_out_28_port, 
      alu_out_27_port, alu_out_26_port, alu_out_25_port, alu_out_24_port, 
      alu_out_23_port, alu_out_22_port, alu_out_21_port, alu_out_20_port, 
      alu_out_19_port, alu_out_18_port, alu_out_17_port, alu_out_16_port, 
      alu_out_15_port, alu_out_14_port, alu_out_13_port, alu_out_12_port, 
      alu_out_11_port, alu_out_10_port, alu_out_9_port, alu_out_8_port, 
      alu_out_7_port, alu_out_6_port, alu_out_5_port, alu_out_4_port, 
      alu_out_3_port, alu_out_2_port, alu_out_1_port, alu_out_0_port, 
      npc_31_port, npc_30_port, npc_29_port, npc_28_port, npc_27_port, 
      npc_26_port, npc_25_port, npc_24_port, npc_23_port, npc_22_port, 
      npc_21_port, npc_20_port, npc_19_port, npc_18_port, npc_17_port, 
      npc_16_port, npc_15_port, npc_14_port, npc_13_port, npc_12_port, 
      npc_11_port, npc_10_port, npc_9_port, npc_8_port, npc_7_port, npc_6_port,
      npc_5_port, npc_4_port, npc_3_port, npc_2_port, npc_1_port, npc_0_port, 
      jr_sel, pc_in_31_port, pc_in_30_port, pc_in_29_port, pc_in_28_port, 
      pc_in_27_port, pc_in_26_port, pc_in_25_port, pc_in_24_port, pc_in_23_port
      , pc_in_22_port, pc_in_21_port, pc_in_20_port, pc_in_19_port, 
      pc_in_18_port, pc_in_17_port, pc_in_16_port, pc_in_15_port, pc_in_14_port
      , pc_in_13_port, pc_in_12_port, pc_in_11_port, pc_in_10_port, 
      pc_in_9_port, pc_in_8_port, pc_in_7_port, pc_in_6_port, pc_in_5_port, 
      pc_in_4_port, pc_in_3_port, pc_in_2_port, pc_in_1_port, pc_in_0_port, 
      pc_out_31_port, pc_out_30_port, pc_out_29_port, pc_out_28_port, 
      pc_out_27_port, pc_out_26_port, pc_out_25_port, pc_out_24_port, 
      pc_out_23_port, pc_out_22_port, pc_out_21_port, pc_out_20_port, 
      pc_out_19_port, pc_out_18_port, pc_out_17_port, pc_out_16_port, 
      pc_out_15_port, pc_out_14_port, pc_out_13_port, pc_out_12_port, 
      pc_out_11_port, pc_out_10_port, pc_out_1, pc_out_0, npc_M_31_port, 
      npc_M_30_port, npc_M_29_port, npc_M_28_port, npc_M_27_port, npc_M_26_port
      , npc_M_25_port, npc_M_24_port, npc_M_23_port, npc_M_22_port, 
      npc_M_21_port, npc_M_20_port, npc_M_19_port, npc_M_18_port, npc_M_17_port
      , npc_M_16_port, npc_M_15_port, npc_M_14_port, npc_M_13_port, 
      npc_M_12_port, npc_M_11_port, npc_M_10_port, npc_M_9_port, npc_M_8_port, 
      npc_M_7_port, npc_M_6_port, npc_M_5_port, npc_M_4_port, npc_M_3_port, 
      npc_M_2_port, npc_M_1_port, npc_M_0_port, ir_E_15_port, ir_E_14_port, 
      ir_E_13_port, ir_E_12_port, ir_E_11_port, ir_E_10_port, ir_E_9_port, 
      ir_E_8_port, ir_E_7_port, ir_E_6_port, ir_E_5_port, ir_E_4_port, 
      ir_E_3_port, ir_E_2_port, ir_E_1_port, ir_E_0_port, wrong_br, right_br, 
      npc_pre_31_port, npc_pre_30_port, npc_pre_29_port, npc_pre_28_port, 
      npc_pre_27_port, npc_pre_26_port, npc_pre_25_port, npc_pre_24_port, 
      npc_pre_23_port, npc_pre_22_port, npc_pre_21_port, npc_pre_20_port, 
      npc_pre_19_port, npc_pre_18_port, npc_pre_17_port, npc_pre_16_port, 
      npc_pre_15_port, npc_pre_14_port, npc_pre_13_port, npc_pre_12_port, 
      npc_pre_11_port, npc_pre_10_port, npc_pre_9_port, npc_pre_8_port, 
      npc_pre_7_port, npc_pre_6_port, npc_pre_5_port, npc_pre_4_port, 
      npc_pre_3_port, npc_pre_2_port, npc_pre_1_port, npc_pre_0_port, 
      link_addr_F_31_port, link_addr_F_30_port, link_addr_F_29_port, 
      link_addr_F_28_port, link_addr_F_27_port, link_addr_F_26_port, 
      link_addr_F_25_port, link_addr_F_24_port, link_addr_F_23_port, 
      link_addr_F_22_port, link_addr_F_21_port, link_addr_F_20_port, 
      link_addr_F_19_port, link_addr_F_18_port, link_addr_F_17_port, 
      link_addr_F_16_port, link_addr_F_15_port, link_addr_F_14_port, 
      link_addr_F_13_port, link_addr_F_12_port, link_addr_F_11_port, 
      link_addr_F_10_port, link_addr_F_9_port, link_addr_F_8_port, 
      link_addr_F_7_port, link_addr_F_6_port, link_addr_F_5_port, 
      link_addr_F_4_port, link_addr_F_3_port, link_addr_F_2_port, 
      link_addr_F_1_port, link_addr_F_0_port, npc_mux_sel, prediction, 
      npc_mux_out_31_port, npc_mux_out_30_port, npc_mux_out_29_port, 
      npc_mux_out_28_port, npc_mux_out_27_port, npc_mux_out_26_port, 
      npc_mux_out_25_port, npc_mux_out_24_port, npc_mux_out_23_port, 
      npc_mux_out_22_port, npc_mux_out_21_port, npc_mux_out_20_port, 
      npc_mux_out_19_port, npc_mux_out_18_port, npc_mux_out_17_port, 
      npc_mux_out_16_port, npc_mux_out_15_port, npc_mux_out_14_port, 
      npc_mux_out_13_port, npc_mux_out_12_port, npc_mux_out_11_port, 
      npc_mux_out_10_port, npc_mux_out_9_port, npc_mux_out_8_port, 
      npc_mux_out_7_port, npc_mux_out_6_port, npc_mux_out_5_port, 
      npc_mux_out_4_port, npc_mux_out_3_port, npc_mux_out_2_port, 
      npc_mux_out_1_port, npc_mux_out_0_port, discard_s, npc_D_31_port, 
      npc_D_30_port, npc_D_29_port, npc_D_28_port, npc_D_27_port, npc_D_26_port
      , npc_D_25_port, npc_D_24_port, npc_D_23_port, npc_D_22_port, 
      npc_D_21_port, npc_D_20_port, npc_D_19_port, npc_D_18_port, npc_D_17_port
      , npc_D_16_port, npc_D_15_port, npc_D_14_port, npc_D_13_port, 
      npc_D_12_port, npc_D_11_port, npc_D_10_port, npc_D_9_port, npc_D_8_port, 
      npc_D_7_port, npc_D_6_port, npc_D_5_port, npc_D_4_port, npc_D_3_port, 
      npc_D_2_port, npc_D_1_port, npc_D_0_port, link_addr_D_31_port, 
      link_addr_D_30_port, link_addr_D_29_port, link_addr_D_28_port, 
      link_addr_D_27_port, link_addr_D_26_port, link_addr_D_25_port, 
      link_addr_D_24_port, link_addr_D_23_port, link_addr_D_22_port, 
      link_addr_D_21_port, link_addr_D_20_port, link_addr_D_19_port, 
      link_addr_D_18_port, link_addr_D_17_port, link_addr_D_16_port, 
      link_addr_D_15_port, link_addr_D_14_port, link_addr_D_13_port, 
      link_addr_D_12_port, link_addr_D_11_port, link_addr_D_10_port, 
      link_addr_D_9_port, link_addr_D_8_port, link_addr_D_7_port, 
      link_addr_D_6_port, link_addr_D_5_port, link_addr_D_4_port, 
      link_addr_D_3_port, link_addr_D_2_port, link_addr_D_1_port, 
      link_addr_D_0_port, pr_D, add_S1_4_port, add_S1_3_port, add_S1_2_port, 
      add_S1_1_port, add_S1_0_port, add_S2_4_port, add_S2_3_port, add_S2_2_port
      , add_S2_1_port, add_S2_0_port, dest_D_4_port, dest_D_3_port, 
      dest_D_2_port, dest_D_1_port, dest_D_0_port, add_D_4_port, add_D_3_port, 
      add_D_2_port, add_D_1_port, add_D_0_port, WB_31_port, WB_30_port, 
      WB_29_port, WB_28_port, WB_27_port, WB_26_port, WB_25_port, WB_24_port, 
      WB_23_port, WB_22_port, WB_21_port, WB_20_port, WB_19_port, WB_18_port, 
      WB_17_port, WB_16_port, WB_15_port, WB_14_port, WB_13_port, WB_12_port, 
      WB_11_port, WB_10_port, WB_9_port, WB_8_port, WB_7_port, WB_6_port, 
      WB_5_port, WB_4_port, WB_3_port, WB_2_port, WB_1_port, WB_0_port, 
      a_out_31_port, a_out_30_port, a_out_29_port, a_out_28_port, a_out_27_port
      , a_out_26_port, a_out_25_port, a_out_24_port, a_out_23_port, 
      a_out_22_port, a_out_21_port, a_out_20_port, a_out_19_port, a_out_18_port
      , a_out_17_port, a_out_16_port, a_out_15_port, a_out_14_port, 
      a_out_13_port, a_out_12_port, a_out_11_port, a_out_10_port, a_out_9_port,
      a_out_8_port, a_out_7_port, a_out_6_port, a_out_5_port, a_out_4_port, 
      a_out_3_port, a_out_2_port, a_out_1_port, a_out_0_port, b_out_31_port, 
      b_out_30_port, b_out_29_port, b_out_28_port, b_out_27_port, b_out_26_port
      , b_out_25_port, b_out_24_port, b_out_23_port, b_out_22_port, 
      b_out_21_port, b_out_20_port, b_out_19_port, b_out_18_port, b_out_17_port
      , b_out_16_port, b_out_15_port, b_out_14_port, b_out_13_port, 
      b_out_12_port, b_out_11_port, b_out_10_port, b_out_9_port, b_out_8_port, 
      b_out_7_port, b_out_6_port, b_out_5_port, b_out_4_port, b_out_3_port, 
      b_out_2_port, b_out_1_port, b_out_0_port, imm_out_31_port, 
      imm_out_30_port, imm_out_29_port, imm_out_28_port, imm_out_27_port, 
      imm_out_26_port, imm_out_25_port, imm_out_24_port, imm_out_23_port, 
      imm_out_22_port, imm_out_21_port, imm_out_20_port, imm_out_19_port, 
      imm_out_18_port, imm_out_17_port, imm_out_16_port, imm_out_15_port, 
      imm_out_14_port, imm_out_13_port, imm_out_12_port, imm_out_11_port, 
      imm_out_10_port, imm_out_9_port, imm_out_8_port, imm_out_7_port, 
      imm_out_6_port, imm_out_5_port, imm_out_4_port, imm_out_3_port, 
      imm_out_2_port, imm_out_1_port, imm_out_0_port, npc_E_31_port, 
      npc_E_30_port, npc_E_29_port, npc_E_28_port, npc_E_27_port, npc_E_26_port
      , npc_E_25_port, npc_E_24_port, npc_E_23_port, npc_E_22_port, 
      npc_E_21_port, npc_E_20_port, npc_E_19_port, npc_E_18_port, npc_E_17_port
      , npc_E_16_port, npc_E_15_port, npc_E_14_port, npc_E_13_port, 
      npc_E_12_port, npc_E_11_port, npc_E_10_port, npc_E_9_port, npc_E_8_port, 
      npc_E_7_port, npc_E_6_port, npc_E_5_port, npc_E_4_port, npc_E_3_port, 
      npc_E_2_port, npc_E_1_port, npc_E_0_port, link_addr_E_31_port, 
      link_addr_E_30_port, link_addr_E_29_port, link_addr_E_28_port, 
      link_addr_E_27_port, link_addr_E_26_port, link_addr_E_25_port, 
      link_addr_E_24_port, link_addr_E_23_port, link_addr_E_22_port, 
      link_addr_E_21_port, link_addr_E_20_port, link_addr_E_19_port, 
      link_addr_E_18_port, link_addr_E_17_port, link_addr_E_16_port, 
      link_addr_E_15_port, link_addr_E_14_port, link_addr_E_13_port, 
      link_addr_E_12_port, link_addr_E_11_port, link_addr_E_10_port, 
      link_addr_E_9_port, link_addr_E_8_port, link_addr_E_7_port, 
      link_addr_E_6_port, link_addr_E_5_port, link_addr_E_4_port, 
      link_addr_E_3_port, link_addr_E_2_port, link_addr_E_1_port, 
      link_addr_E_0_port, A_s_31_port, A_s_30_port, A_s_29_port, A_s_28_port, 
      A_s_27_port, A_s_26_port, A_s_25_port, A_s_24_port, A_s_23_port, 
      A_s_22_port, A_s_21_port, A_s_20_port, A_s_19_port, A_s_18_port, 
      A_s_17_port, A_s_16_port, A_s_15_port, A_s_14_port, A_s_13_port, 
      A_s_12_port, A_s_11_port, A_s_10_port, A_s_9_port, A_s_8_port, A_s_7_port
      , A_s_6_port, A_s_5_port, A_s_4_port, A_s_3_port, A_s_2_port, A_s_1_port,
      A_s_0_port, B_s_31_port, B_s_30_port, B_s_29_port, B_s_28_port, 
      B_s_27_port, B_s_26_port, B_s_25_port, B_s_24_port, B_s_23_port, 
      B_s_22_port, B_s_21_port, B_s_20_port, B_s_19_port, B_s_18_port, 
      B_s_17_port, B_s_16_port, B_s_15_port, B_s_14_port, B_s_13_port, 
      B_s_12_port, B_s_11_port, B_s_10_port, B_s_9_port, B_s_8_port, B_s_7_port
      , B_s_6_port, B_s_5_port, B_s_4_port, B_s_3_port, B_s_2_port, B_s_1_port,
      B_s_0_port, IMM_s_31_port, IMM_s_30_port, IMM_s_29_port, IMM_s_28_port, 
      IMM_s_27_port, IMM_s_26_port, IMM_s_25_port, IMM_s_24_port, IMM_s_23_port
      , IMM_s_22_port, IMM_s_21_port, IMM_s_20_port, IMM_s_19_port, 
      IMM_s_18_port, IMM_s_17_port, IMM_s_16_port, IMM_s_15_port, IMM_s_14_port
      , IMM_s_13_port, IMM_s_12_port, IMM_s_11_port, IMM_s_10_port, 
      IMM_s_9_port, IMM_s_8_port, IMM_s_7_port, IMM_s_6_port, IMM_s_5_port, 
      IMM_s_4_port, IMM_s_3_port, IMM_s_2_port, IMM_s_1_port, IMM_s_0_port, 
      Rs1_4_port, Rs1_3_port, Rs1_2_port, Rs1_1_port, Rs1_0_port, Rs2_4_port, 
      Rs2_3_port, Rs2_2_port, Rs2_1_port, Rs2_0_port, dest_E_4_port, 
      dest_E_3_port, dest_E_2_port, dest_E_1_port, dest_E_0_port, 
      opcode_E_5_port, opcode_E_4_port, opcode_E_3_port, opcode_E_2_port, 
      opcode_E_1_port, opcode_E_0_port, pr_E, mux_a_in_31_port, 
      mux_a_in_30_port, mux_a_in_29_port, mux_a_in_28_port, mux_a_in_27_port, 
      mux_a_in_26_port, mux_a_in_25_port, mux_a_in_24_port, mux_a_in_23_port, 
      mux_a_in_22_port, mux_a_in_21_port, mux_a_in_20_port, mux_a_in_19_port, 
      mux_a_in_18_port, mux_a_in_17_port, mux_a_in_16_port, mux_a_in_15_port, 
      mux_a_in_14_port, mux_a_in_13_port, mux_a_in_12_port, mux_a_in_11_port, 
      mux_a_in_10_port, mux_a_in_9_port, mux_a_in_8_port, mux_a_in_7_port, 
      mux_a_in_6_port, mux_a_in_5_port, mux_a_in_4_port, mux_a_in_3_port, 
      mux_a_in_2_port, mux_a_in_1_port, mux_a_in_0_port, mux_b_in_31_port, 
      mux_b_in_30_port, mux_b_in_29_port, mux_b_in_28_port, mux_b_in_27_port, 
      mux_b_in_26_port, mux_b_in_25_port, mux_b_in_24_port, mux_b_in_23_port, 
      mux_b_in_22_port, mux_b_in_21_port, mux_b_in_20_port, mux_b_in_19_port, 
      mux_b_in_18_port, mux_b_in_17_port, mux_b_in_16_port, mux_b_in_15_port, 
      mux_b_in_14_port, mux_b_in_13_port, mux_b_in_12_port, mux_b_in_11_port, 
      mux_b_in_10_port, mux_b_in_9_port, mux_b_in_8_port, mux_b_in_7_port, 
      mux_b_in_6_port, mux_b_in_5_port, mux_b_in_4_port, mux_b_in_3_port, 
      mux_b_in_2_port, mux_b_in_1_port, mux_b_in_0_port, dest_M_4_port, 
      dest_M_3_port, dest_M_2_port, dest_M_1_port, dest_M_0_port, 
      opcode_M_5_port, opcode_M_4_port, opcode_M_3_port, opcode_M_2_port, 
      opcode_M_1_port, opcode_M_0_port, opcode_W_5_port, opcode_W_4_port, 
      opcode_W_3_port, opcode_W_2_port, opcode_W_1_port, opcode_W_0_port, 
      FWD_MUX_A_S_1_port, FWD_MUX_A_S_0_port, FWD_MUX_B_S_1_port, 
      FWD_MUX_B_S_0_port, alu_out_M_31_port, alu_out_M_30_port, 
      alu_out_M_29_port, alu_out_M_28_port, alu_out_M_27_port, 
      alu_out_M_26_port, alu_out_M_25_port, alu_out_M_24_port, 
      alu_out_M_23_port, alu_out_M_22_port, alu_out_M_21_port, 
      alu_out_M_20_port, alu_out_M_19_port, alu_out_M_18_port, 
      alu_out_M_17_port, alu_out_M_16_port, alu_out_M_15_port, 
      alu_out_M_14_port, alu_out_M_13_port, alu_out_M_12_port, 
      alu_out_W_31_port, alu_out_W_30_port, alu_out_W_29_port, 
      alu_out_W_28_port, alu_out_W_27_port, alu_out_W_26_port, 
      alu_out_W_25_port, alu_out_W_24_port, alu_out_W_23_port, 
      alu_out_W_22_port, alu_out_W_21_port, alu_out_W_20_port, 
      alu_out_W_19_port, alu_out_W_18_port, alu_out_W_17_port, 
      alu_out_W_16_port, alu_out_W_15_port, alu_out_W_14_port, 
      alu_out_W_13_port, alu_out_W_12_port, alu_out_W_11_port, 
      alu_out_W_10_port, alu_out_W_9_port, alu_out_W_8_port, alu_out_W_7_port, 
      alu_out_W_6_port, alu_out_W_5_port, alu_out_W_4_port, alu_out_W_3_port, 
      alu_out_W_2_port, alu_out_W_1_port, alu_out_W_0_port, alu_a_in_31_port, 
      alu_a_in_30_port, alu_a_in_29_port, alu_a_in_28_port, alu_a_in_27_port, 
      alu_a_in_26_port, alu_a_in_25_port, alu_a_in_24_port, alu_a_in_23_port, 
      alu_a_in_22_port, alu_a_in_21_port, alu_a_in_20_port, alu_a_in_19_port, 
      alu_a_in_18_port, alu_a_in_17_port, alu_a_in_16_port, alu_a_in_15_port, 
      alu_a_in_14_port, alu_a_in_13_port, alu_a_in_12_port, alu_a_in_11_port, 
      alu_a_in_10_port, alu_a_in_9_port, alu_a_in_8_port, alu_a_in_7_port, 
      alu_a_in_6_port, alu_a_in_5_port, alu_a_in_4_port, alu_a_in_3_port, 
      alu_a_in_2_port, alu_a_in_1_port, alu_a_in_0_port, alu_b_in_31_port, 
      alu_b_in_30_port, alu_b_in_29_port, alu_b_in_28_port, alu_b_in_27_port, 
      alu_b_in_26_port, alu_b_in_25_port, alu_b_in_24_port, alu_b_in_23_port, 
      alu_b_in_22_port, alu_b_in_21_port, alu_b_in_20_port, alu_b_in_19_port, 
      alu_b_in_18_port, alu_b_in_17_port, alu_b_in_16_port, alu_b_in_15_port, 
      alu_b_in_14_port, alu_b_in_13_port, alu_b_in_12_port, alu_b_in_11_port, 
      alu_b_in_10_port, alu_b_in_9_port, alu_b_in_8_port, alu_b_in_7_port, 
      alu_b_in_6_port, alu_b_in_5_port, alu_b_in_4_port, alu_b_in_3_port, 
      alu_b_in_2_port, alu_b_in_1_port, alu_b_in_0_port, FWD_MUX_BR_S_1_port, 
      FWD_MUX_BR_S_0_port, br_mux_out_31_port, br_mux_out_30_port, 
      br_mux_out_29_port, br_mux_out_28_port, br_mux_out_27_port, 
      br_mux_out_26_port, br_mux_out_25_port, br_mux_out_24_port, 
      br_mux_out_23_port, br_mux_out_22_port, br_mux_out_21_port, 
      br_mux_out_20_port, br_mux_out_19_port, br_mux_out_18_port, 
      br_mux_out_17_port, br_mux_out_16_port, br_mux_out_15_port, 
      br_mux_out_14_port, br_mux_out_13_port, br_mux_out_12_port, 
      br_mux_out_11_port, br_mux_out_10_port, br_mux_out_9_port, 
      br_mux_out_8_port, br_mux_out_7_port, br_mux_out_6_port, 
      br_mux_out_5_port, br_mux_out_4_port, br_mux_out_3_port, 
      br_mux_out_2_port, br_mux_out_1_port, br_mux_out_0_port, 
      link_addr_M_31_port, link_addr_M_30_port, link_addr_M_29_port, 
      link_addr_M_28_port, link_addr_M_27_port, link_addr_M_26_port, 
      link_addr_M_25_port, link_addr_M_24_port, link_addr_M_23_port, 
      link_addr_M_22_port, link_addr_M_21_port, link_addr_M_20_port, 
      link_addr_M_19_port, link_addr_M_18_port, link_addr_M_17_port, 
      link_addr_M_16_port, link_addr_M_15_port, link_addr_M_14_port, 
      link_addr_M_13_port, link_addr_M_12_port, link_addr_M_11_port, 
      link_addr_M_10_port, link_addr_M_9_port, link_addr_M_8_port, 
      link_addr_M_7_port, link_addr_M_6_port, link_addr_M_5_port, 
      link_addr_M_4_port, link_addr_M_3_port, link_addr_M_2_port, 
      link_addr_M_1_port, link_addr_M_0_port, link_addr_W_31_port, 
      link_addr_W_30_port, link_addr_W_29_port, link_addr_W_28_port, 
      link_addr_W_27_port, link_addr_W_26_port, link_addr_W_25_port, 
      link_addr_W_24_port, link_addr_W_23_port, link_addr_W_22_port, 
      link_addr_W_21_port, link_addr_W_20_port, link_addr_W_19_port, 
      link_addr_W_18_port, link_addr_W_17_port, link_addr_W_16_port, 
      link_addr_W_15_port, link_addr_W_14_port, link_addr_W_13_port, 
      link_addr_W_12_port, link_addr_W_11_port, link_addr_W_10_port, 
      link_addr_W_9_port, link_addr_W_8_port, link_addr_W_7_port, 
      link_addr_W_6_port, link_addr_W_5_port, link_addr_W_4_port, 
      link_addr_W_3_port, link_addr_W_2_port, link_addr_W_1_port, 
      link_addr_W_0_port, LMD_out_31_port, LMD_out_30_port, LMD_out_29_port, 
      LMD_out_28_port, LMD_out_27_port, LMD_out_26_port, LMD_out_25_port, 
      LMD_out_24_port, LMD_out_23_port, LMD_out_22_port, LMD_out_21_port, 
      LMD_out_20_port, LMD_out_19_port, LMD_out_18_port, LMD_out_17_port, 
      LMD_out_16_port, LMD_out_15_port, LMD_out_14_port, LMD_out_13_port, 
      LMD_out_12_port, LMD_out_11_port, LMD_out_10_port, LMD_out_9_port, 
      LMD_out_8_port, LMD_out_7_port, LMD_out_6_port, LMD_out_5_port, 
      LMD_out_4_port, LMD_out_3_port, LMD_out_2_port, LMD_out_1_port, 
      LMD_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16 : std_logic;

begin
   IR1 <= ( IR1_31_port, IR1_30_port, IR1_29_port, IR1_28_port, IR1_27_port, 
      IR1_26_port, IR1_25_port, IR1_24_port, IR1_23_port, IR1_22_port, 
      IR1_21_port, IR1_20_port, IR1_19_port, IR1_18_port, IR1_17_port, 
      IR1_16_port, IR1_15_port, IR1_14_port, IR1_13_port, IR1_12_port, 
      IR1_11_port, IR1_10_port, IR1_9_port, IR1_8_port, IR1_7_port, IR1_6_port,
      IR1_5_port, IR1_4_port, IR1_3_port, IR1_2_port, IR1_1_port, IR1_0_port );
   DRAM_ADD <= ( DRAM_ADD_11_port, DRAM_ADD_10_port, DRAM_ADD_9_port, 
      DRAM_ADD_8_port, DRAM_ADD_7_port, DRAM_ADD_6_port, DRAM_ADD_5_port, 
      DRAM_ADD_4_port, DRAM_ADD_3_port, DRAM_ADD_2_port, DRAM_ADD_1_port, 
      DRAM_ADD_0_port );
   IR_ADD <= ( IR_ADD_7_port, IR_ADD_6_port, IR_ADD_5_port, IR_ADD_4_port, 
      IR_ADD_3_port, IR_ADD_2_port, IR_ADD_1_port, IR_ADD_0_port );
   
   X_Logic1_port <= '1';
   NPC_mux : MUX21_GENERIC_N32_0 port map( A(31) => alu_out_31_port, A(30) => 
                           alu_out_30_port, A(29) => alu_out_29_port, A(28) => 
                           alu_out_28_port, A(27) => alu_out_27_port, A(26) => 
                           alu_out_26_port, A(25) => alu_out_25_port, A(24) => 
                           alu_out_24_port, A(23) => alu_out_23_port, A(22) => 
                           alu_out_22_port, A(21) => alu_out_21_port, A(20) => 
                           alu_out_20_port, A(19) => alu_out_19_port, A(18) => 
                           alu_out_18_port, A(17) => alu_out_17_port, A(16) => 
                           alu_out_16_port, A(15) => alu_out_15_port, A(14) => 
                           alu_out_14_port, A(13) => alu_out_13_port, A(12) => 
                           alu_out_12_port, A(11) => alu_out_11_port, A(10) => 
                           alu_out_10_port, A(9) => alu_out_9_port, A(8) => 
                           alu_out_8_port, A(7) => alu_out_7_port, A(6) => 
                           alu_out_6_port, A(5) => alu_out_5_port, A(4) => 
                           alu_out_4_port, A(3) => alu_out_3_port, A(2) => 
                           alu_out_2_port, A(1) => alu_out_1_port, A(0) => 
                           alu_out_0_port, B(31) => npc_31_port, B(30) => 
                           npc_30_port, B(29) => npc_29_port, B(28) => 
                           npc_28_port, B(27) => npc_27_port, B(26) => 
                           npc_26_port, B(25) => npc_25_port, B(24) => 
                           npc_24_port, B(23) => npc_23_port, B(22) => 
                           npc_22_port, B(21) => npc_21_port, B(20) => 
                           npc_20_port, B(19) => npc_19_port, B(18) => 
                           npc_18_port, B(17) => npc_17_port, B(16) => 
                           npc_16_port, B(15) => npc_15_port, B(14) => 
                           npc_14_port, B(13) => npc_13_port, B(12) => 
                           npc_12_port, B(11) => npc_11_port, B(10) => 
                           npc_10_port, B(9) => npc_9_port, B(8) => npc_8_port,
                           B(7) => npc_7_port, B(6) => npc_6_port, B(5) => 
                           npc_5_port, B(4) => npc_4_port, B(3) => npc_3_port, 
                           B(2) => npc_2_port, B(1) => npc_1_port, B(0) => 
                           npc_0_port, SEL => jr_sel, Y(31) => pc_in_31_port, 
                           Y(30) => pc_in_30_port, Y(29) => pc_in_29_port, 
                           Y(28) => pc_in_28_port, Y(27) => pc_in_27_port, 
                           Y(26) => pc_in_26_port, Y(25) => pc_in_25_port, 
                           Y(24) => pc_in_24_port, Y(23) => pc_in_23_port, 
                           Y(22) => pc_in_22_port, Y(21) => pc_in_21_port, 
                           Y(20) => pc_in_20_port, Y(19) => pc_in_19_port, 
                           Y(18) => pc_in_18_port, Y(17) => pc_in_17_port, 
                           Y(16) => pc_in_16_port, Y(15) => pc_in_15_port, 
                           Y(14) => pc_in_14_port, Y(13) => pc_in_13_port, 
                           Y(12) => pc_in_12_port, Y(11) => pc_in_11_port, 
                           Y(10) => pc_in_10_port, Y(9) => pc_in_9_port, Y(8) 
                           => pc_in_8_port, Y(7) => pc_in_7_port, Y(6) => 
                           pc_in_6_port, Y(5) => pc_in_5_port, Y(4) => 
                           pc_in_4_port, Y(3) => pc_in_3_port, Y(2) => 
                           pc_in_2_port, Y(1) => pc_in_1_port, Y(0) => 
                           pc_in_0_port);
   PC_reg : register_e_N32 port map( D(31) => pc_in_31_port, D(30) => 
                           pc_in_30_port, D(29) => pc_in_29_port, D(28) => 
                           pc_in_28_port, D(27) => pc_in_27_port, D(26) => 
                           pc_in_26_port, D(25) => pc_in_25_port, D(24) => 
                           pc_in_24_port, D(23) => pc_in_23_port, D(22) => 
                           pc_in_22_port, D(21) => pc_in_21_port, D(20) => 
                           pc_in_20_port, D(19) => pc_in_19_port, D(18) => 
                           pc_in_18_port, D(17) => pc_in_17_port, D(16) => 
                           pc_in_16_port, D(15) => pc_in_15_port, D(14) => 
                           pc_in_14_port, D(13) => pc_in_13_port, D(12) => 
                           pc_in_12_port, D(11) => pc_in_11_port, D(10) => 
                           pc_in_10_port, D(9) => pc_in_9_port, D(8) => 
                           pc_in_8_port, D(7) => pc_in_7_port, D(6) => 
                           pc_in_6_port, D(5) => pc_in_5_port, D(4) => 
                           pc_in_4_port, D(3) => pc_in_3_port, D(2) => 
                           pc_in_2_port, D(1) => pc_in_1_port, D(0) => 
                           pc_in_0_port, clk => Clk, rst => n16, O(31) => 
                           pc_out_31_port, O(30) => pc_out_30_port, O(29) => 
                           pc_out_29_port, O(28) => pc_out_28_port, O(27) => 
                           pc_out_27_port, O(26) => pc_out_26_port, O(25) => 
                           pc_out_25_port, O(24) => pc_out_24_port, O(23) => 
                           pc_out_23_port, O(22) => pc_out_22_port, O(21) => 
                           pc_out_21_port, O(20) => pc_out_20_port, O(19) => 
                           pc_out_19_port, O(18) => pc_out_18_port, O(17) => 
                           pc_out_17_port, O(16) => pc_out_16_port, O(15) => 
                           pc_out_15_port, O(14) => pc_out_14_port, O(13) => 
                           pc_out_13_port, O(12) => pc_out_12_port, O(11) => 
                           pc_out_11_port, O(10) => pc_out_10_port, O(9) => 
                           IR_ADD_7_port, O(8) => IR_ADD_6_port, O(7) => 
                           IR_ADD_5_port, O(6) => IR_ADD_4_port, O(5) => 
                           IR_ADD_3_port, O(4) => IR_ADD_2_port, O(3) => 
                           IR_ADD_1_port, O(2) => IR_ADD_0_port, O(1) => 
                           pc_out_1, O(0) => pc_out_0);
   BR_pred : branch_predictor port map( RST => n16, PC_IN(31) => pc_out_31_port
                           , PC_IN(30) => pc_out_30_port, PC_IN(29) => 
                           pc_out_29_port, PC_IN(28) => pc_out_28_port, 
                           PC_IN(27) => pc_out_27_port, PC_IN(26) => 
                           pc_out_26_port, PC_IN(25) => pc_out_25_port, 
                           PC_IN(24) => pc_out_24_port, PC_IN(23) => 
                           pc_out_23_port, PC_IN(22) => pc_out_22_port, 
                           PC_IN(21) => pc_out_21_port, PC_IN(20) => 
                           pc_out_20_port, PC_IN(19) => pc_out_19_port, 
                           PC_IN(18) => pc_out_18_port, PC_IN(17) => 
                           pc_out_17_port, PC_IN(16) => pc_out_16_port, 
                           PC_IN(15) => pc_out_15_port, PC_IN(14) => 
                           pc_out_14_port, PC_IN(13) => pc_out_13_port, 
                           PC_IN(12) => pc_out_12_port, PC_IN(11) => 
                           pc_out_11_port, PC_IN(10) => pc_out_10_port, 
                           PC_IN(9) => IR_ADD_7_port, PC_IN(8) => IR_ADD_6_port
                           , PC_IN(7) => IR_ADD_5_port, PC_IN(6) => 
                           IR_ADD_4_port, PC_IN(5) => IR_ADD_3_port, PC_IN(4) 
                           => IR_ADD_2_port, PC_IN(3) => IR_ADD_1_port, 
                           PC_IN(2) => IR_ADD_0_port, PC_IN(1) => pc_out_1, 
                           PC_IN(0) => pc_out_0, PC_FAIL(31) => npc_M_31_port, 
                           PC_FAIL(30) => npc_M_30_port, PC_FAIL(29) => 
                           npc_M_29_port, PC_FAIL(28) => npc_M_28_port, 
                           PC_FAIL(27) => npc_M_27_port, PC_FAIL(26) => 
                           npc_M_26_port, PC_FAIL(25) => npc_M_25_port, 
                           PC_FAIL(24) => npc_M_24_port, PC_FAIL(23) => 
                           npc_M_23_port, PC_FAIL(22) => npc_M_22_port, 
                           PC_FAIL(21) => npc_M_21_port, PC_FAIL(20) => 
                           npc_M_20_port, PC_FAIL(19) => npc_M_19_port, 
                           PC_FAIL(18) => npc_M_18_port, PC_FAIL(17) => 
                           npc_M_17_port, PC_FAIL(16) => npc_M_16_port, 
                           PC_FAIL(15) => npc_M_15_port, PC_FAIL(14) => 
                           npc_M_14_port, PC_FAIL(13) => npc_M_13_port, 
                           PC_FAIL(12) => npc_M_12_port, PC_FAIL(11) => 
                           npc_M_11_port, PC_FAIL(10) => npc_M_10_port, 
                           PC_FAIL(9) => npc_M_9_port, PC_FAIL(8) => 
                           npc_M_8_port, PC_FAIL(7) => npc_M_7_port, PC_FAIL(6)
                           => npc_M_6_port, PC_FAIL(5) => npc_M_5_port, 
                           PC_FAIL(4) => npc_M_4_port, PC_FAIL(3) => 
                           npc_M_3_port, PC_FAIL(2) => npc_M_2_port, PC_FAIL(1)
                           => npc_M_1_port, PC_FAIL(0) => npc_M_0_port, 
                           IR_IN(31) => IRAM_OUT(31), IR_IN(30) => IRAM_OUT(30)
                           , IR_IN(29) => IRAM_OUT(29), IR_IN(28) => 
                           IRAM_OUT(28), IR_IN(27) => IRAM_OUT(27), IR_IN(26) 
                           => IRAM_OUT(26), IR_IN(25) => IRAM_OUT(25), 
                           IR_IN(24) => IRAM_OUT(24), IR_IN(23) => IRAM_OUT(23)
                           , IR_IN(22) => IRAM_OUT(22), IR_IN(21) => 
                           IRAM_OUT(21), IR_IN(20) => IRAM_OUT(20), IR_IN(19) 
                           => IRAM_OUT(19), IR_IN(18) => IRAM_OUT(18), 
                           IR_IN(17) => IRAM_OUT(17), IR_IN(16) => IRAM_OUT(16)
                           , IR_IN(15) => IRAM_OUT(15), IR_IN(14) => 
                           IRAM_OUT(14), IR_IN(13) => IRAM_OUT(13), IR_IN(12) 
                           => IRAM_OUT(12), IR_IN(11) => IRAM_OUT(11), 
                           IR_IN(10) => IRAM_OUT(10), IR_IN(9) => IRAM_OUT(9), 
                           IR_IN(8) => IRAM_OUT(8), IR_IN(7) => IRAM_OUT(7), 
                           IR_IN(6) => IRAM_OUT(6), IR_IN(5) => IRAM_OUT(5), 
                           IR_IN(4) => IRAM_OUT(4), IR_IN(3) => IRAM_OUT(3), 
                           IR_IN(2) => IRAM_OUT(2), IR_IN(1) => IRAM_OUT(1), 
                           IR_IN(0) => IRAM_OUT(0), IR_FAIL(15) => ir_E_15_port
                           , IR_FAIL(14) => ir_E_14_port, IR_FAIL(13) => 
                           ir_E_13_port, IR_FAIL(12) => ir_E_12_port, 
                           IR_FAIL(11) => ir_E_11_port, IR_FAIL(10) => 
                           ir_E_10_port, IR_FAIL(9) => ir_E_9_port, IR_FAIL(8) 
                           => ir_E_8_port, IR_FAIL(7) => ir_E_7_port, 
                           IR_FAIL(6) => ir_E_6_port, IR_FAIL(5) => ir_E_5_port
                           , IR_FAIL(4) => ir_E_4_port, IR_FAIL(3) => 
                           ir_E_3_port, IR_FAIL(2) => ir_E_2_port, IR_FAIL(1) 
                           => ir_E_1_port, IR_FAIL(0) => ir_E_0_port, WRONG_PRE
                           => wrong_br, RIGHT_PRE => right_br, NPC_OUT(31) => 
                           npc_pre_31_port, NPC_OUT(30) => npc_pre_30_port, 
                           NPC_OUT(29) => npc_pre_29_port, NPC_OUT(28) => 
                           npc_pre_28_port, NPC_OUT(27) => npc_pre_27_port, 
                           NPC_OUT(26) => npc_pre_26_port, NPC_OUT(25) => 
                           npc_pre_25_port, NPC_OUT(24) => npc_pre_24_port, 
                           NPC_OUT(23) => npc_pre_23_port, NPC_OUT(22) => 
                           npc_pre_22_port, NPC_OUT(21) => npc_pre_21_port, 
                           NPC_OUT(20) => npc_pre_20_port, NPC_OUT(19) => 
                           npc_pre_19_port, NPC_OUT(18) => npc_pre_18_port, 
                           NPC_OUT(17) => npc_pre_17_port, NPC_OUT(16) => 
                           npc_pre_16_port, NPC_OUT(15) => npc_pre_15_port, 
                           NPC_OUT(14) => npc_pre_14_port, NPC_OUT(13) => 
                           npc_pre_13_port, NPC_OUT(12) => npc_pre_12_port, 
                           NPC_OUT(11) => npc_pre_11_port, NPC_OUT(10) => 
                           npc_pre_10_port, NPC_OUT(9) => npc_pre_9_port, 
                           NPC_OUT(8) => npc_pre_8_port, NPC_OUT(7) => 
                           npc_pre_7_port, NPC_OUT(6) => npc_pre_6_port, 
                           NPC_OUT(5) => npc_pre_5_port, NPC_OUT(4) => 
                           npc_pre_4_port, NPC_OUT(3) => npc_pre_3_port, 
                           NPC_OUT(2) => npc_pre_2_port, NPC_OUT(1) => 
                           npc_pre_1_port, NPC_OUT(0) => npc_pre_0_port, 
                           LINK_ADD(31) => link_addr_F_31_port, LINK_ADD(30) =>
                           link_addr_F_30_port, LINK_ADD(29) => 
                           link_addr_F_29_port, LINK_ADD(28) => 
                           link_addr_F_28_port, LINK_ADD(27) => 
                           link_addr_F_27_port, LINK_ADD(26) => 
                           link_addr_F_26_port, LINK_ADD(25) => 
                           link_addr_F_25_port, LINK_ADD(24) => 
                           link_addr_F_24_port, LINK_ADD(23) => 
                           link_addr_F_23_port, LINK_ADD(22) => 
                           link_addr_F_22_port, LINK_ADD(21) => 
                           link_addr_F_21_port, LINK_ADD(20) => 
                           link_addr_F_20_port, LINK_ADD(19) => 
                           link_addr_F_19_port, LINK_ADD(18) => 
                           link_addr_F_18_port, LINK_ADD(17) => 
                           link_addr_F_17_port, LINK_ADD(16) => 
                           link_addr_F_16_port, LINK_ADD(15) => 
                           link_addr_F_15_port, LINK_ADD(14) => 
                           link_addr_F_14_port, LINK_ADD(13) => 
                           link_addr_F_13_port, LINK_ADD(12) => 
                           link_addr_F_12_port, LINK_ADD(11) => 
                           link_addr_F_11_port, LINK_ADD(10) => 
                           link_addr_F_10_port, LINK_ADD(9) => 
                           link_addr_F_9_port, LINK_ADD(8) => 
                           link_addr_F_8_port, LINK_ADD(7) => 
                           link_addr_F_7_port, LINK_ADD(6) => 
                           link_addr_F_6_port, LINK_ADD(5) => 
                           link_addr_F_5_port, LINK_ADD(4) => 
                           link_addr_F_4_port, LINK_ADD(3) => 
                           link_addr_F_3_port, LINK_ADD(2) => 
                           link_addr_F_2_port, LINK_ADD(1) => 
                           link_addr_F_1_port, LINK_ADD(0) => 
                           link_addr_F_0_port, SEL => npc_mux_sel, TAKEN => 
                           prediction);
   NPC_add_mux : MUX21_GENERIC_N32_3 port map( A(31) => npc_pre_31_port, A(30) 
                           => npc_pre_30_port, A(29) => npc_pre_29_port, A(28) 
                           => npc_pre_28_port, A(27) => npc_pre_27_port, A(26) 
                           => npc_pre_26_port, A(25) => npc_pre_25_port, A(24) 
                           => npc_pre_24_port, A(23) => npc_pre_23_port, A(22) 
                           => npc_pre_22_port, A(21) => npc_pre_21_port, A(20) 
                           => npc_pre_20_port, A(19) => npc_pre_19_port, A(18) 
                           => npc_pre_18_port, A(17) => npc_pre_17_port, A(16) 
                           => npc_pre_16_port, A(15) => npc_pre_15_port, A(14) 
                           => npc_pre_14_port, A(13) => npc_pre_13_port, A(12) 
                           => npc_pre_12_port, A(11) => npc_pre_11_port, A(10) 
                           => npc_pre_10_port, A(9) => npc_pre_9_port, A(8) => 
                           npc_pre_8_port, A(7) => npc_pre_7_port, A(6) => 
                           npc_pre_6_port, A(5) => npc_pre_5_port, A(4) => 
                           npc_pre_4_port, A(3) => npc_pre_3_port, A(2) => 
                           npc_pre_2_port, A(1) => npc_pre_1_port, A(0) => 
                           npc_pre_0_port, B(31) => pc_out_31_port, B(30) => 
                           pc_out_30_port, B(29) => pc_out_29_port, B(28) => 
                           pc_out_28_port, B(27) => pc_out_27_port, B(26) => 
                           pc_out_26_port, B(25) => pc_out_25_port, B(24) => 
                           pc_out_24_port, B(23) => pc_out_23_port, B(22) => 
                           pc_out_22_port, B(21) => pc_out_21_port, B(20) => 
                           pc_out_20_port, B(19) => pc_out_19_port, B(18) => 
                           pc_out_18_port, B(17) => pc_out_17_port, B(16) => 
                           pc_out_16_port, B(15) => pc_out_15_port, B(14) => 
                           pc_out_14_port, B(13) => pc_out_13_port, B(12) => 
                           pc_out_12_port, B(11) => pc_out_11_port, B(10) => 
                           pc_out_10_port, B(9) => IR_ADD_7_port, B(8) => 
                           IR_ADD_6_port, B(7) => IR_ADD_5_port, B(6) => 
                           IR_ADD_4_port, B(5) => IR_ADD_3_port, B(4) => 
                           IR_ADD_2_port, B(3) => IR_ADD_1_port, B(2) => 
                           IR_ADD_0_port, B(1) => pc_out_1, B(0) => pc_out_0, 
                           SEL => npc_mux_sel, Y(31) => npc_mux_out_31_port, 
                           Y(30) => npc_mux_out_30_port, Y(29) => 
                           npc_mux_out_29_port, Y(28) => npc_mux_out_28_port, 
                           Y(27) => npc_mux_out_27_port, Y(26) => 
                           npc_mux_out_26_port, Y(25) => npc_mux_out_25_port, 
                           Y(24) => npc_mux_out_24_port, Y(23) => 
                           npc_mux_out_23_port, Y(22) => npc_mux_out_22_port, 
                           Y(21) => npc_mux_out_21_port, Y(20) => 
                           npc_mux_out_20_port, Y(19) => npc_mux_out_19_port, 
                           Y(18) => npc_mux_out_18_port, Y(17) => 
                           npc_mux_out_17_port, Y(16) => npc_mux_out_16_port, 
                           Y(15) => npc_mux_out_15_port, Y(14) => 
                           npc_mux_out_14_port, Y(13) => npc_mux_out_13_port, 
                           Y(12) => npc_mux_out_12_port, Y(11) => 
                           npc_mux_out_11_port, Y(10) => npc_mux_out_10_port, 
                           Y(9) => npc_mux_out_9_port, Y(8) => 
                           npc_mux_out_8_port, Y(7) => npc_mux_out_7_port, Y(6)
                           => npc_mux_out_6_port, Y(5) => npc_mux_out_5_port, 
                           Y(4) => npc_mux_out_4_port, Y(3) => 
                           npc_mux_out_3_port, Y(2) => npc_mux_out_2_port, Y(1)
                           => npc_mux_out_1_port, Y(0) => npc_mux_out_0_port);
   NPC_add : NPC_adder port map( inPC(31) => npc_mux_out_31_port, inPC(30) => 
                           npc_mux_out_30_port, inPC(29) => npc_mux_out_29_port
                           , inPC(28) => npc_mux_out_28_port, inPC(27) => 
                           npc_mux_out_27_port, inPC(26) => npc_mux_out_26_port
                           , inPC(25) => npc_mux_out_25_port, inPC(24) => 
                           npc_mux_out_24_port, inPC(23) => npc_mux_out_23_port
                           , inPC(22) => npc_mux_out_22_port, inPC(21) => 
                           npc_mux_out_21_port, inPC(20) => npc_mux_out_20_port
                           , inPC(19) => npc_mux_out_19_port, inPC(18) => 
                           npc_mux_out_18_port, inPC(17) => npc_mux_out_17_port
                           , inPC(16) => npc_mux_out_16_port, inPC(15) => 
                           npc_mux_out_15_port, inPC(14) => npc_mux_out_14_port
                           , inPC(13) => npc_mux_out_13_port, inPC(12) => 
                           npc_mux_out_12_port, inPC(11) => npc_mux_out_11_port
                           , inPC(10) => npc_mux_out_10_port, inPC(9) => 
                           npc_mux_out_9_port, inPC(8) => npc_mux_out_8_port, 
                           inPC(7) => npc_mux_out_7_port, inPC(6) => 
                           npc_mux_out_6_port, inPC(5) => npc_mux_out_5_port, 
                           inPC(4) => npc_mux_out_4_port, inPC(3) => 
                           npc_mux_out_3_port, inPC(2) => npc_mux_out_2_port, 
                           inPC(1) => npc_mux_out_1_port, inPC(0) => 
                           npc_mux_out_0_port, outPC(31) => npc_31_port, 
                           outPC(30) => npc_30_port, outPC(29) => npc_29_port, 
                           outPC(28) => npc_28_port, outPC(27) => npc_27_port, 
                           outPC(26) => npc_26_port, outPC(25) => npc_25_port, 
                           outPC(24) => npc_24_port, outPC(23) => npc_23_port, 
                           outPC(22) => npc_22_port, outPC(21) => npc_21_port, 
                           outPC(20) => npc_20_port, outPC(19) => npc_19_port, 
                           outPC(18) => npc_18_port, outPC(17) => npc_17_port, 
                           outPC(16) => npc_16_port, outPC(15) => npc_15_port, 
                           outPC(14) => npc_14_port, outPC(13) => npc_13_port, 
                           outPC(12) => npc_12_port, outPC(11) => npc_11_port, 
                           outPC(10) => npc_10_port, outPC(9) => npc_9_port, 
                           outPC(8) => npc_8_port, outPC(7) => npc_7_port, 
                           outPC(6) => npc_6_port, outPC(5) => npc_5_port, 
                           outPC(4) => npc_4_port, outPC(3) => npc_3_port, 
                           outPC(2) => npc_2_port, outPC(1) => npc_1_port, 
                           outPC(0) => npc_0_port);
   IF_IDs : IF_ID port map( CLK => Clk, RST => n16, DISCARD => discard_s, 
                           NPC_IN(31) => npc_31_port, NPC_IN(30) => npc_30_port
                           , NPC_IN(29) => npc_29_port, NPC_IN(28) => 
                           npc_28_port, NPC_IN(27) => npc_27_port, NPC_IN(26) 
                           => npc_26_port, NPC_IN(25) => npc_25_port, 
                           NPC_IN(24) => npc_24_port, NPC_IN(23) => npc_23_port
                           , NPC_IN(22) => npc_22_port, NPC_IN(21) => 
                           npc_21_port, NPC_IN(20) => npc_20_port, NPC_IN(19) 
                           => npc_19_port, NPC_IN(18) => npc_18_port, 
                           NPC_IN(17) => npc_17_port, NPC_IN(16) => npc_16_port
                           , NPC_IN(15) => npc_15_port, NPC_IN(14) => 
                           npc_14_port, NPC_IN(13) => npc_13_port, NPC_IN(12) 
                           => npc_12_port, NPC_IN(11) => npc_11_port, 
                           NPC_IN(10) => npc_10_port, NPC_IN(9) => npc_9_port, 
                           NPC_IN(8) => npc_8_port, NPC_IN(7) => npc_7_port, 
                           NPC_IN(6) => npc_6_port, NPC_IN(5) => npc_5_port, 
                           NPC_IN(4) => npc_4_port, NPC_IN(3) => npc_3_port, 
                           NPC_IN(2) => npc_2_port, NPC_IN(1) => npc_1_port, 
                           NPC_IN(0) => npc_0_port, NPC_L_IN(31) => 
                           link_addr_F_31_port, NPC_L_IN(30) => 
                           link_addr_F_30_port, NPC_L_IN(29) => 
                           link_addr_F_29_port, NPC_L_IN(28) => 
                           link_addr_F_28_port, NPC_L_IN(27) => 
                           link_addr_F_27_port, NPC_L_IN(26) => 
                           link_addr_F_26_port, NPC_L_IN(25) => 
                           link_addr_F_25_port, NPC_L_IN(24) => 
                           link_addr_F_24_port, NPC_L_IN(23) => 
                           link_addr_F_23_port, NPC_L_IN(22) => 
                           link_addr_F_22_port, NPC_L_IN(21) => 
                           link_addr_F_21_port, NPC_L_IN(20) => 
                           link_addr_F_20_port, NPC_L_IN(19) => 
                           link_addr_F_19_port, NPC_L_IN(18) => 
                           link_addr_F_18_port, NPC_L_IN(17) => 
                           link_addr_F_17_port, NPC_L_IN(16) => 
                           link_addr_F_16_port, NPC_L_IN(15) => 
                           link_addr_F_15_port, NPC_L_IN(14) => 
                           link_addr_F_14_port, NPC_L_IN(13) => 
                           link_addr_F_13_port, NPC_L_IN(12) => 
                           link_addr_F_12_port, NPC_L_IN(11) => 
                           link_addr_F_11_port, NPC_L_IN(10) => 
                           link_addr_F_10_port, NPC_L_IN(9) => 
                           link_addr_F_9_port, NPC_L_IN(8) => 
                           link_addr_F_8_port, NPC_L_IN(7) => 
                           link_addr_F_7_port, NPC_L_IN(6) => 
                           link_addr_F_6_port, NPC_L_IN(5) => 
                           link_addr_F_5_port, NPC_L_IN(4) => 
                           link_addr_F_4_port, NPC_L_IN(3) => 
                           link_addr_F_3_port, NPC_L_IN(2) => 
                           link_addr_F_2_port, NPC_L_IN(1) => 
                           link_addr_F_1_port, NPC_L_IN(0) => 
                           link_addr_F_0_port, IR_IN(31) => IRAM_OUT(31), 
                           IR_IN(30) => IRAM_OUT(30), IR_IN(29) => IRAM_OUT(29)
                           , IR_IN(28) => IRAM_OUT(28), IR_IN(27) => 
                           IRAM_OUT(27), IR_IN(26) => IRAM_OUT(26), IR_IN(25) 
                           => IRAM_OUT(25), IR_IN(24) => IRAM_OUT(24), 
                           IR_IN(23) => IRAM_OUT(23), IR_IN(22) => IRAM_OUT(22)
                           , IR_IN(21) => IRAM_OUT(21), IR_IN(20) => 
                           IRAM_OUT(20), IR_IN(19) => IRAM_OUT(19), IR_IN(18) 
                           => IRAM_OUT(18), IR_IN(17) => IRAM_OUT(17), 
                           IR_IN(16) => IRAM_OUT(16), IR_IN(15) => IRAM_OUT(15)
                           , IR_IN(14) => IRAM_OUT(14), IR_IN(13) => 
                           IRAM_OUT(13), IR_IN(12) => IRAM_OUT(12), IR_IN(11) 
                           => IRAM_OUT(11), IR_IN(10) => IRAM_OUT(10), IR_IN(9)
                           => IRAM_OUT(9), IR_IN(8) => IRAM_OUT(8), IR_IN(7) =>
                           IRAM_OUT(7), IR_IN(6) => IRAM_OUT(6), IR_IN(5) => 
                           IRAM_OUT(5), IR_IN(4) => IRAM_OUT(4), IR_IN(3) => 
                           IRAM_OUT(3), IR_IN(2) => IRAM_OUT(2), IR_IN(1) => 
                           IRAM_OUT(1), IR_IN(0) => IRAM_OUT(0), PR_IN => 
                           prediction, NPC_OUT(31) => npc_D_31_port, 
                           NPC_OUT(30) => npc_D_30_port, NPC_OUT(29) => 
                           npc_D_29_port, NPC_OUT(28) => npc_D_28_port, 
                           NPC_OUT(27) => npc_D_27_port, NPC_OUT(26) => 
                           npc_D_26_port, NPC_OUT(25) => npc_D_25_port, 
                           NPC_OUT(24) => npc_D_24_port, NPC_OUT(23) => 
                           npc_D_23_port, NPC_OUT(22) => npc_D_22_port, 
                           NPC_OUT(21) => npc_D_21_port, NPC_OUT(20) => 
                           npc_D_20_port, NPC_OUT(19) => npc_D_19_port, 
                           NPC_OUT(18) => npc_D_18_port, NPC_OUT(17) => 
                           npc_D_17_port, NPC_OUT(16) => npc_D_16_port, 
                           NPC_OUT(15) => npc_D_15_port, NPC_OUT(14) => 
                           npc_D_14_port, NPC_OUT(13) => npc_D_13_port, 
                           NPC_OUT(12) => npc_D_12_port, NPC_OUT(11) => 
                           npc_D_11_port, NPC_OUT(10) => npc_D_10_port, 
                           NPC_OUT(9) => npc_D_9_port, NPC_OUT(8) => 
                           npc_D_8_port, NPC_OUT(7) => npc_D_7_port, NPC_OUT(6)
                           => npc_D_6_port, NPC_OUT(5) => npc_D_5_port, 
                           NPC_OUT(4) => npc_D_4_port, NPC_OUT(3) => 
                           npc_D_3_port, NPC_OUT(2) => npc_D_2_port, NPC_OUT(1)
                           => npc_D_1_port, NPC_OUT(0) => npc_D_0_port, 
                           NPC_L_OUT(31) => link_addr_D_31_port, NPC_L_OUT(30) 
                           => link_addr_D_30_port, NPC_L_OUT(29) => 
                           link_addr_D_29_port, NPC_L_OUT(28) => 
                           link_addr_D_28_port, NPC_L_OUT(27) => 
                           link_addr_D_27_port, NPC_L_OUT(26) => 
                           link_addr_D_26_port, NPC_L_OUT(25) => 
                           link_addr_D_25_port, NPC_L_OUT(24) => 
                           link_addr_D_24_port, NPC_L_OUT(23) => 
                           link_addr_D_23_port, NPC_L_OUT(22) => 
                           link_addr_D_22_port, NPC_L_OUT(21) => 
                           link_addr_D_21_port, NPC_L_OUT(20) => 
                           link_addr_D_20_port, NPC_L_OUT(19) => 
                           link_addr_D_19_port, NPC_L_OUT(18) => 
                           link_addr_D_18_port, NPC_L_OUT(17) => 
                           link_addr_D_17_port, NPC_L_OUT(16) => 
                           link_addr_D_16_port, NPC_L_OUT(15) => 
                           link_addr_D_15_port, NPC_L_OUT(14) => 
                           link_addr_D_14_port, NPC_L_OUT(13) => 
                           link_addr_D_13_port, NPC_L_OUT(12) => 
                           link_addr_D_12_port, NPC_L_OUT(11) => 
                           link_addr_D_11_port, NPC_L_OUT(10) => 
                           link_addr_D_10_port, NPC_L_OUT(9) => 
                           link_addr_D_9_port, NPC_L_OUT(8) => 
                           link_addr_D_8_port, NPC_L_OUT(7) => 
                           link_addr_D_7_port, NPC_L_OUT(6) => 
                           link_addr_D_6_port, NPC_L_OUT(5) => 
                           link_addr_D_5_port, NPC_L_OUT(4) => 
                           link_addr_D_4_port, NPC_L_OUT(3) => 
                           link_addr_D_3_port, NPC_L_OUT(2) => 
                           link_addr_D_2_port, NPC_L_OUT(1) => 
                           link_addr_D_1_port, NPC_L_OUT(0) => 
                           link_addr_D_0_port, IR_OUT(31) => IR1_31_port, 
                           IR_OUT(30) => IR1_30_port, IR_OUT(29) => IR1_29_port
                           , IR_OUT(28) => IR1_28_port, IR_OUT(27) => 
                           IR1_27_port, IR_OUT(26) => IR1_26_port, IR_OUT(25) 
                           => IR1_25_port, IR_OUT(24) => IR1_24_port, 
                           IR_OUT(23) => IR1_23_port, IR_OUT(22) => IR1_22_port
                           , IR_OUT(21) => IR1_21_port, IR_OUT(20) => 
                           IR1_20_port, IR_OUT(19) => IR1_19_port, IR_OUT(18) 
                           => IR1_18_port, IR_OUT(17) => IR1_17_port, 
                           IR_OUT(16) => IR1_16_port, IR_OUT(15) => IR1_15_port
                           , IR_OUT(14) => IR1_14_port, IR_OUT(13) => 
                           IR1_13_port, IR_OUT(12) => IR1_12_port, IR_OUT(11) 
                           => IR1_11_port, IR_OUT(10) => IR1_10_port, IR_OUT(9)
                           => IR1_9_port, IR_OUT(8) => IR1_8_port, IR_OUT(7) =>
                           IR1_7_port, IR_OUT(6) => IR1_6_port, IR_OUT(5) => 
                           IR1_5_port, IR_OUT(4) => IR1_4_port, IR_OUT(3) => 
                           IR1_3_port, IR_OUT(2) => IR1_2_port, IR_OUT(1) => 
                           IR1_1_port, IR_OUT(0) => IR1_0_port, PR_OUT => pr_D)
                           ;
   dec : IR_decoder port map( rst => n16, IR_OUT(20) => IR1_31_port, IR_OUT(19)
                           => IR1_30_port, IR_OUT(18) => IR1_29_port, 
                           IR_OUT(17) => IR1_28_port, IR_OUT(16) => IR1_27_port
                           , IR_OUT(15) => IR1_26_port, IR_OUT(14) => 
                           IR1_25_port, IR_OUT(13) => IR1_24_port, IR_OUT(12) 
                           => IR1_23_port, IR_OUT(11) => IR1_22_port, 
                           IR_OUT(10) => IR1_21_port, IR_OUT(9) => IR1_20_port,
                           IR_OUT(8) => IR1_19_port, IR_OUT(7) => IR1_18_port, 
                           IR_OUT(6) => IR1_17_port, IR_OUT(5) => IR1_16_port, 
                           IR_OUT(4) => IR1_15_port, IR_OUT(3) => IR1_14_port, 
                           IR_OUT(2) => IR1_13_port, IR_OUT(1) => IR1_12_port, 
                           IR_OUT(0) => IR1_11_port, ADDS1(4) => add_S1_4_port,
                           ADDS1(3) => add_S1_3_port, ADDS1(2) => add_S1_2_port
                           , ADDS1(1) => add_S1_1_port, ADDS1(0) => 
                           add_S1_0_port, ADDS2(4) => add_S2_4_port, ADDS2(3) 
                           => add_S2_3_port, ADDS2(2) => add_S2_2_port, 
                           ADDS2(1) => add_S2_1_port, ADDS2(0) => add_S2_0_port
                           , ADDD(4) => dest_D_4_port, ADDD(3) => dest_D_3_port
                           , ADDD(2) => dest_D_2_port, ADDD(1) => dest_D_1_port
                           , ADDD(0) => dest_D_0_port);
   Reg_F : register_file_N32_addBit5 port map( RESET => n16, RE => 
                           X_Logic1_port, WE => RF_WE, ADD_WR(4) => 
                           add_D_4_port, ADD_WR(3) => add_D_3_port, ADD_WR(2) 
                           => add_D_2_port, ADD_WR(1) => add_D_1_port, 
                           ADD_WR(0) => add_D_0_port, ADD_RDA(4) => 
                           add_S1_4_port, ADD_RDA(3) => add_S1_3_port, 
                           ADD_RDA(2) => add_S1_2_port, ADD_RDA(1) => 
                           add_S1_1_port, ADD_RDA(0) => add_S1_0_port, 
                           ADD_RDB(4) => add_S2_4_port, ADD_RDB(3) => 
                           add_S2_3_port, ADD_RDB(2) => add_S2_2_port, 
                           ADD_RDB(1) => add_S2_1_port, ADD_RDB(0) => 
                           add_S2_0_port, DATAIN(31) => WB_31_port, DATAIN(30) 
                           => WB_30_port, DATAIN(29) => WB_29_port, DATAIN(28) 
                           => WB_28_port, DATAIN(27) => WB_27_port, DATAIN(26) 
                           => WB_26_port, DATAIN(25) => WB_25_port, DATAIN(24) 
                           => WB_24_port, DATAIN(23) => WB_23_port, DATAIN(22) 
                           => WB_22_port, DATAIN(21) => WB_21_port, DATAIN(20) 
                           => WB_20_port, DATAIN(19) => WB_19_port, DATAIN(18) 
                           => WB_18_port, DATAIN(17) => WB_17_port, DATAIN(16) 
                           => WB_16_port, DATAIN(15) => WB_15_port, DATAIN(14) 
                           => WB_14_port, DATAIN(13) => WB_13_port, DATAIN(12) 
                           => WB_12_port, DATAIN(11) => WB_11_port, DATAIN(10) 
                           => WB_10_port, DATAIN(9) => WB_9_port, DATAIN(8) => 
                           WB_8_port, DATAIN(7) => WB_7_port, DATAIN(6) => 
                           WB_6_port, DATAIN(5) => WB_5_port, DATAIN(4) => 
                           WB_4_port, DATAIN(3) => WB_3_port, DATAIN(2) => 
                           WB_2_port, DATAIN(1) => WB_1_port, DATAIN(0) => 
                           WB_0_port, OUTA(31) => a_out_31_port, OUTA(30) => 
                           a_out_30_port, OUTA(29) => a_out_29_port, OUTA(28) 
                           => a_out_28_port, OUTA(27) => a_out_27_port, 
                           OUTA(26) => a_out_26_port, OUTA(25) => a_out_25_port
                           , OUTA(24) => a_out_24_port, OUTA(23) => 
                           a_out_23_port, OUTA(22) => a_out_22_port, OUTA(21) 
                           => a_out_21_port, OUTA(20) => a_out_20_port, 
                           OUTA(19) => a_out_19_port, OUTA(18) => a_out_18_port
                           , OUTA(17) => a_out_17_port, OUTA(16) => 
                           a_out_16_port, OUTA(15) => a_out_15_port, OUTA(14) 
                           => a_out_14_port, OUTA(13) => a_out_13_port, 
                           OUTA(12) => a_out_12_port, OUTA(11) => a_out_11_port
                           , OUTA(10) => a_out_10_port, OUTA(9) => a_out_9_port
                           , OUTA(8) => a_out_8_port, OUTA(7) => a_out_7_port, 
                           OUTA(6) => a_out_6_port, OUTA(5) => a_out_5_port, 
                           OUTA(4) => a_out_4_port, OUTA(3) => a_out_3_port, 
                           OUTA(2) => a_out_2_port, OUTA(1) => a_out_1_port, 
                           OUTA(0) => a_out_0_port, OUTB(31) => b_out_31_port, 
                           OUTB(30) => b_out_30_port, OUTB(29) => b_out_29_port
                           , OUTB(28) => b_out_28_port, OUTB(27) => 
                           b_out_27_port, OUTB(26) => b_out_26_port, OUTB(25) 
                           => b_out_25_port, OUTB(24) => b_out_24_port, 
                           OUTB(23) => b_out_23_port, OUTB(22) => b_out_22_port
                           , OUTB(21) => b_out_21_port, OUTB(20) => 
                           b_out_20_port, OUTB(19) => b_out_19_port, OUTB(18) 
                           => b_out_18_port, OUTB(17) => b_out_17_port, 
                           OUTB(16) => b_out_16_port, OUTB(15) => b_out_15_port
                           , OUTB(14) => b_out_14_port, OUTB(13) => 
                           b_out_13_port, OUTB(12) => b_out_12_port, OUTB(11) 
                           => b_out_11_port, OUTB(10) => b_out_10_port, OUTB(9)
                           => b_out_9_port, OUTB(8) => b_out_8_port, OUTB(7) =>
                           b_out_7_port, OUTB(6) => b_out_6_port, OUTB(5) => 
                           b_out_5_port, OUTB(4) => b_out_4_port, OUTB(3) => 
                           b_out_3_port, OUTB(2) => b_out_2_port, OUTB(1) => 
                           b_out_1_port, OUTB(0) => b_out_0_port);
   sign_ext : sign_extender port map( d_in(31) => IR1_31_port, d_in(30) => 
                           IR1_30_port, d_in(29) => IR1_29_port, d_in(28) => 
                           IR1_28_port, d_in(27) => IR1_27_port, d_in(26) => 
                           IR1_26_port, d_in(25) => IR1_25_port, d_in(24) => 
                           IR1_24_port, d_in(23) => IR1_23_port, d_in(22) => 
                           IR1_22_port, d_in(21) => IR1_21_port, d_in(20) => 
                           IR1_20_port, d_in(19) => IR1_19_port, d_in(18) => 
                           IR1_18_port, d_in(17) => IR1_17_port, d_in(16) => 
                           IR1_16_port, d_in(15) => IR1_15_port, d_in(14) => 
                           IR1_14_port, d_in(13) => IR1_13_port, d_in(12) => 
                           IR1_12_port, d_in(11) => IR1_11_port, d_in(10) => 
                           IR1_10_port, d_in(9) => IR1_9_port, d_in(8) => 
                           IR1_8_port, d_in(7) => IR1_7_port, d_in(6) => 
                           IR1_6_port, d_in(5) => IR1_5_port, d_in(4) => 
                           IR1_4_port, d_in(3) => IR1_3_port, d_in(2) => 
                           IR1_2_port, d_in(1) => IR1_1_port, d_in(0) => 
                           IR1_0_port, rst => n16, d_ext(31) => imm_out_31_port
                           , d_ext(30) => imm_out_30_port, d_ext(29) => 
                           imm_out_29_port, d_ext(28) => imm_out_28_port, 
                           d_ext(27) => imm_out_27_port, d_ext(26) => 
                           imm_out_26_port, d_ext(25) => imm_out_25_port, 
                           d_ext(24) => imm_out_24_port, d_ext(23) => 
                           imm_out_23_port, d_ext(22) => imm_out_22_port, 
                           d_ext(21) => imm_out_21_port, d_ext(20) => 
                           imm_out_20_port, d_ext(19) => imm_out_19_port, 
                           d_ext(18) => imm_out_18_port, d_ext(17) => 
                           imm_out_17_port, d_ext(16) => imm_out_16_port, 
                           d_ext(15) => imm_out_15_port, d_ext(14) => 
                           imm_out_14_port, d_ext(13) => imm_out_13_port, 
                           d_ext(12) => imm_out_12_port, d_ext(11) => 
                           imm_out_11_port, d_ext(10) => imm_out_10_port, 
                           d_ext(9) => imm_out_9_port, d_ext(8) => 
                           imm_out_8_port, d_ext(7) => imm_out_7_port, d_ext(6)
                           => imm_out_6_port, d_ext(5) => imm_out_5_port, 
                           d_ext(4) => imm_out_4_port, d_ext(3) => 
                           imm_out_3_port, d_ext(2) => imm_out_2_port, d_ext(1)
                           => imm_out_1_port, d_ext(0) => imm_out_0_port);
   ID_EXs : ID_EX port map( CLK => Clk, RST => n16, NPC_IN(31) => npc_D_31_port
                           , NPC_IN(30) => npc_D_30_port, NPC_IN(29) => 
                           npc_D_29_port, NPC_IN(28) => npc_D_28_port, 
                           NPC_IN(27) => npc_D_27_port, NPC_IN(26) => 
                           npc_D_26_port, NPC_IN(25) => npc_D_25_port, 
                           NPC_IN(24) => npc_D_24_port, NPC_IN(23) => 
                           npc_D_23_port, NPC_IN(22) => npc_D_22_port, 
                           NPC_IN(21) => npc_D_21_port, NPC_IN(20) => 
                           npc_D_20_port, NPC_IN(19) => npc_D_19_port, 
                           NPC_IN(18) => npc_D_18_port, NPC_IN(17) => 
                           npc_D_17_port, NPC_IN(16) => npc_D_16_port, 
                           NPC_IN(15) => npc_D_15_port, NPC_IN(14) => 
                           npc_D_14_port, NPC_IN(13) => npc_D_13_port, 
                           NPC_IN(12) => npc_D_12_port, NPC_IN(11) => 
                           npc_D_11_port, NPC_IN(10) => npc_D_10_port, 
                           NPC_IN(9) => npc_D_9_port, NPC_IN(8) => npc_D_8_port
                           , NPC_IN(7) => npc_D_7_port, NPC_IN(6) => 
                           npc_D_6_port, NPC_IN(5) => npc_D_5_port, NPC_IN(4) 
                           => npc_D_4_port, NPC_IN(3) => npc_D_3_port, 
                           NPC_IN(2) => npc_D_2_port, NPC_IN(1) => npc_D_1_port
                           , NPC_IN(0) => npc_D_0_port, NPC_L_IN(31) => 
                           link_addr_D_31_port, NPC_L_IN(30) => 
                           link_addr_D_30_port, NPC_L_IN(29) => 
                           link_addr_D_29_port, NPC_L_IN(28) => 
                           link_addr_D_28_port, NPC_L_IN(27) => 
                           link_addr_D_27_port, NPC_L_IN(26) => 
                           link_addr_D_26_port, NPC_L_IN(25) => 
                           link_addr_D_25_port, NPC_L_IN(24) => 
                           link_addr_D_24_port, NPC_L_IN(23) => 
                           link_addr_D_23_port, NPC_L_IN(22) => 
                           link_addr_D_22_port, NPC_L_IN(21) => 
                           link_addr_D_21_port, NPC_L_IN(20) => 
                           link_addr_D_20_port, NPC_L_IN(19) => 
                           link_addr_D_19_port, NPC_L_IN(18) => 
                           link_addr_D_18_port, NPC_L_IN(17) => 
                           link_addr_D_17_port, NPC_L_IN(16) => 
                           link_addr_D_16_port, NPC_L_IN(15) => 
                           link_addr_D_15_port, NPC_L_IN(14) => 
                           link_addr_D_14_port, NPC_L_IN(13) => 
                           link_addr_D_13_port, NPC_L_IN(12) => 
                           link_addr_D_12_port, NPC_L_IN(11) => 
                           link_addr_D_11_port, NPC_L_IN(10) => 
                           link_addr_D_10_port, NPC_L_IN(9) => 
                           link_addr_D_9_port, NPC_L_IN(8) => 
                           link_addr_D_8_port, NPC_L_IN(7) => 
                           link_addr_D_7_port, NPC_L_IN(6) => 
                           link_addr_D_6_port, NPC_L_IN(5) => 
                           link_addr_D_5_port, NPC_L_IN(4) => 
                           link_addr_D_4_port, NPC_L_IN(3) => 
                           link_addr_D_3_port, NPC_L_IN(2) => 
                           link_addr_D_2_port, NPC_L_IN(1) => 
                           link_addr_D_1_port, NPC_L_IN(0) => 
                           link_addr_D_0_port, A_IN(31) => a_out_31_port, 
                           A_IN(30) => a_out_30_port, A_IN(29) => a_out_29_port
                           , A_IN(28) => a_out_28_port, A_IN(27) => 
                           a_out_27_port, A_IN(26) => a_out_26_port, A_IN(25) 
                           => a_out_25_port, A_IN(24) => a_out_24_port, 
                           A_IN(23) => a_out_23_port, A_IN(22) => a_out_22_port
                           , A_IN(21) => a_out_21_port, A_IN(20) => 
                           a_out_20_port, A_IN(19) => a_out_19_port, A_IN(18) 
                           => a_out_18_port, A_IN(17) => a_out_17_port, 
                           A_IN(16) => a_out_16_port, A_IN(15) => a_out_15_port
                           , A_IN(14) => a_out_14_port, A_IN(13) => 
                           a_out_13_port, A_IN(12) => a_out_12_port, A_IN(11) 
                           => a_out_11_port, A_IN(10) => a_out_10_port, A_IN(9)
                           => a_out_9_port, A_IN(8) => a_out_8_port, A_IN(7) =>
                           a_out_7_port, A_IN(6) => a_out_6_port, A_IN(5) => 
                           a_out_5_port, A_IN(4) => a_out_4_port, A_IN(3) => 
                           a_out_3_port, A_IN(2) => a_out_2_port, A_IN(1) => 
                           a_out_1_port, A_IN(0) => a_out_0_port, B_IN(31) => 
                           b_out_31_port, B_IN(30) => b_out_30_port, B_IN(29) 
                           => b_out_29_port, B_IN(28) => b_out_28_port, 
                           B_IN(27) => b_out_27_port, B_IN(26) => b_out_26_port
                           , B_IN(25) => b_out_25_port, B_IN(24) => 
                           b_out_24_port, B_IN(23) => b_out_23_port, B_IN(22) 
                           => b_out_22_port, B_IN(21) => b_out_21_port, 
                           B_IN(20) => b_out_20_port, B_IN(19) => b_out_19_port
                           , B_IN(18) => b_out_18_port, B_IN(17) => 
                           b_out_17_port, B_IN(16) => b_out_16_port, B_IN(15) 
                           => b_out_15_port, B_IN(14) => b_out_14_port, 
                           B_IN(13) => b_out_13_port, B_IN(12) => b_out_12_port
                           , B_IN(11) => b_out_11_port, B_IN(10) => 
                           b_out_10_port, B_IN(9) => b_out_9_port, B_IN(8) => 
                           b_out_8_port, B_IN(7) => b_out_7_port, B_IN(6) => 
                           b_out_6_port, B_IN(5) => b_out_5_port, B_IN(4) => 
                           b_out_4_port, B_IN(3) => b_out_3_port, B_IN(2) => 
                           b_out_2_port, B_IN(1) => b_out_1_port, B_IN(0) => 
                           b_out_0_port, IMM_IN(31) => imm_out_31_port, 
                           IMM_IN(30) => imm_out_30_port, IMM_IN(29) => 
                           imm_out_29_port, IMM_IN(28) => imm_out_28_port, 
                           IMM_IN(27) => imm_out_27_port, IMM_IN(26) => 
                           imm_out_26_port, IMM_IN(25) => imm_out_25_port, 
                           IMM_IN(24) => imm_out_24_port, IMM_IN(23) => 
                           imm_out_23_port, IMM_IN(22) => imm_out_22_port, 
                           IMM_IN(21) => imm_out_21_port, IMM_IN(20) => 
                           imm_out_20_port, IMM_IN(19) => imm_out_19_port, 
                           IMM_IN(18) => imm_out_18_port, IMM_IN(17) => 
                           imm_out_17_port, IMM_IN(16) => imm_out_16_port, 
                           IMM_IN(15) => imm_out_15_port, IMM_IN(14) => 
                           imm_out_14_port, IMM_IN(13) => imm_out_13_port, 
                           IMM_IN(12) => imm_out_12_port, IMM_IN(11) => 
                           imm_out_11_port, IMM_IN(10) => imm_out_10_port, 
                           IMM_IN(9) => imm_out_9_port, IMM_IN(8) => 
                           imm_out_8_port, IMM_IN(7) => imm_out_7_port, 
                           IMM_IN(6) => imm_out_6_port, IMM_IN(5) => 
                           imm_out_5_port, IMM_IN(4) => imm_out_4_port, 
                           IMM_IN(3) => imm_out_3_port, IMM_IN(2) => 
                           imm_out_2_port, IMM_IN(1) => imm_out_1_port, 
                           IMM_IN(0) => imm_out_0_port, RS1_IN(4) => 
                           add_S1_4_port, RS1_IN(3) => add_S1_3_port, RS1_IN(2)
                           => add_S1_2_port, RS1_IN(1) => add_S1_1_port, 
                           RS1_IN(0) => add_S1_0_port, RS2_IN(4) => 
                           add_S2_4_port, RS2_IN(3) => add_S2_3_port, RS2_IN(2)
                           => add_S2_2_port, RS2_IN(1) => add_S2_1_port, 
                           RS2_IN(0) => add_S2_0_port, RD_IN(4) => 
                           dest_D_4_port, RD_IN(3) => dest_D_3_port, RD_IN(2) 
                           => dest_D_2_port, RD_IN(1) => dest_D_1_port, 
                           RD_IN(0) => dest_D_0_port, OPCODE_IN(5) => 
                           IR1_31_port, OPCODE_IN(4) => IR1_30_port, 
                           OPCODE_IN(3) => IR1_29_port, OPCODE_IN(2) => 
                           IR1_28_port, OPCODE_IN(1) => IR1_27_port, 
                           OPCODE_IN(0) => IR1_26_port, IR_IN(15) => 
                           IR1_15_port, IR_IN(14) => IR1_14_port, IR_IN(13) => 
                           IR1_13_port, IR_IN(12) => IR1_12_port, IR_IN(11) => 
                           IR1_11_port, IR_IN(10) => IR1_10_port, IR_IN(9) => 
                           IR1_9_port, IR_IN(8) => IR1_8_port, IR_IN(7) => 
                           IR1_7_port, IR_IN(6) => IR1_6_port, IR_IN(5) => 
                           IR1_5_port, IR_IN(4) => IR1_4_port, IR_IN(3) => 
                           IR1_3_port, IR_IN(2) => IR1_2_port, IR_IN(1) => 
                           IR1_1_port, IR_IN(0) => IR1_0_port, PR_IN => pr_D, 
                           NPC_OUT(31) => npc_E_31_port, NPC_OUT(30) => 
                           npc_E_30_port, NPC_OUT(29) => npc_E_29_port, 
                           NPC_OUT(28) => npc_E_28_port, NPC_OUT(27) => 
                           npc_E_27_port, NPC_OUT(26) => npc_E_26_port, 
                           NPC_OUT(25) => npc_E_25_port, NPC_OUT(24) => 
                           npc_E_24_port, NPC_OUT(23) => npc_E_23_port, 
                           NPC_OUT(22) => npc_E_22_port, NPC_OUT(21) => 
                           npc_E_21_port, NPC_OUT(20) => npc_E_20_port, 
                           NPC_OUT(19) => npc_E_19_port, NPC_OUT(18) => 
                           npc_E_18_port, NPC_OUT(17) => npc_E_17_port, 
                           NPC_OUT(16) => npc_E_16_port, NPC_OUT(15) => 
                           npc_E_15_port, NPC_OUT(14) => npc_E_14_port, 
                           NPC_OUT(13) => npc_E_13_port, NPC_OUT(12) => 
                           npc_E_12_port, NPC_OUT(11) => npc_E_11_port, 
                           NPC_OUT(10) => npc_E_10_port, NPC_OUT(9) => 
                           npc_E_9_port, NPC_OUT(8) => npc_E_8_port, NPC_OUT(7)
                           => npc_E_7_port, NPC_OUT(6) => npc_E_6_port, 
                           NPC_OUT(5) => npc_E_5_port, NPC_OUT(4) => 
                           npc_E_4_port, NPC_OUT(3) => npc_E_3_port, NPC_OUT(2)
                           => npc_E_2_port, NPC_OUT(1) => npc_E_1_port, 
                           NPC_OUT(0) => npc_E_0_port, NPC_L_OUT(31) => 
                           link_addr_E_31_port, NPC_L_OUT(30) => 
                           link_addr_E_30_port, NPC_L_OUT(29) => 
                           link_addr_E_29_port, NPC_L_OUT(28) => 
                           link_addr_E_28_port, NPC_L_OUT(27) => 
                           link_addr_E_27_port, NPC_L_OUT(26) => 
                           link_addr_E_26_port, NPC_L_OUT(25) => 
                           link_addr_E_25_port, NPC_L_OUT(24) => 
                           link_addr_E_24_port, NPC_L_OUT(23) => 
                           link_addr_E_23_port, NPC_L_OUT(22) => 
                           link_addr_E_22_port, NPC_L_OUT(21) => 
                           link_addr_E_21_port, NPC_L_OUT(20) => 
                           link_addr_E_20_port, NPC_L_OUT(19) => 
                           link_addr_E_19_port, NPC_L_OUT(18) => 
                           link_addr_E_18_port, NPC_L_OUT(17) => 
                           link_addr_E_17_port, NPC_L_OUT(16) => 
                           link_addr_E_16_port, NPC_L_OUT(15) => 
                           link_addr_E_15_port, NPC_L_OUT(14) => 
                           link_addr_E_14_port, NPC_L_OUT(13) => 
                           link_addr_E_13_port, NPC_L_OUT(12) => 
                           link_addr_E_12_port, NPC_L_OUT(11) => 
                           link_addr_E_11_port, NPC_L_OUT(10) => 
                           link_addr_E_10_port, NPC_L_OUT(9) => 
                           link_addr_E_9_port, NPC_L_OUT(8) => 
                           link_addr_E_8_port, NPC_L_OUT(7) => 
                           link_addr_E_7_port, NPC_L_OUT(6) => 
                           link_addr_E_6_port, NPC_L_OUT(5) => 
                           link_addr_E_5_port, NPC_L_OUT(4) => 
                           link_addr_E_4_port, NPC_L_OUT(3) => 
                           link_addr_E_3_port, NPC_L_OUT(2) => 
                           link_addr_E_2_port, NPC_L_OUT(1) => 
                           link_addr_E_1_port, NPC_L_OUT(0) => 
                           link_addr_E_0_port, A_OUT(31) => A_s_31_port, 
                           A_OUT(30) => A_s_30_port, A_OUT(29) => A_s_29_port, 
                           A_OUT(28) => A_s_28_port, A_OUT(27) => A_s_27_port, 
                           A_OUT(26) => A_s_26_port, A_OUT(25) => A_s_25_port, 
                           A_OUT(24) => A_s_24_port, A_OUT(23) => A_s_23_port, 
                           A_OUT(22) => A_s_22_port, A_OUT(21) => A_s_21_port, 
                           A_OUT(20) => A_s_20_port, A_OUT(19) => A_s_19_port, 
                           A_OUT(18) => A_s_18_port, A_OUT(17) => A_s_17_port, 
                           A_OUT(16) => A_s_16_port, A_OUT(15) => A_s_15_port, 
                           A_OUT(14) => A_s_14_port, A_OUT(13) => A_s_13_port, 
                           A_OUT(12) => A_s_12_port, A_OUT(11) => A_s_11_port, 
                           A_OUT(10) => A_s_10_port, A_OUT(9) => A_s_9_port, 
                           A_OUT(8) => A_s_8_port, A_OUT(7) => A_s_7_port, 
                           A_OUT(6) => A_s_6_port, A_OUT(5) => A_s_5_port, 
                           A_OUT(4) => A_s_4_port, A_OUT(3) => A_s_3_port, 
                           A_OUT(2) => A_s_2_port, A_OUT(1) => A_s_1_port, 
                           A_OUT(0) => A_s_0_port, B_OUT(31) => B_s_31_port, 
                           B_OUT(30) => B_s_30_port, B_OUT(29) => B_s_29_port, 
                           B_OUT(28) => B_s_28_port, B_OUT(27) => B_s_27_port, 
                           B_OUT(26) => B_s_26_port, B_OUT(25) => B_s_25_port, 
                           B_OUT(24) => B_s_24_port, B_OUT(23) => B_s_23_port, 
                           B_OUT(22) => B_s_22_port, B_OUT(21) => B_s_21_port, 
                           B_OUT(20) => B_s_20_port, B_OUT(19) => B_s_19_port, 
                           B_OUT(18) => B_s_18_port, B_OUT(17) => B_s_17_port, 
                           B_OUT(16) => B_s_16_port, B_OUT(15) => B_s_15_port, 
                           B_OUT(14) => B_s_14_port, B_OUT(13) => B_s_13_port, 
                           B_OUT(12) => B_s_12_port, B_OUT(11) => B_s_11_port, 
                           B_OUT(10) => B_s_10_port, B_OUT(9) => B_s_9_port, 
                           B_OUT(8) => B_s_8_port, B_OUT(7) => B_s_7_port, 
                           B_OUT(6) => B_s_6_port, B_OUT(5) => B_s_5_port, 
                           B_OUT(4) => B_s_4_port, B_OUT(3) => B_s_3_port, 
                           B_OUT(2) => B_s_2_port, B_OUT(1) => B_s_1_port, 
                           B_OUT(0) => B_s_0_port, IMM_OUT(31) => IMM_s_31_port
                           , IMM_OUT(30) => IMM_s_30_port, IMM_OUT(29) => 
                           IMM_s_29_port, IMM_OUT(28) => IMM_s_28_port, 
                           IMM_OUT(27) => IMM_s_27_port, IMM_OUT(26) => 
                           IMM_s_26_port, IMM_OUT(25) => IMM_s_25_port, 
                           IMM_OUT(24) => IMM_s_24_port, IMM_OUT(23) => 
                           IMM_s_23_port, IMM_OUT(22) => IMM_s_22_port, 
                           IMM_OUT(21) => IMM_s_21_port, IMM_OUT(20) => 
                           IMM_s_20_port, IMM_OUT(19) => IMM_s_19_port, 
                           IMM_OUT(18) => IMM_s_18_port, IMM_OUT(17) => 
                           IMM_s_17_port, IMM_OUT(16) => IMM_s_16_port, 
                           IMM_OUT(15) => IMM_s_15_port, IMM_OUT(14) => 
                           IMM_s_14_port, IMM_OUT(13) => IMM_s_13_port, 
                           IMM_OUT(12) => IMM_s_12_port, IMM_OUT(11) => 
                           IMM_s_11_port, IMM_OUT(10) => IMM_s_10_port, 
                           IMM_OUT(9) => IMM_s_9_port, IMM_OUT(8) => 
                           IMM_s_8_port, IMM_OUT(7) => IMM_s_7_port, IMM_OUT(6)
                           => IMM_s_6_port, IMM_OUT(5) => IMM_s_5_port, 
                           IMM_OUT(4) => IMM_s_4_port, IMM_OUT(3) => 
                           IMM_s_3_port, IMM_OUT(2) => IMM_s_2_port, IMM_OUT(1)
                           => IMM_s_1_port, IMM_OUT(0) => IMM_s_0_port, 
                           RS1_OUT(4) => Rs1_4_port, RS1_OUT(3) => Rs1_3_port, 
                           RS1_OUT(2) => Rs1_2_port, RS1_OUT(1) => Rs1_1_port, 
                           RS1_OUT(0) => Rs1_0_port, RS2_OUT(4) => Rs2_4_port, 
                           RS2_OUT(3) => Rs2_3_port, RS2_OUT(2) => Rs2_2_port, 
                           RS2_OUT(1) => Rs2_1_port, RS2_OUT(0) => Rs2_0_port, 
                           RD_OUT(4) => dest_E_4_port, RD_OUT(3) => 
                           dest_E_3_port, RD_OUT(2) => dest_E_2_port, RD_OUT(1)
                           => dest_E_1_port, RD_OUT(0) => dest_E_0_port, 
                           OPCODE_OUT(5) => opcode_E_5_port, OPCODE_OUT(4) => 
                           opcode_E_4_port, OPCODE_OUT(3) => opcode_E_3_port, 
                           OPCODE_OUT(2) => opcode_E_2_port, OPCODE_OUT(1) => 
                           opcode_E_1_port, OPCODE_OUT(0) => opcode_E_0_port, 
                           IR_OUT(15) => ir_E_15_port, IR_OUT(14) => 
                           ir_E_14_port, IR_OUT(13) => ir_E_13_port, IR_OUT(12)
                           => ir_E_12_port, IR_OUT(11) => ir_E_11_port, 
                           IR_OUT(10) => ir_E_10_port, IR_OUT(9) => ir_E_9_port
                           , IR_OUT(8) => ir_E_8_port, IR_OUT(7) => ir_E_7_port
                           , IR_OUT(6) => ir_E_6_port, IR_OUT(5) => ir_E_5_port
                           , IR_OUT(4) => ir_E_4_port, IR_OUT(3) => ir_E_3_port
                           , IR_OUT(2) => ir_E_2_port, IR_OUT(1) => ir_E_1_port
                           , IR_OUT(0) => ir_E_0_port, PR_OUT => pr_E);
   A_mux : MUX21_GENERIC_N32_2 port map( A(31) => npc_E_31_port, A(30) => 
                           npc_E_30_port, A(29) => npc_E_29_port, A(28) => 
                           npc_E_28_port, A(27) => npc_E_27_port, A(26) => 
                           npc_E_26_port, A(25) => npc_E_25_port, A(24) => 
                           npc_E_24_port, A(23) => npc_E_23_port, A(22) => 
                           npc_E_22_port, A(21) => npc_E_21_port, A(20) => 
                           npc_E_20_port, A(19) => npc_E_19_port, A(18) => 
                           npc_E_18_port, A(17) => npc_E_17_port, A(16) => 
                           npc_E_16_port, A(15) => npc_E_15_port, A(14) => 
                           npc_E_14_port, A(13) => npc_E_13_port, A(12) => 
                           npc_E_12_port, A(11) => npc_E_11_port, A(10) => 
                           npc_E_10_port, A(9) => npc_E_9_port, A(8) => 
                           npc_E_8_port, A(7) => npc_E_7_port, A(6) => 
                           npc_E_6_port, A(5) => npc_E_5_port, A(4) => 
                           npc_E_4_port, A(3) => npc_E_3_port, A(2) => 
                           npc_E_2_port, A(1) => npc_E_1_port, A(0) => 
                           npc_E_0_port, B(31) => A_s_31_port, B(30) => 
                           A_s_30_port, B(29) => A_s_29_port, B(28) => 
                           A_s_28_port, B(27) => A_s_27_port, B(26) => 
                           A_s_26_port, B(25) => A_s_25_port, B(24) => 
                           A_s_24_port, B(23) => A_s_23_port, B(22) => 
                           A_s_22_port, B(21) => A_s_21_port, B(20) => 
                           A_s_20_port, B(19) => A_s_19_port, B(18) => 
                           A_s_18_port, B(17) => A_s_17_port, B(16) => 
                           A_s_16_port, B(15) => A_s_15_port, B(14) => 
                           A_s_14_port, B(13) => A_s_13_port, B(12) => 
                           A_s_12_port, B(11) => A_s_11_port, B(10) => 
                           A_s_10_port, B(9) => A_s_9_port, B(8) => A_s_8_port,
                           B(7) => A_s_7_port, B(6) => A_s_6_port, B(5) => 
                           A_s_5_port, B(4) => A_s_4_port, B(3) => A_s_3_port, 
                           B(2) => A_s_2_port, B(1) => A_s_1_port, B(0) => 
                           A_s_0_port, SEL => MUXA_SEL, Y(31) => 
                           mux_a_in_31_port, Y(30) => mux_a_in_30_port, Y(29) 
                           => mux_a_in_29_port, Y(28) => mux_a_in_28_port, 
                           Y(27) => mux_a_in_27_port, Y(26) => mux_a_in_26_port
                           , Y(25) => mux_a_in_25_port, Y(24) => 
                           mux_a_in_24_port, Y(23) => mux_a_in_23_port, Y(22) 
                           => mux_a_in_22_port, Y(21) => mux_a_in_21_port, 
                           Y(20) => mux_a_in_20_port, Y(19) => mux_a_in_19_port
                           , Y(18) => mux_a_in_18_port, Y(17) => 
                           mux_a_in_17_port, Y(16) => mux_a_in_16_port, Y(15) 
                           => mux_a_in_15_port, Y(14) => mux_a_in_14_port, 
                           Y(13) => mux_a_in_13_port, Y(12) => mux_a_in_12_port
                           , Y(11) => mux_a_in_11_port, Y(10) => 
                           mux_a_in_10_port, Y(9) => mux_a_in_9_port, Y(8) => 
                           mux_a_in_8_port, Y(7) => mux_a_in_7_port, Y(6) => 
                           mux_a_in_6_port, Y(5) => mux_a_in_5_port, Y(4) => 
                           mux_a_in_4_port, Y(3) => mux_a_in_3_port, Y(2) => 
                           mux_a_in_2_port, Y(1) => mux_a_in_1_port, Y(0) => 
                           mux_a_in_0_port);
   B_mux : MUX21_GENERIC_N32_1 port map( A(31) => IMM_s_31_port, A(30) => 
                           IMM_s_30_port, A(29) => IMM_s_29_port, A(28) => 
                           IMM_s_28_port, A(27) => IMM_s_27_port, A(26) => 
                           IMM_s_26_port, A(25) => IMM_s_25_port, A(24) => 
                           IMM_s_24_port, A(23) => IMM_s_23_port, A(22) => 
                           IMM_s_22_port, A(21) => IMM_s_21_port, A(20) => 
                           IMM_s_20_port, A(19) => IMM_s_19_port, A(18) => 
                           IMM_s_18_port, A(17) => IMM_s_17_port, A(16) => 
                           IMM_s_16_port, A(15) => IMM_s_15_port, A(14) => 
                           IMM_s_14_port, A(13) => IMM_s_13_port, A(12) => 
                           IMM_s_12_port, A(11) => IMM_s_11_port, A(10) => 
                           IMM_s_10_port, A(9) => IMM_s_9_port, A(8) => 
                           IMM_s_8_port, A(7) => IMM_s_7_port, A(6) => 
                           IMM_s_6_port, A(5) => IMM_s_5_port, A(4) => 
                           IMM_s_4_port, A(3) => IMM_s_3_port, A(2) => 
                           IMM_s_2_port, A(1) => IMM_s_1_port, A(0) => 
                           IMM_s_0_port, B(31) => B_s_31_port, B(30) => 
                           B_s_30_port, B(29) => B_s_29_port, B(28) => 
                           B_s_28_port, B(27) => B_s_27_port, B(26) => 
                           B_s_26_port, B(25) => B_s_25_port, B(24) => 
                           B_s_24_port, B(23) => B_s_23_port, B(22) => 
                           B_s_22_port, B(21) => B_s_21_port, B(20) => 
                           B_s_20_port, B(19) => B_s_19_port, B(18) => 
                           B_s_18_port, B(17) => B_s_17_port, B(16) => 
                           B_s_16_port, B(15) => B_s_15_port, B(14) => 
                           B_s_14_port, B(13) => B_s_13_port, B(12) => 
                           B_s_12_port, B(11) => B_s_11_port, B(10) => 
                           B_s_10_port, B(9) => B_s_9_port, B(8) => B_s_8_port,
                           B(7) => B_s_7_port, B(6) => B_s_6_port, B(5) => 
                           B_s_5_port, B(4) => B_s_4_port, B(3) => B_s_3_port, 
                           B(2) => B_s_2_port, B(1) => B_s_1_port, B(0) => 
                           B_s_0_port, SEL => MUXB_SEL, Y(31) => 
                           mux_b_in_31_port, Y(30) => mux_b_in_30_port, Y(29) 
                           => mux_b_in_29_port, Y(28) => mux_b_in_28_port, 
                           Y(27) => mux_b_in_27_port, Y(26) => mux_b_in_26_port
                           , Y(25) => mux_b_in_25_port, Y(24) => 
                           mux_b_in_24_port, Y(23) => mux_b_in_23_port, Y(22) 
                           => mux_b_in_22_port, Y(21) => mux_b_in_21_port, 
                           Y(20) => mux_b_in_20_port, Y(19) => mux_b_in_19_port
                           , Y(18) => mux_b_in_18_port, Y(17) => 
                           mux_b_in_17_port, Y(16) => mux_b_in_16_port, Y(15) 
                           => mux_b_in_15_port, Y(14) => mux_b_in_14_port, 
                           Y(13) => mux_b_in_13_port, Y(12) => mux_b_in_12_port
                           , Y(11) => mux_b_in_11_port, Y(10) => 
                           mux_b_in_10_port, Y(9) => mux_b_in_9_port, Y(8) => 
                           mux_b_in_8_port, Y(7) => mux_b_in_7_port, Y(6) => 
                           mux_b_in_6_port, Y(5) => mux_b_in_5_port, Y(4) => 
                           mux_b_in_4_port, Y(3) => mux_b_in_3_port, Y(2) => 
                           mux_b_in_2_port, Y(1) => mux_b_in_1_port, Y(0) => 
                           mux_b_in_0_port);
   FORWARDING : FWD_UNIT port map( Rst => n16, Rs1(4) => Rs1_4_port, Rs1(3) => 
                           Rs1_3_port, Rs1(2) => Rs1_2_port, Rs1(1) => 
                           Rs1_1_port, Rs1(0) => Rs1_0_port, Rs2(4) => 
                           Rs2_4_port, Rs2(3) => Rs2_3_port, Rs2(2) => 
                           Rs2_2_port, Rs2(1) => Rs2_1_port, Rs2(0) => 
                           Rs2_0_port, Rd_M(4) => dest_M_4_port, Rd_M(3) => 
                           dest_M_3_port, Rd_M(2) => dest_M_2_port, Rd_M(1) => 
                           dest_M_1_port, Rd_M(0) => dest_M_0_port, Rd_W(4) => 
                           add_D_4_port, Rd_W(3) => add_D_3_port, Rd_W(2) => 
                           add_D_2_port, Rd_W(1) => add_D_1_port, Rd_W(0) => 
                           add_D_0_port, ICODE(5) => opcode_E_5_port, ICODE(4) 
                           => opcode_E_4_port, ICODE(3) => opcode_E_3_port, 
                           ICODE(2) => opcode_E_2_port, ICODE(1) => 
                           opcode_E_1_port, ICODE(0) => opcode_E_0_port, 
                           ICODE_M(5) => opcode_M_5_port, ICODE_M(4) => 
                           opcode_M_4_port, ICODE_M(3) => opcode_M_3_port, 
                           ICODE_M(2) => opcode_M_2_port, ICODE_M(1) => 
                           opcode_M_1_port, ICODE_M(0) => opcode_M_0_port, 
                           ICODE_W(5) => opcode_W_5_port, ICODE_W(4) => 
                           opcode_W_4_port, ICODE_W(3) => opcode_W_3_port, 
                           ICODE_W(2) => opcode_W_2_port, ICODE_W(1) => 
                           opcode_W_1_port, ICODE_W(0) => opcode_W_0_port, 
                           SEL_A(1) => FWD_MUX_A_S_1_port, SEL_A(0) => 
                           FWD_MUX_A_S_0_port, SEL_B(1) => FWD_MUX_B_S_1_port, 
                           SEL_B(0) => FWD_MUX_B_S_0_port);
   FWD_MUX_A : mux_3to1_N32_0 port map( A(31) => mux_a_in_31_port, A(30) => 
                           mux_a_in_30_port, A(29) => mux_a_in_29_port, A(28) 
                           => mux_a_in_28_port, A(27) => mux_a_in_27_port, 
                           A(26) => mux_a_in_26_port, A(25) => mux_a_in_25_port
                           , A(24) => mux_a_in_24_port, A(23) => 
                           mux_a_in_23_port, A(22) => mux_a_in_22_port, A(21) 
                           => mux_a_in_21_port, A(20) => mux_a_in_20_port, 
                           A(19) => mux_a_in_19_port, A(18) => mux_a_in_18_port
                           , A(17) => mux_a_in_17_port, A(16) => 
                           mux_a_in_16_port, A(15) => mux_a_in_15_port, A(14) 
                           => mux_a_in_14_port, A(13) => mux_a_in_13_port, 
                           A(12) => mux_a_in_12_port, A(11) => mux_a_in_11_port
                           , A(10) => mux_a_in_10_port, A(9) => mux_a_in_9_port
                           , A(8) => mux_a_in_8_port, A(7) => mux_a_in_7_port, 
                           A(6) => mux_a_in_6_port, A(5) => mux_a_in_5_port, 
                           A(4) => mux_a_in_4_port, A(3) => mux_a_in_3_port, 
                           A(2) => mux_a_in_2_port, A(1) => mux_a_in_1_port, 
                           A(0) => mux_a_in_0_port, B(31) => alu_out_M_31_port,
                           B(30) => alu_out_M_30_port, B(29) => 
                           alu_out_M_29_port, B(28) => alu_out_M_28_port, B(27)
                           => alu_out_M_27_port, B(26) => alu_out_M_26_port, 
                           B(25) => alu_out_M_25_port, B(24) => 
                           alu_out_M_24_port, B(23) => alu_out_M_23_port, B(22)
                           => alu_out_M_22_port, B(21) => alu_out_M_21_port, 
                           B(20) => alu_out_M_20_port, B(19) => 
                           alu_out_M_19_port, B(18) => alu_out_M_18_port, B(17)
                           => alu_out_M_17_port, B(16) => alu_out_M_16_port, 
                           B(15) => alu_out_M_15_port, B(14) => 
                           alu_out_M_14_port, B(13) => alu_out_M_13_port, B(12)
                           => alu_out_M_12_port, B(11) => DRAM_ADD_11_port, 
                           B(10) => DRAM_ADD_10_port, B(9) => DRAM_ADD_9_port, 
                           B(8) => DRAM_ADD_8_port, B(7) => DRAM_ADD_7_port, 
                           B(6) => DRAM_ADD_6_port, B(5) => DRAM_ADD_5_port, 
                           B(4) => DRAM_ADD_4_port, B(3) => DRAM_ADD_3_port, 
                           B(2) => DRAM_ADD_2_port, B(1) => DRAM_ADD_1_port, 
                           B(0) => DRAM_ADD_0_port, C(31) => alu_out_W_31_port,
                           C(30) => alu_out_W_30_port, C(29) => 
                           alu_out_W_29_port, C(28) => alu_out_W_28_port, C(27)
                           => alu_out_W_27_port, C(26) => alu_out_W_26_port, 
                           C(25) => alu_out_W_25_port, C(24) => 
                           alu_out_W_24_port, C(23) => alu_out_W_23_port, C(22)
                           => alu_out_W_22_port, C(21) => alu_out_W_21_port, 
                           C(20) => alu_out_W_20_port, C(19) => 
                           alu_out_W_19_port, C(18) => alu_out_W_18_port, C(17)
                           => alu_out_W_17_port, C(16) => alu_out_W_16_port, 
                           C(15) => alu_out_W_15_port, C(14) => 
                           alu_out_W_14_port, C(13) => alu_out_W_13_port, C(12)
                           => alu_out_W_12_port, C(11) => alu_out_W_11_port, 
                           C(10) => alu_out_W_10_port, C(9) => alu_out_W_9_port
                           , C(8) => alu_out_W_8_port, C(7) => alu_out_W_7_port
                           , C(6) => alu_out_W_6_port, C(5) => alu_out_W_5_port
                           , C(4) => alu_out_W_4_port, C(3) => alu_out_W_3_port
                           , C(2) => alu_out_W_2_port, C(1) => alu_out_W_1_port
                           , C(0) => alu_out_W_0_port, SEL(1) => 
                           FWD_MUX_A_S_1_port, SEL(0) => FWD_MUX_A_S_0_port, 
                           Y(31) => alu_a_in_31_port, Y(30) => alu_a_in_30_port
                           , Y(29) => alu_a_in_29_port, Y(28) => 
                           alu_a_in_28_port, Y(27) => alu_a_in_27_port, Y(26) 
                           => alu_a_in_26_port, Y(25) => alu_a_in_25_port, 
                           Y(24) => alu_a_in_24_port, Y(23) => alu_a_in_23_port
                           , Y(22) => alu_a_in_22_port, Y(21) => 
                           alu_a_in_21_port, Y(20) => alu_a_in_20_port, Y(19) 
                           => alu_a_in_19_port, Y(18) => alu_a_in_18_port, 
                           Y(17) => alu_a_in_17_port, Y(16) => alu_a_in_16_port
                           , Y(15) => alu_a_in_15_port, Y(14) => 
                           alu_a_in_14_port, Y(13) => alu_a_in_13_port, Y(12) 
                           => alu_a_in_12_port, Y(11) => alu_a_in_11_port, 
                           Y(10) => alu_a_in_10_port, Y(9) => alu_a_in_9_port, 
                           Y(8) => alu_a_in_8_port, Y(7) => alu_a_in_7_port, 
                           Y(6) => alu_a_in_6_port, Y(5) => alu_a_in_5_port, 
                           Y(4) => alu_a_in_4_port, Y(3) => alu_a_in_3_port, 
                           Y(2) => alu_a_in_2_port, Y(1) => alu_a_in_1_port, 
                           Y(0) => alu_a_in_0_port);
   FWD_MUX_B : mux_3to1_N32_3 port map( A(31) => mux_b_in_31_port, A(30) => 
                           mux_b_in_30_port, A(29) => mux_b_in_29_port, A(28) 
                           => mux_b_in_28_port, A(27) => mux_b_in_27_port, 
                           A(26) => mux_b_in_26_port, A(25) => mux_b_in_25_port
                           , A(24) => mux_b_in_24_port, A(23) => 
                           mux_b_in_23_port, A(22) => mux_b_in_22_port, A(21) 
                           => mux_b_in_21_port, A(20) => mux_b_in_20_port, 
                           A(19) => mux_b_in_19_port, A(18) => mux_b_in_18_port
                           , A(17) => mux_b_in_17_port, A(16) => 
                           mux_b_in_16_port, A(15) => mux_b_in_15_port, A(14) 
                           => mux_b_in_14_port, A(13) => mux_b_in_13_port, 
                           A(12) => mux_b_in_12_port, A(11) => mux_b_in_11_port
                           , A(10) => mux_b_in_10_port, A(9) => mux_b_in_9_port
                           , A(8) => mux_b_in_8_port, A(7) => mux_b_in_7_port, 
                           A(6) => mux_b_in_6_port, A(5) => mux_b_in_5_port, 
                           A(4) => mux_b_in_4_port, A(3) => mux_b_in_3_port, 
                           A(2) => mux_b_in_2_port, A(1) => mux_b_in_1_port, 
                           A(0) => mux_b_in_0_port, B(31) => alu_out_M_31_port,
                           B(30) => alu_out_M_30_port, B(29) => 
                           alu_out_M_29_port, B(28) => alu_out_M_28_port, B(27)
                           => alu_out_M_27_port, B(26) => alu_out_M_26_port, 
                           B(25) => alu_out_M_25_port, B(24) => 
                           alu_out_M_24_port, B(23) => alu_out_M_23_port, B(22)
                           => alu_out_M_22_port, B(21) => alu_out_M_21_port, 
                           B(20) => alu_out_M_20_port, B(19) => 
                           alu_out_M_19_port, B(18) => alu_out_M_18_port, B(17)
                           => alu_out_M_17_port, B(16) => alu_out_M_16_port, 
                           B(15) => alu_out_M_15_port, B(14) => 
                           alu_out_M_14_port, B(13) => alu_out_M_13_port, B(12)
                           => alu_out_M_12_port, B(11) => DRAM_ADD_11_port, 
                           B(10) => DRAM_ADD_10_port, B(9) => DRAM_ADD_9_port, 
                           B(8) => DRAM_ADD_8_port, B(7) => DRAM_ADD_7_port, 
                           B(6) => DRAM_ADD_6_port, B(5) => DRAM_ADD_5_port, 
                           B(4) => DRAM_ADD_4_port, B(3) => DRAM_ADD_3_port, 
                           B(2) => DRAM_ADD_2_port, B(1) => DRAM_ADD_1_port, 
                           B(0) => DRAM_ADD_0_port, C(31) => alu_out_W_31_port,
                           C(30) => alu_out_W_30_port, C(29) => 
                           alu_out_W_29_port, C(28) => alu_out_W_28_port, C(27)
                           => alu_out_W_27_port, C(26) => alu_out_W_26_port, 
                           C(25) => alu_out_W_25_port, C(24) => 
                           alu_out_W_24_port, C(23) => alu_out_W_23_port, C(22)
                           => alu_out_W_22_port, C(21) => alu_out_W_21_port, 
                           C(20) => alu_out_W_20_port, C(19) => 
                           alu_out_W_19_port, C(18) => alu_out_W_18_port, C(17)
                           => alu_out_W_17_port, C(16) => alu_out_W_16_port, 
                           C(15) => alu_out_W_15_port, C(14) => 
                           alu_out_W_14_port, C(13) => alu_out_W_13_port, C(12)
                           => alu_out_W_12_port, C(11) => alu_out_W_11_port, 
                           C(10) => alu_out_W_10_port, C(9) => alu_out_W_9_port
                           , C(8) => alu_out_W_8_port, C(7) => alu_out_W_7_port
                           , C(6) => alu_out_W_6_port, C(5) => alu_out_W_5_port
                           , C(4) => alu_out_W_4_port, C(3) => alu_out_W_3_port
                           , C(2) => alu_out_W_2_port, C(1) => alu_out_W_1_port
                           , C(0) => alu_out_W_0_port, SEL(1) => 
                           FWD_MUX_B_S_1_port, SEL(0) => FWD_MUX_B_S_0_port, 
                           Y(31) => alu_b_in_31_port, Y(30) => alu_b_in_30_port
                           , Y(29) => alu_b_in_29_port, Y(28) => 
                           alu_b_in_28_port, Y(27) => alu_b_in_27_port, Y(26) 
                           => alu_b_in_26_port, Y(25) => alu_b_in_25_port, 
                           Y(24) => alu_b_in_24_port, Y(23) => alu_b_in_23_port
                           , Y(22) => alu_b_in_22_port, Y(21) => 
                           alu_b_in_21_port, Y(20) => alu_b_in_20_port, Y(19) 
                           => alu_b_in_19_port, Y(18) => alu_b_in_18_port, 
                           Y(17) => alu_b_in_17_port, Y(16) => alu_b_in_16_port
                           , Y(15) => alu_b_in_15_port, Y(14) => 
                           alu_b_in_14_port, Y(13) => alu_b_in_13_port, Y(12) 
                           => alu_b_in_12_port, Y(11) => alu_b_in_11_port, 
                           Y(10) => alu_b_in_10_port, Y(9) => alu_b_in_9_port, 
                           Y(8) => alu_b_in_8_port, Y(7) => alu_b_in_7_port, 
                           Y(6) => alu_b_in_6_port, Y(5) => alu_b_in_5_port, 
                           Y(4) => alu_b_in_4_port, Y(3) => alu_b_in_3_port, 
                           Y(2) => alu_b_in_2_port, Y(1) => alu_b_in_1_port, 
                           Y(0) => alu_b_in_0_port);
   ALU_C : ALU_N32 port map( INA(31) => alu_a_in_31_port, INA(30) => 
                           alu_a_in_30_port, INA(29) => alu_a_in_29_port, 
                           INA(28) => alu_a_in_28_port, INA(27) => 
                           alu_a_in_27_port, INA(26) => alu_a_in_26_port, 
                           INA(25) => alu_a_in_25_port, INA(24) => 
                           alu_a_in_24_port, INA(23) => alu_a_in_23_port, 
                           INA(22) => alu_a_in_22_port, INA(21) => 
                           alu_a_in_21_port, INA(20) => alu_a_in_20_port, 
                           INA(19) => alu_a_in_19_port, INA(18) => 
                           alu_a_in_18_port, INA(17) => alu_a_in_17_port, 
                           INA(16) => alu_a_in_16_port, INA(15) => 
                           alu_a_in_15_port, INA(14) => alu_a_in_14_port, 
                           INA(13) => alu_a_in_13_port, INA(12) => 
                           alu_a_in_12_port, INA(11) => alu_a_in_11_port, 
                           INA(10) => alu_a_in_10_port, INA(9) => 
                           alu_a_in_9_port, INA(8) => alu_a_in_8_port, INA(7) 
                           => alu_a_in_7_port, INA(6) => alu_a_in_6_port, 
                           INA(5) => alu_a_in_5_port, INA(4) => alu_a_in_4_port
                           , INA(3) => alu_a_in_3_port, INA(2) => 
                           alu_a_in_2_port, INA(1) => alu_a_in_1_port, INA(0) 
                           => alu_a_in_0_port, INB(31) => alu_b_in_31_port, 
                           INB(30) => alu_b_in_30_port, INB(29) => 
                           alu_b_in_29_port, INB(28) => alu_b_in_28_port, 
                           INB(27) => alu_b_in_27_port, INB(26) => 
                           alu_b_in_26_port, INB(25) => alu_b_in_25_port, 
                           INB(24) => alu_b_in_24_port, INB(23) => 
                           alu_b_in_23_port, INB(22) => alu_b_in_22_port, 
                           INB(21) => alu_b_in_21_port, INB(20) => 
                           alu_b_in_20_port, INB(19) => alu_b_in_19_port, 
                           INB(18) => alu_b_in_18_port, INB(17) => 
                           alu_b_in_17_port, INB(16) => alu_b_in_16_port, 
                           INB(15) => alu_b_in_15_port, INB(14) => 
                           alu_b_in_14_port, INB(13) => alu_b_in_13_port, 
                           INB(12) => alu_b_in_12_port, INB(11) => 
                           alu_b_in_11_port, INB(10) => alu_b_in_10_port, 
                           INB(9) => alu_b_in_9_port, INB(8) => alu_b_in_8_port
                           , INB(7) => alu_b_in_7_port, INB(6) => 
                           alu_b_in_6_port, INB(5) => alu_b_in_5_port, INB(4) 
                           => alu_b_in_4_port, INB(3) => alu_b_in_3_port, 
                           INB(2) => alu_b_in_2_port, INB(1) => alu_b_in_1_port
                           , INB(0) => alu_b_in_0_port, OP(0) => ALU_OPCODE(0),
                           OP(1) => ALU_OPCODE(1), OP(2) => ALU_OPCODE(2), 
                           OP(3) => ALU_OPCODE(3), OP(4) => ALU_OPCODE(4), 
                           alu_out(31) => alu_out_31_port, alu_out(30) => 
                           alu_out_30_port, alu_out(29) => alu_out_29_port, 
                           alu_out(28) => alu_out_28_port, alu_out(27) => 
                           alu_out_27_port, alu_out(26) => alu_out_26_port, 
                           alu_out(25) => alu_out_25_port, alu_out(24) => 
                           alu_out_24_port, alu_out(23) => alu_out_23_port, 
                           alu_out(22) => alu_out_22_port, alu_out(21) => 
                           alu_out_21_port, alu_out(20) => alu_out_20_port, 
                           alu_out(19) => alu_out_19_port, alu_out(18) => 
                           alu_out_18_port, alu_out(17) => alu_out_17_port, 
                           alu_out(16) => alu_out_16_port, alu_out(15) => 
                           alu_out_15_port, alu_out(14) => alu_out_14_port, 
                           alu_out(13) => alu_out_13_port, alu_out(12) => 
                           alu_out_12_port, alu_out(11) => alu_out_11_port, 
                           alu_out(10) => alu_out_10_port, alu_out(9) => 
                           alu_out_9_port, alu_out(8) => alu_out_8_port, 
                           alu_out(7) => alu_out_7_port, alu_out(6) => 
                           alu_out_6_port, alu_out(5) => alu_out_5_port, 
                           alu_out(4) => alu_out_4_port, alu_out(3) => 
                           alu_out_3_port, alu_out(2) => alu_out_2_port, 
                           alu_out(1) => alu_out_1_port, alu_out(0) => 
                           alu_out_0_port);
   FORWARDING_BR : FWD_UNIT_BRANCH port map( Rst => n16, Rs1(4) => Rs1_4_port, 
                           Rs1(3) => Rs1_3_port, Rs1(2) => Rs1_2_port, Rs1(1) 
                           => Rs1_1_port, Rs1(0) => Rs1_0_port, Rd_M(4) => 
                           dest_M_4_port, Rd_M(3) => dest_M_3_port, Rd_M(2) => 
                           dest_M_2_port, Rd_M(1) => dest_M_1_port, Rd_M(0) => 
                           dest_M_0_port, Rd_W(4) => add_D_4_port, Rd_W(3) => 
                           add_D_3_port, Rd_W(2) => add_D_2_port, Rd_W(1) => 
                           add_D_1_port, Rd_W(0) => add_D_0_port, ICODE(5) => 
                           opcode_E_5_port, ICODE(4) => n9, ICODE(3) => n3, 
                           ICODE(2) => opcode_E_2_port, ICODE(1) => n13, 
                           ICODE(0) => n7, ICODE_M(5) => opcode_M_5_port, 
                           ICODE_M(4) => n8, ICODE_M(3) => n15, ICODE_M(2) => 
                           n5, ICODE_M(1) => n14, ICODE_M(0) => n10, ICODE_W(5)
                           => opcode_W_5_port, ICODE_W(4) => n11, ICODE_W(3) =>
                           n6, ICODE_W(2) => n4, ICODE_W(1) => n12, ICODE_W(0) 
                           => opcode_W_0_port, SEL(1) => FWD_MUX_BR_S_1_port, 
                           SEL(0) => FWD_MUX_BR_S_0_port);
   FWD_MUX_BRANCH : mux_3to1_N32_2 port map( A(31) => A_s_31_port, A(30) => 
                           A_s_30_port, A(29) => A_s_29_port, A(28) => 
                           A_s_28_port, A(27) => A_s_27_port, A(26) => 
                           A_s_26_port, A(25) => A_s_25_port, A(24) => 
                           A_s_24_port, A(23) => A_s_23_port, A(22) => 
                           A_s_22_port, A(21) => A_s_21_port, A(20) => 
                           A_s_20_port, A(19) => A_s_19_port, A(18) => 
                           A_s_18_port, A(17) => A_s_17_port, A(16) => 
                           A_s_16_port, A(15) => A_s_15_port, A(14) => 
                           A_s_14_port, A(13) => A_s_13_port, A(12) => 
                           A_s_12_port, A(11) => A_s_11_port, A(10) => 
                           A_s_10_port, A(9) => A_s_9_port, A(8) => A_s_8_port,
                           A(7) => A_s_7_port, A(6) => A_s_6_port, A(5) => 
                           A_s_5_port, A(4) => A_s_4_port, A(3) => A_s_3_port, 
                           A(2) => A_s_2_port, A(1) => A_s_1_port, A(0) => 
                           A_s_0_port, B(31) => alu_out_M_31_port, B(30) => 
                           alu_out_M_30_port, B(29) => alu_out_M_29_port, B(28)
                           => alu_out_M_28_port, B(27) => alu_out_M_27_port, 
                           B(26) => alu_out_M_26_port, B(25) => 
                           alu_out_M_25_port, B(24) => alu_out_M_24_port, B(23)
                           => alu_out_M_23_port, B(22) => alu_out_M_22_port, 
                           B(21) => alu_out_M_21_port, B(20) => 
                           alu_out_M_20_port, B(19) => alu_out_M_19_port, B(18)
                           => alu_out_M_18_port, B(17) => alu_out_M_17_port, 
                           B(16) => alu_out_M_16_port, B(15) => 
                           alu_out_M_15_port, B(14) => alu_out_M_14_port, B(13)
                           => alu_out_M_13_port, B(12) => alu_out_M_12_port, 
                           B(11) => DRAM_ADD_11_port, B(10) => DRAM_ADD_10_port
                           , B(9) => DRAM_ADD_9_port, B(8) => DRAM_ADD_8_port, 
                           B(7) => DRAM_ADD_7_port, B(6) => DRAM_ADD_6_port, 
                           B(5) => DRAM_ADD_5_port, B(4) => DRAM_ADD_4_port, 
                           B(3) => DRAM_ADD_3_port, B(2) => DRAM_ADD_2_port, 
                           B(1) => DRAM_ADD_1_port, B(0) => DRAM_ADD_0_port, 
                           C(31) => alu_out_W_31_port, C(30) => 
                           alu_out_W_30_port, C(29) => alu_out_W_29_port, C(28)
                           => alu_out_W_28_port, C(27) => alu_out_W_27_port, 
                           C(26) => alu_out_W_26_port, C(25) => 
                           alu_out_W_25_port, C(24) => alu_out_W_24_port, C(23)
                           => alu_out_W_23_port, C(22) => alu_out_W_22_port, 
                           C(21) => alu_out_W_21_port, C(20) => 
                           alu_out_W_20_port, C(19) => alu_out_W_19_port, C(18)
                           => alu_out_W_18_port, C(17) => alu_out_W_17_port, 
                           C(16) => alu_out_W_16_port, C(15) => 
                           alu_out_W_15_port, C(14) => alu_out_W_14_port, C(13)
                           => alu_out_W_13_port, C(12) => alu_out_W_12_port, 
                           C(11) => alu_out_W_11_port, C(10) => 
                           alu_out_W_10_port, C(9) => alu_out_W_9_port, C(8) =>
                           alu_out_W_8_port, C(7) => alu_out_W_7_port, C(6) => 
                           alu_out_W_6_port, C(5) => alu_out_W_5_port, C(4) => 
                           alu_out_W_4_port, C(3) => alu_out_W_3_port, C(2) => 
                           alu_out_W_2_port, C(1) => alu_out_W_1_port, C(0) => 
                           alu_out_W_0_port, SEL(1) => FWD_MUX_BR_S_1_port, 
                           SEL(0) => FWD_MUX_BR_S_0_port, Y(31) => 
                           br_mux_out_31_port, Y(30) => br_mux_out_30_port, 
                           Y(29) => br_mux_out_29_port, Y(28) => 
                           br_mux_out_28_port, Y(27) => br_mux_out_27_port, 
                           Y(26) => br_mux_out_26_port, Y(25) => 
                           br_mux_out_25_port, Y(24) => br_mux_out_24_port, 
                           Y(23) => br_mux_out_23_port, Y(22) => 
                           br_mux_out_22_port, Y(21) => br_mux_out_21_port, 
                           Y(20) => br_mux_out_20_port, Y(19) => 
                           br_mux_out_19_port, Y(18) => br_mux_out_18_port, 
                           Y(17) => br_mux_out_17_port, Y(16) => 
                           br_mux_out_16_port, Y(15) => br_mux_out_15_port, 
                           Y(14) => br_mux_out_14_port, Y(13) => 
                           br_mux_out_13_port, Y(12) => br_mux_out_12_port, 
                           Y(11) => br_mux_out_11_port, Y(10) => 
                           br_mux_out_10_port, Y(9) => br_mux_out_9_port, Y(8) 
                           => br_mux_out_8_port, Y(7) => br_mux_out_7_port, 
                           Y(6) => br_mux_out_6_port, Y(5) => br_mux_out_5_port
                           , Y(4) => br_mux_out_4_port, Y(3) => 
                           br_mux_out_3_port, Y(2) => br_mux_out_2_port, Y(1) 
                           => br_mux_out_1_port, Y(0) => br_mux_out_0_port);
   branch : branch_cond_N32 port map( A(31) => br_mux_out_31_port, A(30) => 
                           br_mux_out_30_port, A(29) => br_mux_out_29_port, 
                           A(28) => br_mux_out_28_port, A(27) => 
                           br_mux_out_27_port, A(26) => br_mux_out_26_port, 
                           A(25) => br_mux_out_25_port, A(24) => 
                           br_mux_out_24_port, A(23) => br_mux_out_23_port, 
                           A(22) => br_mux_out_22_port, A(21) => 
                           br_mux_out_21_port, A(20) => br_mux_out_20_port, 
                           A(19) => br_mux_out_19_port, A(18) => 
                           br_mux_out_18_port, A(17) => br_mux_out_17_port, 
                           A(16) => br_mux_out_16_port, A(15) => 
                           br_mux_out_15_port, A(14) => br_mux_out_14_port, 
                           A(13) => br_mux_out_13_port, A(12) => 
                           br_mux_out_12_port, A(11) => br_mux_out_11_port, 
                           A(10) => br_mux_out_10_port, A(9) => 
                           br_mux_out_9_port, A(8) => br_mux_out_8_port, A(7) 
                           => br_mux_out_7_port, A(6) => br_mux_out_6_port, 
                           A(5) => br_mux_out_5_port, A(4) => br_mux_out_4_port
                           , A(3) => br_mux_out_3_port, A(2) => 
                           br_mux_out_2_port, A(1) => br_mux_out_1_port, A(0) 
                           => br_mux_out_0_port, EN => BR_EN, OP(0) => 
                           ALU_OPCODE(0), OP(1) => ALU_OPCODE(1), OP(2) => 
                           ALU_OPCODE(2), OP(3) => n2, OP(4) => ALU_OPCODE(4), 
                           PRE => pr_E, DISCARD => discard_s, WRONG => wrong_br
                           , RIGHT => right_br, SEL => jr_sel);
   EX_MEM_s : EX_MEM port map( CLK => Clk, RST => n16, NPC_IN(31) => 
                           npc_E_31_port, NPC_IN(30) => npc_E_30_port, 
                           NPC_IN(29) => npc_E_29_port, NPC_IN(28) => 
                           npc_E_28_port, NPC_IN(27) => npc_E_27_port, 
                           NPC_IN(26) => npc_E_26_port, NPC_IN(25) => 
                           npc_E_25_port, NPC_IN(24) => npc_E_24_port, 
                           NPC_IN(23) => npc_E_23_port, NPC_IN(22) => 
                           npc_E_22_port, NPC_IN(21) => npc_E_21_port, 
                           NPC_IN(20) => npc_E_20_port, NPC_IN(19) => 
                           npc_E_19_port, NPC_IN(18) => npc_E_18_port, 
                           NPC_IN(17) => npc_E_17_port, NPC_IN(16) => 
                           npc_E_16_port, NPC_IN(15) => npc_E_15_port, 
                           NPC_IN(14) => npc_E_14_port, NPC_IN(13) => 
                           npc_E_13_port, NPC_IN(12) => npc_E_12_port, 
                           NPC_IN(11) => npc_E_11_port, NPC_IN(10) => 
                           npc_E_10_port, NPC_IN(9) => npc_E_9_port, NPC_IN(8) 
                           => npc_E_8_port, NPC_IN(7) => npc_E_7_port, 
                           NPC_IN(6) => npc_E_6_port, NPC_IN(5) => npc_E_5_port
                           , NPC_IN(4) => npc_E_4_port, NPC_IN(3) => 
                           npc_E_3_port, NPC_IN(2) => npc_E_2_port, NPC_IN(1) 
                           => npc_E_1_port, NPC_IN(0) => npc_E_0_port, 
                           NPC_L_IN(31) => link_addr_E_31_port, NPC_L_IN(30) =>
                           link_addr_E_30_port, NPC_L_IN(29) => 
                           link_addr_E_29_port, NPC_L_IN(28) => 
                           link_addr_E_28_port, NPC_L_IN(27) => 
                           link_addr_E_27_port, NPC_L_IN(26) => 
                           link_addr_E_26_port, NPC_L_IN(25) => 
                           link_addr_E_25_port, NPC_L_IN(24) => 
                           link_addr_E_24_port, NPC_L_IN(23) => 
                           link_addr_E_23_port, NPC_L_IN(22) => 
                           link_addr_E_22_port, NPC_L_IN(21) => 
                           link_addr_E_21_port, NPC_L_IN(20) => 
                           link_addr_E_20_port, NPC_L_IN(19) => 
                           link_addr_E_19_port, NPC_L_IN(18) => 
                           link_addr_E_18_port, NPC_L_IN(17) => 
                           link_addr_E_17_port, NPC_L_IN(16) => 
                           link_addr_E_16_port, NPC_L_IN(15) => 
                           link_addr_E_15_port, NPC_L_IN(14) => 
                           link_addr_E_14_port, NPC_L_IN(13) => 
                           link_addr_E_13_port, NPC_L_IN(12) => 
                           link_addr_E_12_port, NPC_L_IN(11) => 
                           link_addr_E_11_port, NPC_L_IN(10) => 
                           link_addr_E_10_port, NPC_L_IN(9) => 
                           link_addr_E_9_port, NPC_L_IN(8) => 
                           link_addr_E_8_port, NPC_L_IN(7) => 
                           link_addr_E_7_port, NPC_L_IN(6) => 
                           link_addr_E_6_port, NPC_L_IN(5) => 
                           link_addr_E_5_port, NPC_L_IN(4) => 
                           link_addr_E_4_port, NPC_L_IN(3) => 
                           link_addr_E_3_port, NPC_L_IN(2) => 
                           link_addr_E_2_port, NPC_L_IN(1) => 
                           link_addr_E_1_port, NPC_L_IN(0) => 
                           link_addr_E_0_port, ALU_IN(31) => alu_out_31_port, 
                           ALU_IN(30) => alu_out_30_port, ALU_IN(29) => n1, 
                           ALU_IN(28) => alu_out_28_port, ALU_IN(27) => 
                           alu_out_27_port, ALU_IN(26) => alu_out_26_port, 
                           ALU_IN(25) => alu_out_25_port, ALU_IN(24) => 
                           alu_out_24_port, ALU_IN(23) => alu_out_23_port, 
                           ALU_IN(22) => alu_out_22_port, ALU_IN(21) => 
                           alu_out_21_port, ALU_IN(20) => alu_out_20_port, 
                           ALU_IN(19) => alu_out_19_port, ALU_IN(18) => 
                           alu_out_18_port, ALU_IN(17) => alu_out_17_port, 
                           ALU_IN(16) => alu_out_16_port, ALU_IN(15) => 
                           alu_out_15_port, ALU_IN(14) => alu_out_14_port, 
                           ALU_IN(13) => alu_out_13_port, ALU_IN(12) => 
                           alu_out_12_port, ALU_IN(11) => alu_out_11_port, 
                           ALU_IN(10) => alu_out_10_port, ALU_IN(9) => 
                           alu_out_9_port, ALU_IN(8) => alu_out_8_port, 
                           ALU_IN(7) => alu_out_7_port, ALU_IN(6) => 
                           alu_out_6_port, ALU_IN(5) => alu_out_5_port, 
                           ALU_IN(4) => alu_out_4_port, ALU_IN(3) => 
                           alu_out_3_port, ALU_IN(2) => alu_out_2_port, 
                           ALU_IN(1) => alu_out_1_port, ALU_IN(0) => 
                           alu_out_0_port, B_IN(31) => B_s_31_port, B_IN(30) =>
                           B_s_30_port, B_IN(29) => B_s_29_port, B_IN(28) => 
                           B_s_28_port, B_IN(27) => B_s_27_port, B_IN(26) => 
                           B_s_26_port, B_IN(25) => B_s_25_port, B_IN(24) => 
                           B_s_24_port, B_IN(23) => B_s_23_port, B_IN(22) => 
                           B_s_22_port, B_IN(21) => B_s_21_port, B_IN(20) => 
                           B_s_20_port, B_IN(19) => B_s_19_port, B_IN(18) => 
                           B_s_18_port, B_IN(17) => B_s_17_port, B_IN(16) => 
                           B_s_16_port, B_IN(15) => B_s_15_port, B_IN(14) => 
                           B_s_14_port, B_IN(13) => B_s_13_port, B_IN(12) => 
                           B_s_12_port, B_IN(11) => B_s_11_port, B_IN(10) => 
                           B_s_10_port, B_IN(9) => B_s_9_port, B_IN(8) => 
                           B_s_8_port, B_IN(7) => B_s_7_port, B_IN(6) => 
                           B_s_6_port, B_IN(5) => B_s_5_port, B_IN(4) => 
                           B_s_4_port, B_IN(3) => B_s_3_port, B_IN(2) => 
                           B_s_2_port, B_IN(1) => B_s_1_port, B_IN(0) => 
                           B_s_0_port, RD_IN(4) => dest_E_4_port, RD_IN(3) => 
                           dest_E_3_port, RD_IN(2) => dest_E_2_port, RD_IN(1) 
                           => dest_E_1_port, RD_IN(0) => dest_E_0_port, 
                           OPCODE_IN(5) => opcode_E_5_port, OPCODE_IN(4) => n9,
                           OPCODE_IN(3) => n3, OPCODE_IN(2) => opcode_E_2_port,
                           OPCODE_IN(1) => n13, OPCODE_IN(0) => n7, NPC_OUT(31)
                           => npc_M_31_port, NPC_OUT(30) => npc_M_30_port, 
                           NPC_OUT(29) => npc_M_29_port, NPC_OUT(28) => 
                           npc_M_28_port, NPC_OUT(27) => npc_M_27_port, 
                           NPC_OUT(26) => npc_M_26_port, NPC_OUT(25) => 
                           npc_M_25_port, NPC_OUT(24) => npc_M_24_port, 
                           NPC_OUT(23) => npc_M_23_port, NPC_OUT(22) => 
                           npc_M_22_port, NPC_OUT(21) => npc_M_21_port, 
                           NPC_OUT(20) => npc_M_20_port, NPC_OUT(19) => 
                           npc_M_19_port, NPC_OUT(18) => npc_M_18_port, 
                           NPC_OUT(17) => npc_M_17_port, NPC_OUT(16) => 
                           npc_M_16_port, NPC_OUT(15) => npc_M_15_port, 
                           NPC_OUT(14) => npc_M_14_port, NPC_OUT(13) => 
                           npc_M_13_port, NPC_OUT(12) => npc_M_12_port, 
                           NPC_OUT(11) => npc_M_11_port, NPC_OUT(10) => 
                           npc_M_10_port, NPC_OUT(9) => npc_M_9_port, 
                           NPC_OUT(8) => npc_M_8_port, NPC_OUT(7) => 
                           npc_M_7_port, NPC_OUT(6) => npc_M_6_port, NPC_OUT(5)
                           => npc_M_5_port, NPC_OUT(4) => npc_M_4_port, 
                           NPC_OUT(3) => npc_M_3_port, NPC_OUT(2) => 
                           npc_M_2_port, NPC_OUT(1) => npc_M_1_port, NPC_OUT(0)
                           => npc_M_0_port, NPC_L_OUT(31) => 
                           link_addr_M_31_port, NPC_L_OUT(30) => 
                           link_addr_M_30_port, NPC_L_OUT(29) => 
                           link_addr_M_29_port, NPC_L_OUT(28) => 
                           link_addr_M_28_port, NPC_L_OUT(27) => 
                           link_addr_M_27_port, NPC_L_OUT(26) => 
                           link_addr_M_26_port, NPC_L_OUT(25) => 
                           link_addr_M_25_port, NPC_L_OUT(24) => 
                           link_addr_M_24_port, NPC_L_OUT(23) => 
                           link_addr_M_23_port, NPC_L_OUT(22) => 
                           link_addr_M_22_port, NPC_L_OUT(21) => 
                           link_addr_M_21_port, NPC_L_OUT(20) => 
                           link_addr_M_20_port, NPC_L_OUT(19) => 
                           link_addr_M_19_port, NPC_L_OUT(18) => 
                           link_addr_M_18_port, NPC_L_OUT(17) => 
                           link_addr_M_17_port, NPC_L_OUT(16) => 
                           link_addr_M_16_port, NPC_L_OUT(15) => 
                           link_addr_M_15_port, NPC_L_OUT(14) => 
                           link_addr_M_14_port, NPC_L_OUT(13) => 
                           link_addr_M_13_port, NPC_L_OUT(12) => 
                           link_addr_M_12_port, NPC_L_OUT(11) => 
                           link_addr_M_11_port, NPC_L_OUT(10) => 
                           link_addr_M_10_port, NPC_L_OUT(9) => 
                           link_addr_M_9_port, NPC_L_OUT(8) => 
                           link_addr_M_8_port, NPC_L_OUT(7) => 
                           link_addr_M_7_port, NPC_L_OUT(6) => 
                           link_addr_M_6_port, NPC_L_OUT(5) => 
                           link_addr_M_5_port, NPC_L_OUT(4) => 
                           link_addr_M_4_port, NPC_L_OUT(3) => 
                           link_addr_M_3_port, NPC_L_OUT(2) => 
                           link_addr_M_2_port, NPC_L_OUT(1) => 
                           link_addr_M_1_port, NPC_L_OUT(0) => 
                           link_addr_M_0_port, ALU_OUT(31) => alu_out_M_31_port
                           , ALU_OUT(30) => alu_out_M_30_port, ALU_OUT(29) => 
                           alu_out_M_29_port, ALU_OUT(28) => alu_out_M_28_port,
                           ALU_OUT(27) => alu_out_M_27_port, ALU_OUT(26) => 
                           alu_out_M_26_port, ALU_OUT(25) => alu_out_M_25_port,
                           ALU_OUT(24) => alu_out_M_24_port, ALU_OUT(23) => 
                           alu_out_M_23_port, ALU_OUT(22) => alu_out_M_22_port,
                           ALU_OUT(21) => alu_out_M_21_port, ALU_OUT(20) => 
                           alu_out_M_20_port, ALU_OUT(19) => alu_out_M_19_port,
                           ALU_OUT(18) => alu_out_M_18_port, ALU_OUT(17) => 
                           alu_out_M_17_port, ALU_OUT(16) => alu_out_M_16_port,
                           ALU_OUT(15) => alu_out_M_15_port, ALU_OUT(14) => 
                           alu_out_M_14_port, ALU_OUT(13) => alu_out_M_13_port,
                           ALU_OUT(12) => alu_out_M_12_port, ALU_OUT(11) => 
                           DRAM_ADD_11_port, ALU_OUT(10) => DRAM_ADD_10_port, 
                           ALU_OUT(9) => DRAM_ADD_9_port, ALU_OUT(8) => 
                           DRAM_ADD_8_port, ALU_OUT(7) => DRAM_ADD_7_port, 
                           ALU_OUT(6) => DRAM_ADD_6_port, ALU_OUT(5) => 
                           DRAM_ADD_5_port, ALU_OUT(4) => DRAM_ADD_4_port, 
                           ALU_OUT(3) => DRAM_ADD_3_port, ALU_OUT(2) => 
                           DRAM_ADD_2_port, ALU_OUT(1) => DRAM_ADD_1_port, 
                           ALU_OUT(0) => DRAM_ADD_0_port, B_OUT(31) => 
                           DRAM_IN(31), B_OUT(30) => DRAM_IN(30), B_OUT(29) => 
                           DRAM_IN(29), B_OUT(28) => DRAM_IN(28), B_OUT(27) => 
                           DRAM_IN(27), B_OUT(26) => DRAM_IN(26), B_OUT(25) => 
                           DRAM_IN(25), B_OUT(24) => DRAM_IN(24), B_OUT(23) => 
                           DRAM_IN(23), B_OUT(22) => DRAM_IN(22), B_OUT(21) => 
                           DRAM_IN(21), B_OUT(20) => DRAM_IN(20), B_OUT(19) => 
                           DRAM_IN(19), B_OUT(18) => DRAM_IN(18), B_OUT(17) => 
                           DRAM_IN(17), B_OUT(16) => DRAM_IN(16), B_OUT(15) => 
                           DRAM_IN(15), B_OUT(14) => DRAM_IN(14), B_OUT(13) => 
                           DRAM_IN(13), B_OUT(12) => DRAM_IN(12), B_OUT(11) => 
                           DRAM_IN(11), B_OUT(10) => DRAM_IN(10), B_OUT(9) => 
                           DRAM_IN(9), B_OUT(8) => DRAM_IN(8), B_OUT(7) => 
                           DRAM_IN(7), B_OUT(6) => DRAM_IN(6), B_OUT(5) => 
                           DRAM_IN(5), B_OUT(4) => DRAM_IN(4), B_OUT(3) => 
                           DRAM_IN(3), B_OUT(2) => DRAM_IN(2), B_OUT(1) => 
                           DRAM_IN(1), B_OUT(0) => DRAM_IN(0), RD_OUT(4) => 
                           dest_M_4_port, RD_OUT(3) => dest_M_3_port, RD_OUT(2)
                           => dest_M_2_port, RD_OUT(1) => dest_M_1_port, 
                           RD_OUT(0) => dest_M_0_port, OPCODE_OUT(5) => 
                           opcode_M_5_port, OPCODE_OUT(4) => opcode_M_4_port, 
                           OPCODE_OUT(3) => opcode_M_3_port, OPCODE_OUT(2) => 
                           opcode_M_2_port, OPCODE_OUT(1) => opcode_M_1_port, 
                           OPCODE_OUT(0) => opcode_M_0_port);
   MEM_WB_s : MEM_WB port map( CLK => Clk, RST => n16, NPC_L_IN(31) => 
                           link_addr_M_31_port, NPC_L_IN(30) => 
                           link_addr_M_30_port, NPC_L_IN(29) => 
                           link_addr_M_29_port, NPC_L_IN(28) => 
                           link_addr_M_28_port, NPC_L_IN(27) => 
                           link_addr_M_27_port, NPC_L_IN(26) => 
                           link_addr_M_26_port, NPC_L_IN(25) => 
                           link_addr_M_25_port, NPC_L_IN(24) => 
                           link_addr_M_24_port, NPC_L_IN(23) => 
                           link_addr_M_23_port, NPC_L_IN(22) => 
                           link_addr_M_22_port, NPC_L_IN(21) => 
                           link_addr_M_21_port, NPC_L_IN(20) => 
                           link_addr_M_20_port, NPC_L_IN(19) => 
                           link_addr_M_19_port, NPC_L_IN(18) => 
                           link_addr_M_18_port, NPC_L_IN(17) => 
                           link_addr_M_17_port, NPC_L_IN(16) => 
                           link_addr_M_16_port, NPC_L_IN(15) => 
                           link_addr_M_15_port, NPC_L_IN(14) => 
                           link_addr_M_14_port, NPC_L_IN(13) => 
                           link_addr_M_13_port, NPC_L_IN(12) => 
                           link_addr_M_12_port, NPC_L_IN(11) => 
                           link_addr_M_11_port, NPC_L_IN(10) => 
                           link_addr_M_10_port, NPC_L_IN(9) => 
                           link_addr_M_9_port, NPC_L_IN(8) => 
                           link_addr_M_8_port, NPC_L_IN(7) => 
                           link_addr_M_7_port, NPC_L_IN(6) => 
                           link_addr_M_6_port, NPC_L_IN(5) => 
                           link_addr_M_5_port, NPC_L_IN(4) => 
                           link_addr_M_4_port, NPC_L_IN(3) => 
                           link_addr_M_3_port, NPC_L_IN(2) => 
                           link_addr_M_2_port, NPC_L_IN(1) => 
                           link_addr_M_1_port, NPC_L_IN(0) => 
                           link_addr_M_0_port, ALU_IN(31) => alu_out_M_31_port,
                           ALU_IN(30) => alu_out_M_30_port, ALU_IN(29) => 
                           alu_out_M_29_port, ALU_IN(28) => alu_out_M_28_port, 
                           ALU_IN(27) => alu_out_M_27_port, ALU_IN(26) => 
                           alu_out_M_26_port, ALU_IN(25) => alu_out_M_25_port, 
                           ALU_IN(24) => alu_out_M_24_port, ALU_IN(23) => 
                           alu_out_M_23_port, ALU_IN(22) => alu_out_M_22_port, 
                           ALU_IN(21) => alu_out_M_21_port, ALU_IN(20) => 
                           alu_out_M_20_port, ALU_IN(19) => alu_out_M_19_port, 
                           ALU_IN(18) => alu_out_M_18_port, ALU_IN(17) => 
                           alu_out_M_17_port, ALU_IN(16) => alu_out_M_16_port, 
                           ALU_IN(15) => alu_out_M_15_port, ALU_IN(14) => 
                           alu_out_M_14_port, ALU_IN(13) => alu_out_M_13_port, 
                           ALU_IN(12) => alu_out_M_12_port, ALU_IN(11) => 
                           DRAM_ADD_11_port, ALU_IN(10) => DRAM_ADD_10_port, 
                           ALU_IN(9) => DRAM_ADD_9_port, ALU_IN(8) => 
                           DRAM_ADD_8_port, ALU_IN(7) => DRAM_ADD_7_port, 
                           ALU_IN(6) => DRAM_ADD_6_port, ALU_IN(5) => 
                           DRAM_ADD_5_port, ALU_IN(4) => DRAM_ADD_4_port, 
                           ALU_IN(3) => DRAM_ADD_3_port, ALU_IN(2) => 
                           DRAM_ADD_2_port, ALU_IN(1) => DRAM_ADD_1_port, 
                           ALU_IN(0) => DRAM_ADD_0_port, LMD_IN(31) => 
                           DRAM_OUT(31), LMD_IN(30) => DRAM_OUT(30), LMD_IN(29)
                           => DRAM_OUT(29), LMD_IN(28) => DRAM_OUT(28), 
                           LMD_IN(27) => DRAM_OUT(27), LMD_IN(26) => 
                           DRAM_OUT(26), LMD_IN(25) => DRAM_OUT(25), LMD_IN(24)
                           => DRAM_OUT(24), LMD_IN(23) => DRAM_OUT(23), 
                           LMD_IN(22) => DRAM_OUT(22), LMD_IN(21) => 
                           DRAM_OUT(21), LMD_IN(20) => DRAM_OUT(20), LMD_IN(19)
                           => DRAM_OUT(19), LMD_IN(18) => DRAM_OUT(18), 
                           LMD_IN(17) => DRAM_OUT(17), LMD_IN(16) => 
                           DRAM_OUT(16), LMD_IN(15) => DRAM_OUT(15), LMD_IN(14)
                           => DRAM_OUT(14), LMD_IN(13) => DRAM_OUT(13), 
                           LMD_IN(12) => DRAM_OUT(12), LMD_IN(11) => 
                           DRAM_OUT(11), LMD_IN(10) => DRAM_OUT(10), LMD_IN(9) 
                           => DRAM_OUT(9), LMD_IN(8) => DRAM_OUT(8), LMD_IN(7) 
                           => DRAM_OUT(7), LMD_IN(6) => DRAM_OUT(6), LMD_IN(5) 
                           => DRAM_OUT(5), LMD_IN(4) => DRAM_OUT(4), LMD_IN(3) 
                           => DRAM_OUT(3), LMD_IN(2) => DRAM_OUT(2), LMD_IN(1) 
                           => DRAM_OUT(1), LMD_IN(0) => DRAM_OUT(0), RD_IN(4) 
                           => dest_M_4_port, RD_IN(3) => dest_M_3_port, 
                           RD_IN(2) => dest_M_2_port, RD_IN(1) => dest_M_1_port
                           , RD_IN(0) => dest_M_0_port, OPCODE_IN(5) => 
                           opcode_M_5_port, OPCODE_IN(4) => opcode_M_4_port, 
                           OPCODE_IN(3) => n15, OPCODE_IN(2) => n5, 
                           OPCODE_IN(1) => n14, OPCODE_IN(0) => n10, 
                           NPC_L_OUT(31) => link_addr_W_31_port, NPC_L_OUT(30) 
                           => link_addr_W_30_port, NPC_L_OUT(29) => 
                           link_addr_W_29_port, NPC_L_OUT(28) => 
                           link_addr_W_28_port, NPC_L_OUT(27) => 
                           link_addr_W_27_port, NPC_L_OUT(26) => 
                           link_addr_W_26_port, NPC_L_OUT(25) => 
                           link_addr_W_25_port, NPC_L_OUT(24) => 
                           link_addr_W_24_port, NPC_L_OUT(23) => 
                           link_addr_W_23_port, NPC_L_OUT(22) => 
                           link_addr_W_22_port, NPC_L_OUT(21) => 
                           link_addr_W_21_port, NPC_L_OUT(20) => 
                           link_addr_W_20_port, NPC_L_OUT(19) => 
                           link_addr_W_19_port, NPC_L_OUT(18) => 
                           link_addr_W_18_port, NPC_L_OUT(17) => 
                           link_addr_W_17_port, NPC_L_OUT(16) => 
                           link_addr_W_16_port, NPC_L_OUT(15) => 
                           link_addr_W_15_port, NPC_L_OUT(14) => 
                           link_addr_W_14_port, NPC_L_OUT(13) => 
                           link_addr_W_13_port, NPC_L_OUT(12) => 
                           link_addr_W_12_port, NPC_L_OUT(11) => 
                           link_addr_W_11_port, NPC_L_OUT(10) => 
                           link_addr_W_10_port, NPC_L_OUT(9) => 
                           link_addr_W_9_port, NPC_L_OUT(8) => 
                           link_addr_W_8_port, NPC_L_OUT(7) => 
                           link_addr_W_7_port, NPC_L_OUT(6) => 
                           link_addr_W_6_port, NPC_L_OUT(5) => 
                           link_addr_W_5_port, NPC_L_OUT(4) => 
                           link_addr_W_4_port, NPC_L_OUT(3) => 
                           link_addr_W_3_port, NPC_L_OUT(2) => 
                           link_addr_W_2_port, NPC_L_OUT(1) => 
                           link_addr_W_1_port, NPC_L_OUT(0) => 
                           link_addr_W_0_port, ALU_OUT(31) => alu_out_W_31_port
                           , ALU_OUT(30) => alu_out_W_30_port, ALU_OUT(29) => 
                           alu_out_W_29_port, ALU_OUT(28) => alu_out_W_28_port,
                           ALU_OUT(27) => alu_out_W_27_port, ALU_OUT(26) => 
                           alu_out_W_26_port, ALU_OUT(25) => alu_out_W_25_port,
                           ALU_OUT(24) => alu_out_W_24_port, ALU_OUT(23) => 
                           alu_out_W_23_port, ALU_OUT(22) => alu_out_W_22_port,
                           ALU_OUT(21) => alu_out_W_21_port, ALU_OUT(20) => 
                           alu_out_W_20_port, ALU_OUT(19) => alu_out_W_19_port,
                           ALU_OUT(18) => alu_out_W_18_port, ALU_OUT(17) => 
                           alu_out_W_17_port, ALU_OUT(16) => alu_out_W_16_port,
                           ALU_OUT(15) => alu_out_W_15_port, ALU_OUT(14) => 
                           alu_out_W_14_port, ALU_OUT(13) => alu_out_W_13_port,
                           ALU_OUT(12) => alu_out_W_12_port, ALU_OUT(11) => 
                           alu_out_W_11_port, ALU_OUT(10) => alu_out_W_10_port,
                           ALU_OUT(9) => alu_out_W_9_port, ALU_OUT(8) => 
                           alu_out_W_8_port, ALU_OUT(7) => alu_out_W_7_port, 
                           ALU_OUT(6) => alu_out_W_6_port, ALU_OUT(5) => 
                           alu_out_W_5_port, ALU_OUT(4) => alu_out_W_4_port, 
                           ALU_OUT(3) => alu_out_W_3_port, ALU_OUT(2) => 
                           alu_out_W_2_port, ALU_OUT(1) => alu_out_W_1_port, 
                           ALU_OUT(0) => alu_out_W_0_port, LMD_OUT(31) => 
                           LMD_out_31_port, LMD_OUT(30) => LMD_out_30_port, 
                           LMD_OUT(29) => LMD_out_29_port, LMD_OUT(28) => 
                           LMD_out_28_port, LMD_OUT(27) => LMD_out_27_port, 
                           LMD_OUT(26) => LMD_out_26_port, LMD_OUT(25) => 
                           LMD_out_25_port, LMD_OUT(24) => LMD_out_24_port, 
                           LMD_OUT(23) => LMD_out_23_port, LMD_OUT(22) => 
                           LMD_out_22_port, LMD_OUT(21) => LMD_out_21_port, 
                           LMD_OUT(20) => LMD_out_20_port, LMD_OUT(19) => 
                           LMD_out_19_port, LMD_OUT(18) => LMD_out_18_port, 
                           LMD_OUT(17) => LMD_out_17_port, LMD_OUT(16) => 
                           LMD_out_16_port, LMD_OUT(15) => LMD_out_15_port, 
                           LMD_OUT(14) => LMD_out_14_port, LMD_OUT(13) => 
                           LMD_out_13_port, LMD_OUT(12) => LMD_out_12_port, 
                           LMD_OUT(11) => LMD_out_11_port, LMD_OUT(10) => 
                           LMD_out_10_port, LMD_OUT(9) => LMD_out_9_port, 
                           LMD_OUT(8) => LMD_out_8_port, LMD_OUT(7) => 
                           LMD_out_7_port, LMD_OUT(6) => LMD_out_6_port, 
                           LMD_OUT(5) => LMD_out_5_port, LMD_OUT(4) => 
                           LMD_out_4_port, LMD_OUT(3) => LMD_out_3_port, 
                           LMD_OUT(2) => LMD_out_2_port, LMD_OUT(1) => 
                           LMD_out_1_port, LMD_OUT(0) => LMD_out_0_port, 
                           RD_OUT(4) => add_D_4_port, RD_OUT(3) => add_D_3_port
                           , RD_OUT(2) => add_D_2_port, RD_OUT(1) => 
                           add_D_1_port, RD_OUT(0) => add_D_0_port, 
                           OPCODE_OUT(5) => opcode_W_5_port, OPCODE_OUT(4) => 
                           opcode_W_4_port, OPCODE_OUT(3) => opcode_W_3_port, 
                           OPCODE_OUT(2) => opcode_W_2_port, OPCODE_OUT(1) => 
                           opcode_W_1_port, OPCODE_OUT(0) => opcode_W_0_port);
   RF_in_mux : mux_3to1_N32_1 port map( A(31) => alu_out_W_31_port, A(30) => 
                           alu_out_W_30_port, A(29) => alu_out_W_29_port, A(28)
                           => alu_out_W_28_port, A(27) => alu_out_W_27_port, 
                           A(26) => alu_out_W_26_port, A(25) => 
                           alu_out_W_25_port, A(24) => alu_out_W_24_port, A(23)
                           => alu_out_W_23_port, A(22) => alu_out_W_22_port, 
                           A(21) => alu_out_W_21_port, A(20) => 
                           alu_out_W_20_port, A(19) => alu_out_W_19_port, A(18)
                           => alu_out_W_18_port, A(17) => alu_out_W_17_port, 
                           A(16) => alu_out_W_16_port, A(15) => 
                           alu_out_W_15_port, A(14) => alu_out_W_14_port, A(13)
                           => alu_out_W_13_port, A(12) => alu_out_W_12_port, 
                           A(11) => alu_out_W_11_port, A(10) => 
                           alu_out_W_10_port, A(9) => alu_out_W_9_port, A(8) =>
                           alu_out_W_8_port, A(7) => alu_out_W_7_port, A(6) => 
                           alu_out_W_6_port, A(5) => alu_out_W_5_port, A(4) => 
                           alu_out_W_4_port, A(3) => alu_out_W_3_port, A(2) => 
                           alu_out_W_2_port, A(1) => alu_out_W_1_port, A(0) => 
                           alu_out_W_0_port, B(31) => LMD_out_31_port, B(30) =>
                           LMD_out_30_port, B(29) => LMD_out_29_port, B(28) => 
                           LMD_out_28_port, B(27) => LMD_out_27_port, B(26) => 
                           LMD_out_26_port, B(25) => LMD_out_25_port, B(24) => 
                           LMD_out_24_port, B(23) => LMD_out_23_port, B(22) => 
                           LMD_out_22_port, B(21) => LMD_out_21_port, B(20) => 
                           LMD_out_20_port, B(19) => LMD_out_19_port, B(18) => 
                           LMD_out_18_port, B(17) => LMD_out_17_port, B(16) => 
                           LMD_out_16_port, B(15) => LMD_out_15_port, B(14) => 
                           LMD_out_14_port, B(13) => LMD_out_13_port, B(12) => 
                           LMD_out_12_port, B(11) => LMD_out_11_port, B(10) => 
                           LMD_out_10_port, B(9) => LMD_out_9_port, B(8) => 
                           LMD_out_8_port, B(7) => LMD_out_7_port, B(6) => 
                           LMD_out_6_port, B(5) => LMD_out_5_port, B(4) => 
                           LMD_out_4_port, B(3) => LMD_out_3_port, B(2) => 
                           LMD_out_2_port, B(1) => LMD_out_1_port, B(0) => 
                           LMD_out_0_port, C(31) => link_addr_W_31_port, C(30) 
                           => link_addr_W_30_port, C(29) => link_addr_W_29_port
                           , C(28) => link_addr_W_28_port, C(27) => 
                           link_addr_W_27_port, C(26) => link_addr_W_26_port, 
                           C(25) => link_addr_W_25_port, C(24) => 
                           link_addr_W_24_port, C(23) => link_addr_W_23_port, 
                           C(22) => link_addr_W_22_port, C(21) => 
                           link_addr_W_21_port, C(20) => link_addr_W_20_port, 
                           C(19) => link_addr_W_19_port, C(18) => 
                           link_addr_W_18_port, C(17) => link_addr_W_17_port, 
                           C(16) => link_addr_W_16_port, C(15) => 
                           link_addr_W_15_port, C(14) => link_addr_W_14_port, 
                           C(13) => link_addr_W_13_port, C(12) => 
                           link_addr_W_12_port, C(11) => link_addr_W_11_port, 
                           C(10) => link_addr_W_10_port, C(9) => 
                           link_addr_W_9_port, C(8) => link_addr_W_8_port, C(7)
                           => link_addr_W_7_port, C(6) => link_addr_W_6_port, 
                           C(5) => link_addr_W_5_port, C(4) => 
                           link_addr_W_4_port, C(3) => link_addr_W_3_port, C(2)
                           => link_addr_W_2_port, C(1) => link_addr_W_1_port, 
                           C(0) => link_addr_W_0_port, SEL(1) => WB_MUX_SEL(1),
                           SEL(0) => WB_MUX_SEL(0), Y(31) => WB_31_port, Y(30) 
                           => WB_30_port, Y(29) => WB_29_port, Y(28) => 
                           WB_28_port, Y(27) => WB_27_port, Y(26) => WB_26_port
                           , Y(25) => WB_25_port, Y(24) => WB_24_port, Y(23) =>
                           WB_23_port, Y(22) => WB_22_port, Y(21) => WB_21_port
                           , Y(20) => WB_20_port, Y(19) => WB_19_port, Y(18) =>
                           WB_18_port, Y(17) => WB_17_port, Y(16) => WB_16_port
                           , Y(15) => WB_15_port, Y(14) => WB_14_port, Y(13) =>
                           WB_13_port, Y(12) => WB_12_port, Y(11) => WB_11_port
                           , Y(10) => WB_10_port, Y(9) => WB_9_port, Y(8) => 
                           WB_8_port, Y(7) => WB_7_port, Y(6) => WB_6_port, 
                           Y(5) => WB_5_port, Y(4) => WB_4_port, Y(3) => 
                           WB_3_port, Y(2) => WB_2_port, Y(1) => WB_1_port, 
                           Y(0) => WB_0_port);
   U2 : CLKBUF_X1 port map( A => alu_out_29_port, Z => n1);
   U3 : CLKBUF_X1 port map( A => ALU_OPCODE(3), Z => n2);
   U4 : CLKBUF_X1 port map( A => opcode_E_3_port, Z => n3);
   U5 : CLKBUF_X1 port map( A => opcode_W_2_port, Z => n4);
   U6 : CLKBUF_X1 port map( A => opcode_M_2_port, Z => n5);
   U7 : CLKBUF_X1 port map( A => opcode_W_3_port, Z => n6);
   U8 : CLKBUF_X1 port map( A => opcode_E_0_port, Z => n7);
   U9 : CLKBUF_X1 port map( A => opcode_M_4_port, Z => n8);
   U10 : CLKBUF_X1 port map( A => opcode_E_4_port, Z => n9);
   U11 : BUF_X1 port map( A => Rst, Z => n16);
   U12 : CLKBUF_X1 port map( A => opcode_M_0_port, Z => n10);
   U13 : CLKBUF_X1 port map( A => opcode_W_4_port, Z => n11);
   U14 : CLKBUF_X1 port map( A => opcode_W_1_port, Z => n12);
   U15 : CLKBUF_X1 port map( A => opcode_E_1_port, Z => n13);
   U16 : CLKBUF_X1 port map( A => opcode_M_1_port, Z => n14);
   U17 : CLKBUF_X1 port map( A => opcode_M_3_port, Z => n15);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11 is

   port( Clk, Rst : in std_logic;  OPCODE_IN : in std_logic_vector (5 downto 0)
         ;  FUNC_IN : in std_logic_vector (10 downto 0);  MUXA_SEL, MUXB_SEL, 
         BR_EN : out std_logic;  ALU_OPCODE : out std_logic_vector (0 to 4);  
         DRAM_RW, DRAM_EN : out std_logic;  DRAM_SEL : out std_logic_vector (2 
         downto 0);  WB_MUX_SEL : out std_logic_vector (1 downto 0);  RF_WE : 
         out std_logic);

end dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal cw_10_port, cw_9_port, cw_8_port, cw_5_port, cw_4_port, cw_3_port, 
      cw_1_port, cw_0_port, cw1_7_port, cw1_6_port, cw1_5_port, cw1_4_port, 
      cw1_3_port, cw1_2_port, cw1_1_port, cw1_0_port, cw2_2_port, cw2_1_port, 
      cw2_0_port, aluOpcode_i_4_port, aluOpcode_i_3_port, aluOpcode_i_2_port, 
      aluOpcode_i_1_port, aluOpcode_i_0_port, n1, n38, n39, n40, n41, n42, n43,
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n138, n139, n140, n141, n_1756, n_1757, n_1758
      , n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767,
      n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, 
      n_1777, n_1778, n_1779, n_1780, n_1781, n_1782 : std_logic;

begin
   
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => aluOpcode_i_4_port, CK => Clk
                           , RN => n4, Q => ALU_OPCODE(0), QN => n_1756);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => n6, Q => ALU_OPCODE(1), QN => n_1757);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => n6, Q => ALU_OPCODE(2), QN => n_1758);
   cw1_reg_10_inst : DFFR_X1 port map( D => cw_10_port, CK => Clk, RN => n5, Q 
                           => MUXA_SEL, QN => n_1759);
   cw1_reg_9_inst : DFFR_X1 port map( D => cw_9_port, CK => Clk, RN => n5, Q =>
                           MUXB_SEL, QN => n_1760);
   cw1_reg_8_inst : DFFR_X1 port map( D => cw_8_port, CK => Clk, RN => n5, Q =>
                           BR_EN, QN => n_1761);
   cw1_reg_7_inst : SDFFR_X1 port map( D => n110, SI => n1, SE => n47, CK => 
                           Clk, RN => n6, Q => cw1_7_port, QN => n_1762);
   cw1_reg_6_inst : DFFR_X1 port map( D => n12, CK => Clk, RN => n5, Q => 
                           cw1_6_port, QN => n_1763);
   cw1_reg_5_inst : DFFR_X1 port map( D => cw_5_port, CK => Clk, RN => n5, Q =>
                           cw1_5_port, QN => n_1764);
   cw1_reg_4_inst : DFFR_X1 port map( D => cw_4_port, CK => Clk, RN => n5, Q =>
                           cw1_4_port, QN => n_1765);
   cw1_reg_3_inst : DFFR_X1 port map( D => cw_3_port, CK => Clk, RN => n5, Q =>
                           cw1_3_port, QN => n_1766);
   cw1_reg_2_inst : DFFR_X1 port map( D => n11, CK => Clk, RN => n5, Q => 
                           cw1_2_port, QN => n_1767);
   cw1_reg_1_inst : DFFR_X1 port map( D => cw_1_port, CK => Clk, RN => n5, Q =>
                           cw1_1_port, QN => n_1768);
   cw1_reg_0_inst : DFFR_X1 port map( D => cw_0_port, CK => Clk, RN => n4, Q =>
                           cw1_0_port, QN => n_1769);
   cw2_reg_7_inst : DFFR_X1 port map( D => cw1_7_port, CK => Clk, RN => n4, Q 
                           => DRAM_RW, QN => n_1770);
   cw2_reg_6_inst : DFFR_X1 port map( D => cw1_6_port, CK => Clk, RN => n4, Q 
                           => DRAM_EN, QN => n_1771);
   cw2_reg_5_inst : DFFR_X1 port map( D => cw1_5_port, CK => Clk, RN => n4, Q 
                           => DRAM_SEL(2), QN => n_1772);
   cw2_reg_4_inst : DFFR_X1 port map( D => cw1_4_port, CK => Clk, RN => n4, Q 
                           => DRAM_SEL(1), QN => n_1773);
   cw2_reg_3_inst : DFFR_X1 port map( D => cw1_3_port, CK => Clk, RN => n4, Q 
                           => DRAM_SEL(0), QN => n_1774);
   cw2_reg_2_inst : DFFR_X1 port map( D => cw1_2_port, CK => Clk, RN => n4, Q 
                           => cw2_2_port, QN => n_1775);
   cw2_reg_1_inst : DFFR_X1 port map( D => cw1_1_port, CK => Clk, RN => n4, Q 
                           => cw2_1_port, QN => n_1776);
   cw2_reg_0_inst : DFFR_X1 port map( D => cw1_0_port, CK => Clk, RN => n4, Q 
                           => cw2_0_port, QN => n_1777);
   cw3_reg_2_inst : DFFR_X1 port map( D => cw2_2_port, CK => Clk, RN => n4, Q 
                           => WB_MUX_SEL(1), QN => n_1778);
   cw3_reg_1_inst : DFFR_X1 port map( D => cw2_1_port, CK => Clk, RN => n4, Q 
                           => WB_MUX_SEL(0), QN => n_1779);
   cw3_reg_0_inst : DFFR_X1 port map( D => cw2_0_port, CK => Clk, RN => n5, Q 
                           => RF_WE, QN => n_1780);
   n1 <= '0';
   U132 : NAND3_X1 port map( A1 => n52, A2 => n28, A3 => n30, ZN => n49);
   U133 : XOR2_X1 port map( A => n31, B => OPCODE_IN(2), Z => n42);
   U134 : OAI33_X1 port map( A1 => n45, A2 => n3, A3 => OPCODE_IN(2), B1 => n62
                           , B2 => n31, B3 => n24, ZN => n61);
   U135 : NAND3_X1 port map( A1 => OPCODE_IN(2), A2 => n3, A3 => n30, ZN => n64
                           );
   U136 : NAND3_X1 port map( A1 => n31, A2 => n27, A3 => n52, ZN => n58);
   U137 : NAND3_X1 port map( A1 => n91, A2 => n140, A3 => n16, ZN => n80);
   U138 : NAND3_X1 port map( A1 => n103, A2 => n33, A3 => n19, ZN => n102);
   U139 : OAI33_X1 port map( A1 => n92, A2 => FUNC_IN(1), A3 => n104, B1 => 
                           n105, B2 => n106, B3 => n37, ZN => n96);
   U140 : NAND3_X1 port map( A1 => n30, A2 => n20, A3 => n25, ZN => n88);
   U141 : NAND3_X1 port map( A1 => n77, A2 => n141, A3 => n15, ZN => n113);
   U142 : NAND3_X1 port map( A1 => n101, A2 => n100, A3 => n127, ZN => n126);
   U143 : NAND3_X1 port map( A1 => n15, A2 => FUNC_IN(4), A3 => n78, ZN => n127
                           );
   U144 : NAND3_X1 port map( A1 => n128, A2 => n22, A3 => n32, ZN => n100);
   U145 : NAND3_X1 port map( A1 => n26, A2 => n30, A3 => n19, ZN => n101);
   U146 : NAND3_X1 port map( A1 => OPCODE_IN(2), A2 => n3, A3 => OPCODE_IN(3), 
                           ZN => n121);
   U147 : NAND3_X1 port map( A1 => n3, A2 => n20, A3 => n103, ZN => n73);
   U148 : NAND3_X1 port map( A1 => n3, A2 => n20, A3 => n128, ZN => n72);
   U149 : NAND3_X1 port map( A1 => n128, A2 => n22, A3 => n33, ZN => n66);
   U150 : NAND3_X1 port map( A1 => n3, A2 => n20, A3 => n26, ZN => n90);
   U151 : NAND3_X1 port map( A1 => n17, A2 => n141, A3 => n109, ZN => n112);
   U152 : OAI33_X1 port map( A1 => n141, A2 => n108, A3 => n139, B1 => n86, B2 
                           => FUNC_IN(3), B3 => FUNC_IN(2), ZN => n135);
   U153 : NAND3_X1 port map( A1 => OPCODE_IN(3), A2 => OPCODE_IN(2), A3 => n19,
                           ZN => n111);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => n5, Q => ALU_OPCODE(4), QN => n_1781);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => n5, Q => ALU_OPCODE(3), QN => n_1782);
   U4 : OR2_X1 port map( A1 => n47, A2 => n32, ZN => n2);
   U5 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n74);
   U6 : OAI21_X1 port map( B1 => n45, B2 => n72, A => n100, ZN => n70);
   U7 : INV_X1 port map( A => n57, ZN => n19);
   U8 : INV_X1 port map( A => n72, ZN => n9);
   U9 : INV_X1 port map( A => n45, ZN => n30);
   U10 : OAI21_X1 port map( B1 => n45, B2 => n46, A => n2, ZN => cw_5_port);
   U11 : NAND2_X1 port map( A1 => n26, A2 => n52, ZN => n46);
   U12 : OR4_X1 port map( A1 => n98, A2 => n99, A3 => n89, A4 => n70, ZN => n97
                           );
   U13 : AND3_X1 port map( A1 => n120, A2 => n46, A3 => n130, ZN => n129);
   U14 : INV_X1 port map( A => n56, ZN => n23);
   U15 : INV_X1 port map( A => n90, ZN => n7);
   U16 : AND2_X1 port map( A1 => n51, A2 => n47, ZN => n130);
   U17 : INV_X1 port map( A => n88, ZN => n10);
   U18 : NOR2_X1 port map( A1 => n20, A2 => n3, ZN => n52);
   U19 : NOR4_X1 port map( A1 => n28, A2 => n60, A3 => n27, A4 => n48, ZN => 
                           n75);
   U20 : NOR3_X1 port map( A1 => n48, A2 => n62, A3 => n57, ZN => n84);
   U21 : OAI221_X1 port map( B1 => n112, B2 => n116, C1 => n45, C2 => n90, A =>
                           n117, ZN => n98);
   U22 : NAND2_X1 port map( A1 => n37, A2 => n35, ZN => n116);
   U23 : NOR2_X1 port map( A1 => n21, A2 => n84, ZN => n117);
   U24 : INV_X1 port map( A => n65, ZN => n21);
   U25 : OAI221_X1 port map( B1 => n86, B2 => n87, C1 => n74, C2 => n90, A => 
                           n66, ZN => n99);
   U26 : NOR3_X1 port map( A1 => n60, A2 => n42, A3 => n27, ZN => n56);
   U27 : NAND4_X1 port map( A1 => n113, A2 => n88, A3 => n18, A4 => n114, ZN =>
                           aluOpcode_i_1_port);
   U28 : INV_X1 port map( A => n118, ZN => n18);
   U29 : AOI211_X1 port map( C1 => n32, C2 => n9, A => n115, B => n98, ZN => 
                           n114);
   U30 : NAND2_X1 port map( A1 => n31, A2 => n34, ZN => n45);
   U31 : OAI211_X1 port map( C1 => n45, C2 => n111, A => n8, B => n132, ZN => 
                           n115);
   U32 : INV_X1 port map( A => n99, ZN => n8);
   U33 : AOI221_X1 port map( B1 => n9, B2 => n33, C1 => n133, C2 => n78, A => 
                           n83, ZN => n132);
   U34 : NOR2_X1 port map( A1 => n105, A2 => n141, ZN => n133);
   U35 : INV_X1 port map( A => n110, ZN => n32);
   U36 : NOR3_X1 port map( A1 => n141, A2 => n86, A3 => n87, ZN => n85);
   U37 : INV_X1 port map( A => n50, ZN => n33);
   U38 : NAND2_X1 port map( A1 => n128, A2 => n52, ZN => n47);
   U39 : NAND2_X1 port map( A1 => n20, A2 => n24, ZN => n57);
   U40 : NAND2_X1 port map( A1 => n103, A2 => n52, ZN => n51);
   U41 : INV_X1 port map( A => n3, ZN => n24);
   U42 : OAI211_X1 port map( C1 => n34, C2 => n51, A => n58, B => n53, ZN => 
                           cw_0_port);
   U43 : INV_X1 port map( A => n121, ZN => n25);
   U44 : INV_X1 port map( A => n62, ZN => n26);
   U45 : INV_X1 port map( A => n86, ZN => n17);
   U46 : NAND2_X1 port map( A1 => n19, A2 => n128, ZN => n120);
   U47 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           aluOpcode_i_4_port);
   U48 : AOI211_X1 port map( C1 => n36, C2 => n69, A => n70, B => n71, ZN => 
                           n68);
   U49 : AOI21_X1 port map( B1 => n15, B2 => n138, A => n75, ZN => n67);
   U50 : AOI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n71);
   U51 : INV_X1 port map( A => n111, ZN => n13);
   U52 : AND3_X1 port map( A1 => n19, A2 => n103, A3 => n32, ZN => n83);
   U53 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           aluOpcode_i_3_port);
   U54 : OAI21_X1 port map( B1 => n25, B2 => n9, A => n29, ZN => n79);
   U55 : AOI21_X1 port map( B1 => n7, B2 => n33, A => n89, ZN => n81);
   U56 : NOR4_X1 port map( A1 => n10, A2 => n83, A3 => n84, A4 => n85, ZN => 
                           n82);
   U57 : INV_X1 port map( A => n60, ZN => n22);
   U58 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => n89);
   U59 : INV_X1 port map( A => n105, ZN => n15);
   U60 : NAND2_X1 port map( A1 => n122, A2 => n123, ZN => aluOpcode_i_0_port);
   U61 : AOI221_X1 port map( B1 => n33, B2 => n124, C1 => n29, C2 => n125, A =>
                           n126, ZN => n123);
   U62 : AOI211_X1 port map( C1 => n13, C2 => n32, A => n131, B => n115, ZN => 
                           n122);
   U63 : NAND2_X1 port map( A1 => n130, A2 => n73, ZN => n124);
   U64 : INV_X1 port map( A => n108, ZN => n16);
   U65 : OAI22_X1 port map( A1 => n119, A2 => n92, B1 => n120, B2 => n74, ZN =>
                           n118);
   U66 : OR2_X1 port map( A1 => n106, A2 => n86, ZN => n119);
   U67 : INV_X1 port map( A => n39, ZN => n12);
   U68 : INV_X1 port map( A => n53, ZN => n11);
   U69 : AOI21_X1 port map( B1 => n141, B2 => n77, A => n78, ZN => n106);
   U70 : INV_X1 port map( A => n48, ZN => n29);
   U71 : INV_X1 port map( A => n92, ZN => n36);
   U72 : NOR2_X1 port map( A1 => OPCODE_IN(2), A2 => OPCODE_IN(3), ZN => n103);
   U73 : NOR2_X1 port map( A1 => n27, A2 => OPCODE_IN(2), ZN => n128);
   U74 : NOR3_X1 port map( A1 => FUNC_IN(0), A2 => FUNC_IN(2), A3 => n108, ZN 
                           => n69);
   U75 : NAND2_X1 port map( A1 => OPCODE_IN(2), A2 => n27, ZN => n62);
   U76 : NAND4_X1 port map( A1 => n19, A2 => n103, A3 => n136, A4 => n137, ZN 
                           => n86);
   U77 : NOR4_X1 port map( A1 => FUNC_IN(9), A2 => FUNC_IN(8), A3 => FUNC_IN(7)
                           , A4 => FUNC_IN(6), ZN => n137);
   U78 : NOR2_X1 port map( A1 => FUNC_IN(10), A2 => n45, ZN => n136);
   U79 : INV_X1 port map( A => OPCODE_IN(1), ZN => n31);
   U80 : INV_X1 port map( A => OPCODE_IN(2), ZN => n28);
   U81 : NOR3_X1 port map( A1 => n43, A2 => OPCODE_IN(5), A3 => OPCODE_IN(3), 
                           ZN => cw_8_port);
   U82 : AOI22_X1 port map( A1 => n44, A2 => OPCODE_IN(2), B1 => OPCODE_IN(1), 
                           B2 => n28, ZN => n43);
   U83 : NOR2_X1 port map( A1 => n3, A2 => OPCODE_IN(1), ZN => n44);
   U84 : INV_X1 port map( A => OPCODE_IN(3), ZN => n27);
   U85 : AOI21_X1 port map( B1 => n20, B2 => n59, A => n56, ZN => n53);
   U86 : OAI21_X1 port map( B1 => n50, B2 => OPCODE_IN(2), A => n54, ZN => n59)
                           ;
   U87 : NAND4_X1 port map( A1 => n30, A2 => OPCODE_IN(3), A3 => n22, A4 => 
                           OPCODE_IN(2), ZN => n65);
   U88 : NAND2_X1 port map( A1 => OPCODE_IN(1), A2 => n34, ZN => n110);
   U89 : OAI221_X1 port map( B1 => n47, B2 => n50, C1 => OPCODE_IN(1), C2 => 
                           n51, A => n49, ZN => cw_3_port);
   U90 : OAI221_X1 port map( B1 => n46, B2 => n48, C1 => OPCODE_IN(1), C2 => 
                           n47, A => n49, ZN => cw_4_port);
   U91 : NAND2_X1 port map( A1 => OPCODE_IN(0), A2 => n31, ZN => n48);
   U92 : INV_X1 port map( A => OPCODE_IN(5), ZN => n20);
   U93 : OAI22_X1 port map( A1 => n129, A2 => n45, B1 => n134, B2 => n92, ZN =>
                           n131);
   U94 : AOI21_X1 port map( B1 => n135, B2 => n140, A => n14, ZN => n134);
   U95 : INV_X1 port map( A => n112, ZN => n14);
   U96 : OAI21_X1 port map( B1 => n63, B2 => n27, A => n64, ZN => n41);
   U97 : AOI211_X1 port map( C1 => n34, C2 => n24, A => n28, B => n31, ZN => 
                           n63);
   U98 : NAND2_X1 port map( A1 => OPCODE_IN(0), A2 => OPCODE_IN(1), ZN => n50);
   U99 : OAI211_X1 port map( C1 => OPCODE_IN(5), C2 => n54, A => n23, B => n39,
                           ZN => cw_1_port);
   U100 : OAI211_X1 port map( C1 => OPCODE_IN(5), C2 => n38, A => n23, B => n39
                           , ZN => cw_9_port);
   U101 : AOI21_X1 port map( B1 => n40, B2 => n27, A => n41, ZN => n38);
   U102 : OAI22_X1 port map( A1 => n31, A2 => n24, B1 => n3, B2 => n42, ZN => 
                           n40);
   U103 : OAI21_X1 port map( B1 => OPCODE_IN(5), B2 => n121, A => n129, ZN => 
                           n125);
   U104 : NOR2_X1 port map( A1 => n41, A2 => n61, ZN => n54);
   U105 : NAND2_X1 port map( A1 => n3, A2 => OPCODE_IN(5), ZN => n60);
   U106 : NOR3_X1 port map( A1 => n57, A2 => OPCODE_IN(3), A3 => n42, ZN => 
                           cw_10_port);
   U107 : INV_X1 port map( A => OPCODE_IN(0), ZN => n34);
   U108 : NAND2_X1 port map( A1 => n52, A2 => n55, ZN => n39);
   U109 : OAI22_X1 port map( A1 => OPCODE_IN(3), A2 => OPCODE_IN(1), B1 => 
                           OPCODE_IN(2), B2 => n32, ZN => n55);
   U110 : NAND2_X1 port map( A1 => FUNC_IN(5), A2 => n16, ZN => n105);
   U111 : OAI22_X1 port map( A1 => n92, A2 => n141, B1 => n93, B2 => n139, ZN 
                           => n91);
   U112 : AOI21_X1 port map( B1 => FUNC_IN(0), B2 => FUNC_IN(5), A => n36, ZN 
                           => n93);
   U113 : NAND2_X1 port map( A1 => FUNC_IN(3), A2 => n17, ZN => n108);
   U114 : OR4_X1 port map( A1 => n94, A2 => n95, A3 => n96, A4 => n97, ZN => 
                           aluOpcode_i_2_port);
   U115 : AOI21_X1 port map( B1 => n110, B2 => n48, A => n111, ZN => n95);
   U116 : NOR3_X1 port map( A1 => n112, A2 => FUNC_IN(4), A3 => n140, ZN => n94
                           );
   U117 : NOR2_X1 port map( A1 => n107, A2 => n69, ZN => n104);
   U118 : AND3_X1 port map( A1 => FUNC_IN(0), A2 => n17, A3 => n109, ZN => n107
                           );
   U119 : BUF_X1 port map( A => OPCODE_IN(4), Z => n3);
   U120 : NOR2_X1 port map( A1 => n140, A2 => FUNC_IN(2), ZN => n78);
   U121 : NOR2_X1 port map( A1 => n139, A2 => FUNC_IN(1), ZN => n77);
   U122 : INV_X1 port map( A => FUNC_IN(0), ZN => n141);
   U123 : NAND4_X1 port map( A1 => n109, A2 => FUNC_IN(1), A3 => n37, A4 => n35
                           , ZN => n87);
   U124 : NOR2_X1 port map( A1 => n139, A2 => FUNC_IN(3), ZN => n109);
   U125 : NAND2_X1 port map( A1 => FUNC_IN(5), A2 => n37, ZN => n92);
   U126 : INV_X1 port map( A => n76, ZN => n138);
   U127 : AOI21_X1 port map( B1 => n77, B2 => FUNC_IN(4), A => n78, ZN => n76);
   U128 : INV_X1 port map( A => FUNC_IN(1), ZN => n140);
   U129 : INV_X1 port map( A => FUNC_IN(4), ZN => n37);
   U130 : INV_X1 port map( A => FUNC_IN(2), ZN => n139);
   U131 : INV_X1 port map( A => FUNC_IN(5), ZN => n35);
   U154 : BUF_X1 port map( A => Rst, Z => n5);
   U155 : BUF_X1 port map( A => Rst, Z => n4);
   U156 : BUF_X1 port map( A => Rst, Z => n6);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity DLX_syn is

   port( Clk, Rst : in std_logic;  IRAM_DATA_OUT, DRAM_DATA_OUT : in 
         std_logic_vector (31 downto 0);  DRAM_DATA_IN : out std_logic_vector 
         (31 downto 0);  DRAM_ADDRESS : out std_logic_vector (11 downto 0);  
         DRAM_ENABLE, DRAM_RW : out std_logic;  DRAM_SEL : out std_logic_vector
         (2 downto 0);  IRAM_ADDRESS : out std_logic_vector (7 downto 0));

end DLX_syn;

architecture SYN_structural of DLX_syn is

   component DPATH
      port( Clk, Rst, MUXA_SEL, MUXB_SEL, BR_EN : in std_logic;  ALU_OPCODE : 
            in std_logic_vector (0 to 4);  WB_MUX_SEL : in std_logic_vector (1 
            downto 0);  RF_WE : in std_logic;  DRAM_OUT, IRAM_OUT : in 
            std_logic_vector (31 downto 0);  IR1, DRAM_IN : out 
            std_logic_vector (31 downto 0);  DRAM_ADD : out std_logic_vector 
            (11 downto 0);  IR_ADD : out std_logic_vector (7 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11
      port( Clk, Rst : in std_logic;  OPCODE_IN : in std_logic_vector (5 downto
            0);  FUNC_IN : in std_logic_vector (10 downto 0);  MUXA_SEL, 
            MUXB_SEL, BR_EN : out std_logic;  ALU_OPCODE : out std_logic_vector
            (0 to 4);  DRAM_RW, DRAM_EN : out std_logic;  DRAM_SEL : out 
            std_logic_vector (2 downto 0);  WB_MUX_SEL : out std_logic_vector 
            (1 downto 0);  RF_WE : out std_logic);
   end component;
   
   signal IR_CU_31, IR_CU_30, IR_CU_29, IR_CU_28, IR_CU_27, IR_CU_26, 
      IR_CU_10_port, IR_CU_9_port, IR_CU_8_port, IR_CU_7_port, IR_CU_6_port, 
      IR_CU_5_port, IR_CU_4_port, IR_CU_3_port, IR_CU_2_port, IR_CU_1_port, 
      IR_CU_0_port, MUXA_SEL_i, MUXB_SEL_i, BR_EN_i, ALU_OPCODE_i_4_port, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, 
      ALU_OPCODE_i_0_port, WB_MUX_SEL_i_1_port, WB_MUX_SEL_i_0_port, RF_WE_i, 
      n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, 
      n_1792, n_1793, n_1794, n_1795, n_1796, n_1797 : std_logic;

begin
   
   CU_I : 
                           dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11 
                           port map( Clk => Clk, Rst => Rst, OPCODE_IN(5) => 
                           IR_CU_31, OPCODE_IN(4) => IR_CU_30, OPCODE_IN(3) => 
                           IR_CU_29, OPCODE_IN(2) => IR_CU_28, OPCODE_IN(1) => 
                           IR_CU_27, OPCODE_IN(0) => IR_CU_26, FUNC_IN(10) => 
                           IR_CU_10_port, FUNC_IN(9) => IR_CU_9_port, 
                           FUNC_IN(8) => IR_CU_8_port, FUNC_IN(7) => 
                           IR_CU_7_port, FUNC_IN(6) => IR_CU_6_port, FUNC_IN(5)
                           => IR_CU_5_port, FUNC_IN(4) => IR_CU_4_port, 
                           FUNC_IN(3) => IR_CU_3_port, FUNC_IN(2) => 
                           IR_CU_2_port, FUNC_IN(1) => IR_CU_1_port, FUNC_IN(0)
                           => IR_CU_0_port, MUXA_SEL => MUXA_SEL_i, MUXB_SEL =>
                           MUXB_SEL_i, BR_EN => BR_EN_i, ALU_OPCODE(0) => 
                           ALU_OPCODE_i_4_port, ALU_OPCODE(1) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_0_port, DRAM_RW => DRAM_RW, DRAM_EN => 
                           DRAM_ENABLE, DRAM_SEL(2) => DRAM_SEL(2), DRAM_SEL(1)
                           => DRAM_SEL(1), DRAM_SEL(0) => DRAM_SEL(0), 
                           WB_MUX_SEL(1) => WB_MUX_SEL_i_1_port, WB_MUX_SEL(0) 
                           => WB_MUX_SEL_i_0_port, RF_WE => RF_WE_i);
   DataP : DPATH port map( Clk => Clk, Rst => Rst, MUXA_SEL => MUXA_SEL_i, 
                           MUXB_SEL => MUXB_SEL_i, BR_EN => BR_EN_i, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_4_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_3_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_0_port, WB_MUX_SEL(1) => 
                           WB_MUX_SEL_i_1_port, WB_MUX_SEL(0) => 
                           WB_MUX_SEL_i_0_port, RF_WE => RF_WE_i, DRAM_OUT(31) 
                           => DRAM_DATA_OUT(31), DRAM_OUT(30) => 
                           DRAM_DATA_OUT(30), DRAM_OUT(29) => DRAM_DATA_OUT(29)
                           , DRAM_OUT(28) => DRAM_DATA_OUT(28), DRAM_OUT(27) =>
                           DRAM_DATA_OUT(27), DRAM_OUT(26) => DRAM_DATA_OUT(26)
                           , DRAM_OUT(25) => DRAM_DATA_OUT(25), DRAM_OUT(24) =>
                           DRAM_DATA_OUT(24), DRAM_OUT(23) => DRAM_DATA_OUT(23)
                           , DRAM_OUT(22) => DRAM_DATA_OUT(22), DRAM_OUT(21) =>
                           DRAM_DATA_OUT(21), DRAM_OUT(20) => DRAM_DATA_OUT(20)
                           , DRAM_OUT(19) => DRAM_DATA_OUT(19), DRAM_OUT(18) =>
                           DRAM_DATA_OUT(18), DRAM_OUT(17) => DRAM_DATA_OUT(17)
                           , DRAM_OUT(16) => DRAM_DATA_OUT(16), DRAM_OUT(15) =>
                           DRAM_DATA_OUT(15), DRAM_OUT(14) => DRAM_DATA_OUT(14)
                           , DRAM_OUT(13) => DRAM_DATA_OUT(13), DRAM_OUT(12) =>
                           DRAM_DATA_OUT(12), DRAM_OUT(11) => DRAM_DATA_OUT(11)
                           , DRAM_OUT(10) => DRAM_DATA_OUT(10), DRAM_OUT(9) => 
                           DRAM_DATA_OUT(9), DRAM_OUT(8) => DRAM_DATA_OUT(8), 
                           DRAM_OUT(7) => DRAM_DATA_OUT(7), DRAM_OUT(6) => 
                           DRAM_DATA_OUT(6), DRAM_OUT(5) => DRAM_DATA_OUT(5), 
                           DRAM_OUT(4) => DRAM_DATA_OUT(4), DRAM_OUT(3) => 
                           DRAM_DATA_OUT(3), DRAM_OUT(2) => DRAM_DATA_OUT(2), 
                           DRAM_OUT(1) => DRAM_DATA_OUT(1), DRAM_OUT(0) => 
                           DRAM_DATA_OUT(0), IRAM_OUT(31) => IRAM_DATA_OUT(31),
                           IRAM_OUT(30) => IRAM_DATA_OUT(30), IRAM_OUT(29) => 
                           IRAM_DATA_OUT(29), IRAM_OUT(28) => IRAM_DATA_OUT(28)
                           , IRAM_OUT(27) => IRAM_DATA_OUT(27), IRAM_OUT(26) =>
                           IRAM_DATA_OUT(26), IRAM_OUT(25) => IRAM_DATA_OUT(25)
                           , IRAM_OUT(24) => IRAM_DATA_OUT(24), IRAM_OUT(23) =>
                           IRAM_DATA_OUT(23), IRAM_OUT(22) => IRAM_DATA_OUT(22)
                           , IRAM_OUT(21) => IRAM_DATA_OUT(21), IRAM_OUT(20) =>
                           IRAM_DATA_OUT(20), IRAM_OUT(19) => IRAM_DATA_OUT(19)
                           , IRAM_OUT(18) => IRAM_DATA_OUT(18), IRAM_OUT(17) =>
                           IRAM_DATA_OUT(17), IRAM_OUT(16) => IRAM_DATA_OUT(16)
                           , IRAM_OUT(15) => IRAM_DATA_OUT(15), IRAM_OUT(14) =>
                           IRAM_DATA_OUT(14), IRAM_OUT(13) => IRAM_DATA_OUT(13)
                           , IRAM_OUT(12) => IRAM_DATA_OUT(12), IRAM_OUT(11) =>
                           IRAM_DATA_OUT(11), IRAM_OUT(10) => IRAM_DATA_OUT(10)
                           , IRAM_OUT(9) => IRAM_DATA_OUT(9), IRAM_OUT(8) => 
                           IRAM_DATA_OUT(8), IRAM_OUT(7) => IRAM_DATA_OUT(7), 
                           IRAM_OUT(6) => IRAM_DATA_OUT(6), IRAM_OUT(5) => 
                           IRAM_DATA_OUT(5), IRAM_OUT(4) => IRAM_DATA_OUT(4), 
                           IRAM_OUT(3) => IRAM_DATA_OUT(3), IRAM_OUT(2) => 
                           IRAM_DATA_OUT(2), IRAM_OUT(1) => IRAM_DATA_OUT(1), 
                           IRAM_OUT(0) => IRAM_DATA_OUT(0), IR1(31) => IR_CU_31
                           , IR1(30) => IR_CU_30, IR1(29) => IR_CU_29, IR1(28) 
                           => IR_CU_28, IR1(27) => IR_CU_27, IR1(26) => 
                           IR_CU_26, IR1(25) => n_1783, IR1(24) => n_1784, 
                           IR1(23) => n_1785, IR1(22) => n_1786, IR1(21) => 
                           n_1787, IR1(20) => n_1788, IR1(19) => n_1789, 
                           IR1(18) => n_1790, IR1(17) => n_1791, IR1(16) => 
                           n_1792, IR1(15) => n_1793, IR1(14) => n_1794, 
                           IR1(13) => n_1795, IR1(12) => n_1796, IR1(11) => 
                           n_1797, IR1(10) => IR_CU_10_port, IR1(9) => 
                           IR_CU_9_port, IR1(8) => IR_CU_8_port, IR1(7) => 
                           IR_CU_7_port, IR1(6) => IR_CU_6_port, IR1(5) => 
                           IR_CU_5_port, IR1(4) => IR_CU_4_port, IR1(3) => 
                           IR_CU_3_port, IR1(2) => IR_CU_2_port, IR1(1) => 
                           IR_CU_1_port, IR1(0) => IR_CU_0_port, DRAM_IN(31) =>
                           DRAM_DATA_IN(31), DRAM_IN(30) => DRAM_DATA_IN(30), 
                           DRAM_IN(29) => DRAM_DATA_IN(29), DRAM_IN(28) => 
                           DRAM_DATA_IN(28), DRAM_IN(27) => DRAM_DATA_IN(27), 
                           DRAM_IN(26) => DRAM_DATA_IN(26), DRAM_IN(25) => 
                           DRAM_DATA_IN(25), DRAM_IN(24) => DRAM_DATA_IN(24), 
                           DRAM_IN(23) => DRAM_DATA_IN(23), DRAM_IN(22) => 
                           DRAM_DATA_IN(22), DRAM_IN(21) => DRAM_DATA_IN(21), 
                           DRAM_IN(20) => DRAM_DATA_IN(20), DRAM_IN(19) => 
                           DRAM_DATA_IN(19), DRAM_IN(18) => DRAM_DATA_IN(18), 
                           DRAM_IN(17) => DRAM_DATA_IN(17), DRAM_IN(16) => 
                           DRAM_DATA_IN(16), DRAM_IN(15) => DRAM_DATA_IN(15), 
                           DRAM_IN(14) => DRAM_DATA_IN(14), DRAM_IN(13) => 
                           DRAM_DATA_IN(13), DRAM_IN(12) => DRAM_DATA_IN(12), 
                           DRAM_IN(11) => DRAM_DATA_IN(11), DRAM_IN(10) => 
                           DRAM_DATA_IN(10), DRAM_IN(9) => DRAM_DATA_IN(9), 
                           DRAM_IN(8) => DRAM_DATA_IN(8), DRAM_IN(7) => 
                           DRAM_DATA_IN(7), DRAM_IN(6) => DRAM_DATA_IN(6), 
                           DRAM_IN(5) => DRAM_DATA_IN(5), DRAM_IN(4) => 
                           DRAM_DATA_IN(4), DRAM_IN(3) => DRAM_DATA_IN(3), 
                           DRAM_IN(2) => DRAM_DATA_IN(2), DRAM_IN(1) => 
                           DRAM_DATA_IN(1), DRAM_IN(0) => DRAM_DATA_IN(0), 
                           DRAM_ADD(11) => DRAM_ADDRESS(11), DRAM_ADD(10) => 
                           DRAM_ADDRESS(10), DRAM_ADD(9) => DRAM_ADDRESS(9), 
                           DRAM_ADD(8) => DRAM_ADDRESS(8), DRAM_ADD(7) => 
                           DRAM_ADDRESS(7), DRAM_ADD(6) => DRAM_ADDRESS(6), 
                           DRAM_ADD(5) => DRAM_ADDRESS(5), DRAM_ADD(4) => 
                           DRAM_ADDRESS(4), DRAM_ADD(3) => DRAM_ADDRESS(3), 
                           DRAM_ADD(2) => DRAM_ADDRESS(2), DRAM_ADD(1) => 
                           DRAM_ADDRESS(1), DRAM_ADD(0) => DRAM_ADDRESS(0), 
                           IR_ADD(7) => IRAM_ADDRESS(7), IR_ADD(6) => 
                           IRAM_ADDRESS(6), IR_ADD(5) => IRAM_ADDRESS(5), 
                           IR_ADD(4) => IRAM_ADDRESS(4), IR_ADD(3) => 
                           IRAM_ADDRESS(3), IR_ADD(2) => IRAM_ADDRESS(2), 
                           IR_ADD(1) => IRAM_ADDRESS(1), IR_ADD(0) => 
                           IRAM_ADDRESS(0));

end SYN_structural;
