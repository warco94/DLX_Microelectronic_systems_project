
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_syn is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_syn;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity branch_predictor is

   port( RST : in std_logic;  PC_IN, PC_FAIL, IR_IN : in std_logic_vector (31 
         downto 0);  IR_FAIL : in std_logic_vector (15 downto 0);  WRONG_PRE, 
         RIGHT_PRE : in std_logic;  NPC_OUT, LINK_ADD : out std_logic_vector 
         (31 downto 0);  SEL, TAKEN : out std_logic);

end branch_predictor;

architecture SYN_Behavioral of branch_predictor is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal CACHE_mem_0_1_port, CACHE_mem_0_0_port, CACHE_mem_1_1_port, 
      CACHE_mem_1_0_port, CACHE_mem_2_1_port, CACHE_mem_2_0_port, 
      CACHE_mem_3_1_port, CACHE_mem_3_0_port, CACHE_mem_4_1_port, 
      CACHE_mem_4_0_port, CACHE_mem_5_1_port, CACHE_mem_5_0_port, 
      CACHE_mem_6_1_port, CACHE_mem_6_0_port, CACHE_mem_7_1_port, 
      CACHE_mem_7_0_port, CACHE_mem_8_1_port, CACHE_mem_8_0_port, 
      CACHE_mem_9_1_port, CACHE_mem_9_0_port, CACHE_mem_10_1_port, 
      CACHE_mem_10_0_port, CACHE_mem_11_1_port, CACHE_mem_11_0_port, 
      CACHE_mem_12_1_port, CACHE_mem_12_0_port, CACHE_mem_13_1_port, 
      CACHE_mem_13_0_port, CACHE_mem_14_1_port, CACHE_mem_14_0_port, 
      CACHE_mem_15_1_port, CACHE_mem_15_0_port, CACHE_mem_16_1_port, 
      CACHE_mem_16_0_port, CACHE_mem_17_1_port, CACHE_mem_17_0_port, 
      CACHE_mem_18_1_port, CACHE_mem_18_0_port, CACHE_mem_19_1_port, 
      CACHE_mem_19_0_port, CACHE_mem_20_1_port, CACHE_mem_20_0_port, 
      CACHE_mem_21_1_port, CACHE_mem_21_0_port, CACHE_mem_22_1_port, 
      CACHE_mem_22_0_port, CACHE_mem_23_1_port, CACHE_mem_23_0_port, 
      CACHE_mem_24_1_port, CACHE_mem_24_0_port, CACHE_mem_25_1_port, 
      CACHE_mem_25_0_port, CACHE_mem_26_1_port, CACHE_mem_26_0_port, 
      CACHE_mem_27_1_port, CACHE_mem_27_0_port, CACHE_mem_28_1_port, 
      CACHE_mem_28_0_port, CACHE_mem_29_1_port, CACHE_mem_29_0_port, 
      CACHE_mem_30_1_port, CACHE_mem_30_0_port, CACHE_mem_31_1_port, 
      CACHE_mem_31_0_port, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, 
      N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71
      , N72, N73, N74, N75, N76, N77, N82, N83, N84, N85, N86, N87, N88, N89, 
      N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
      N104, N105, N106, N107, N108, N109, N110, N111, N112, N220, N221, N222, 
      N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, 
      N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, 
      N247, N248, N249, N250, N323, N356, N357, N358, N362, N387, N388, N612, 
      N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, 
      N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, 
      N637, N638, N639, N640, N641, N642, N643, N644, N645, n5, n6, n7, n8, n9,
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n60_port, 
      add_65_carry_2_port, add_65_carry_3_port, add_65_carry_4_port, 
      add_65_carry_5_port, add_65_carry_6_port, add_65_carry_7_port, 
      add_65_carry_8_port, add_65_carry_9_port, add_65_carry_10_port, 
      add_65_carry_11_port, add_65_carry_12_port, add_65_carry_13_port, 
      add_65_carry_14_port, add_65_carry_15_port, add_65_carry_16_port, 
      add_65_carry_17_port, add_65_carry_18_port, add_65_carry_19_port, 
      add_65_carry_20_port, add_65_carry_21_port, add_65_carry_22_port, 
      add_65_carry_23_port, add_65_carry_24_port, add_65_carry_25_port, 
      add_65_carry_26_port, add_65_carry_27_port, add_65_carry_28_port, 
      add_65_carry_29_port, add_65_carry_30_port, add_65_carry_31_port, 
      add_59_n1, add_59_carry_2_port, add_59_carry_3_port, add_59_carry_4_port,
      add_59_carry_5_port, add_59_carry_6_port, add_59_carry_7_port, 
      add_59_carry_8_port, add_59_carry_9_port, add_59_carry_10_port, 
      add_59_carry_11_port, add_59_carry_12_port, add_59_carry_13_port, 
      add_59_carry_14_port, add_59_carry_15_port, add_59_carry_16_port, 
      add_59_carry_17_port, add_59_carry_18_port, add_59_carry_19_port, 
      add_59_carry_20_port, add_59_carry_21_port, add_59_carry_22_port, 
      add_59_carry_23_port, add_59_carry_24_port, add_59_carry_25_port, 
      add_59_carry_26_port, add_59_carry_27_port, add_59_carry_28_port, 
      add_59_carry_29_port, add_59_carry_30_port, add_59_carry_31_port, 
      add_53_aco_n2, add_53_aco_carry_2_port, add_53_aco_carry_3_port, 
      add_53_aco_carry_4_port, add_53_aco_carry_5_port, add_53_aco_carry_6_port
      , add_53_aco_carry_7_port, add_53_aco_carry_8_port, 
      add_53_aco_carry_9_port, add_53_aco_carry_10_port, 
      add_53_aco_carry_11_port, add_53_aco_carry_12_port, 
      add_53_aco_carry_13_port, add_53_aco_carry_14_port, 
      add_53_aco_carry_15_port, add_53_aco_carry_16_port, 
      add_53_aco_carry_17_port, add_53_aco_carry_18_port, 
      add_53_aco_carry_19_port, add_53_aco_carry_20_port, 
      add_53_aco_carry_21_port, add_53_aco_carry_22_port, 
      add_53_aco_carry_23_port, add_53_aco_carry_24_port, 
      add_53_aco_carry_25_port, add_53_aco_carry_26_port, 
      add_53_aco_carry_27_port, add_53_aco_carry_28_port, 
      add_53_aco_carry_29_port, add_53_aco_carry_30_port, 
      add_53_aco_carry_31_port, n62_port, n286, n291, n59_port, n1, n2, n3, n4,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48_port, 
      n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, 
      n56_port, n57_port, n58_port, n61_port, n281, n282, n283, n284, n285, 
      n287, n288, n289, n290, n292, n293, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
      n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, 
      n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, 
      n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
      n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, 
      n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, 
      n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
      n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n_1001, n_1002, n_1003 : std_logic;

begin
   
   NPC_OUT_reg_31_inst : DLH_X1 port map( G => N323, D => n1, Q => NPC_OUT(31))
                           ;
   NPC_OUT_reg_30_inst : DLH_X1 port map( G => N323, D => n2, Q => NPC_OUT(30))
                           ;
   NPC_OUT_reg_29_inst : DLH_X1 port map( G => N323, D => n3, Q => NPC_OUT(29))
                           ;
   NPC_OUT_reg_28_inst : DLH_X1 port map( G => N323, D => n4, Q => NPC_OUT(28))
                           ;
   NPC_OUT_reg_27_inst : DLH_X1 port map( G => N323, D => n20, Q => NPC_OUT(27)
                           );
   NPC_OUT_reg_26_inst : DLH_X1 port map( G => N323, D => n21, Q => NPC_OUT(26)
                           );
   NPC_OUT_reg_25_inst : DLH_X1 port map( G => N323, D => n22, Q => NPC_OUT(25)
                           );
   NPC_OUT_reg_24_inst : DLH_X1 port map( G => N323, D => n23, Q => NPC_OUT(24)
                           );
   NPC_OUT_reg_23_inst : DLH_X1 port map( G => N323, D => n24, Q => NPC_OUT(23)
                           );
   NPC_OUT_reg_22_inst : DLH_X1 port map( G => N323, D => n25, Q => NPC_OUT(22)
                           );
   NPC_OUT_reg_21_inst : DLH_X1 port map( G => N323, D => n26, Q => NPC_OUT(21)
                           );
   NPC_OUT_reg_20_inst : DLH_X1 port map( G => N323, D => n27, Q => NPC_OUT(20)
                           );
   NPC_OUT_reg_19_inst : DLH_X1 port map( G => N323, D => n28, Q => NPC_OUT(19)
                           );
   NPC_OUT_reg_18_inst : DLH_X1 port map( G => N323, D => n29, Q => NPC_OUT(18)
                           );
   NPC_OUT_reg_17_inst : DLH_X1 port map( G => N323, D => n30, Q => NPC_OUT(17)
                           );
   NPC_OUT_reg_16_inst : DLH_X1 port map( G => N323, D => n31, Q => NPC_OUT(16)
                           );
   NPC_OUT_reg_15_inst : DLH_X1 port map( G => N323, D => n32, Q => NPC_OUT(15)
                           );
   NPC_OUT_reg_14_inst : DLH_X1 port map( G => N323, D => n33, Q => NPC_OUT(14)
                           );
   NPC_OUT_reg_13_inst : DLH_X1 port map( G => N323, D => n34, Q => NPC_OUT(13)
                           );
   NPC_OUT_reg_12_inst : DLH_X1 port map( G => N323, D => n35, Q => NPC_OUT(12)
                           );
   NPC_OUT_reg_11_inst : DLH_X1 port map( G => N323, D => n36, Q => NPC_OUT(11)
                           );
   NPC_OUT_reg_10_inst : DLH_X1 port map( G => N323, D => n37, Q => NPC_OUT(10)
                           );
   NPC_OUT_reg_9_inst : DLH_X1 port map( G => N323, D => n38, Q => NPC_OUT(9));
   NPC_OUT_reg_8_inst : DLH_X1 port map( G => N323, D => n39, Q => NPC_OUT(8));
   NPC_OUT_reg_7_inst : DLH_X1 port map( G => N323, D => n40, Q => NPC_OUT(7));
   NPC_OUT_reg_6_inst : DLH_X1 port map( G => N323, D => n41, Q => NPC_OUT(6));
   NPC_OUT_reg_5_inst : DLH_X1 port map( G => N323, D => n42, Q => NPC_OUT(5));
   NPC_OUT_reg_4_inst : DLH_X1 port map( G => N323, D => n43, Q => NPC_OUT(4));
   NPC_OUT_reg_3_inst : DLH_X1 port map( G => N323, D => n44, Q => NPC_OUT(3));
   NPC_OUT_reg_2_inst : DLH_X1 port map( G => N323, D => n45, Q => NPC_OUT(2));
   NPC_OUT_reg_1_inst : DLH_X1 port map( G => N323, D => n46, Q => NPC_OUT(1));
   NPC_OUT_reg_0_inst : DLH_X1 port map( G => N323, D => n60_port, Q => 
                           NPC_OUT(0));
   LINK_ADD_reg_31_inst : DLH_X1 port map( G => N356, D => N388, Q => 
                           LINK_ADD(31));
   LINK_ADD_reg_30_inst : DLH_X1 port map( G => N356, D => N387, Q => 
                           LINK_ADD(30));
   LINK_ADD_reg_29_inst : DLH_X1 port map( G => n5092, D => n48_port, Q => 
                           LINK_ADD(29));
   LINK_ADD_reg_28_inst : DLH_X1 port map( G => n5092, D => n287, Q => 
                           LINK_ADD(28));
   LINK_ADD_reg_27_inst : DLH_X1 port map( G => n5092, D => n49_port, Q => 
                           LINK_ADD(27));
   LINK_ADD_reg_26_inst : DLH_X1 port map( G => n5092, D => n283, Q => 
                           LINK_ADD(26));
   LINK_ADD_reg_25_inst : DLH_X1 port map( G => n5092, D => n50_port, Q => 
                           LINK_ADD(25));
   LINK_ADD_reg_24_inst : DLH_X1 port map( G => n5092, D => n293, Q => 
                           LINK_ADD(24));
   LINK_ADD_reg_23_inst : DLH_X1 port map( G => n5092, D => n51_port, Q => 
                           LINK_ADD(23));
   LINK_ADD_reg_22_inst : DLH_X1 port map( G => n5092, D => n290, Q => 
                           LINK_ADD(22));
   LINK_ADD_reg_21_inst : DLH_X1 port map( G => n5092, D => n52_port, Q => 
                           LINK_ADD(21));
   LINK_ADD_reg_20_inst : DLH_X1 port map( G => n5092, D => n289, Q => 
                           LINK_ADD(20));
   LINK_ADD_reg_19_inst : DLH_X1 port map( G => n5092, D => n53_port, Q => 
                           LINK_ADD(19));
   LINK_ADD_reg_18_inst : DLH_X1 port map( G => n5092, D => n288, Q => 
                           LINK_ADD(18));
   LINK_ADD_reg_17_inst : DLH_X1 port map( G => n5092, D => n54_port, Q => 
                           LINK_ADD(17));
   LINK_ADD_reg_16_inst : DLH_X1 port map( G => n5092, D => n285, Q => 
                           LINK_ADD(16));
   LINK_ADD_reg_15_inst : DLH_X1 port map( G => n5092, D => n55_port, Q => 
                           LINK_ADD(15));
   LINK_ADD_reg_14_inst : DLH_X1 port map( G => n5092, D => n284, Q => 
                           LINK_ADD(14));
   LINK_ADD_reg_13_inst : DLH_X1 port map( G => n5092, D => n56_port, Q => 
                           LINK_ADD(13));
   LINK_ADD_reg_12_inst : DLH_X1 port map( G => n5092, D => n292, Q => 
                           LINK_ADD(12));
   LINK_ADD_reg_11_inst : DLH_X1 port map( G => n5092, D => n57_port, Q => 
                           LINK_ADD(11));
   LINK_ADD_reg_10_inst : DLH_X1 port map( G => n5092, D => n281, Q => 
                           LINK_ADD(10));
   LINK_ADD_reg_9_inst : DLH_X1 port map( G => n5092, D => n58_port, Q => 
                           LINK_ADD(9));
   LINK_ADD_reg_8_inst : DLH_X1 port map( G => n5092, D => n282, Q => 
                           LINK_ADD(8));
   LINK_ADD_reg_7_inst : DLH_X1 port map( G => N356, D => n61_port, Q => 
                           LINK_ADD(7));
   LINK_ADD_reg_6_inst : DLH_X1 port map( G => N356, D => n291, Q => 
                           LINK_ADD(6));
   LINK_ADD_reg_5_inst : DLH_X1 port map( G => N356, D => N362, Q => 
                           LINK_ADD(5));
   LINK_ADD_reg_4_inst : DLH_X1 port map( G => N356, D => n286, Q => 
                           LINK_ADD(4));
   LINK_ADD_reg_3_inst : DLH_X1 port map( G => N356, D => n59_port, Q => 
                           LINK_ADD(3));
   LINK_ADD_reg_2_inst : DLH_X1 port map( G => N356, D => n62_port, Q => 
                           LINK_ADD(2));
   LINK_ADD_reg_1_inst : DLH_X1 port map( G => N356, D => N358, Q => 
                           LINK_ADD(1));
   LINK_ADD_reg_0_inst : DLH_X1 port map( G => N356, D => N357, Q => 
                           LINK_ADD(0));
   CACHE_mem_reg_0_1_inst : DLH_X1 port map( G => N643, D => N645, Q => 
                           CACHE_mem_0_1_port);
   CACHE_mem_reg_0_0_inst : DLH_X1 port map( G => N643, D => N644, Q => 
                           CACHE_mem_0_0_port);
   CACHE_mem_reg_1_1_inst : DLH_X1 port map( G => N642, D => N645, Q => 
                           CACHE_mem_1_1_port);
   CACHE_mem_reg_1_0_inst : DLH_X1 port map( G => N642, D => N644, Q => 
                           CACHE_mem_1_0_port);
   CACHE_mem_reg_2_1_inst : DLH_X1 port map( G => N641, D => N645, Q => 
                           CACHE_mem_2_1_port);
   CACHE_mem_reg_2_0_inst : DLH_X1 port map( G => N641, D => N644, Q => 
                           CACHE_mem_2_0_port);
   CACHE_mem_reg_3_1_inst : DLH_X1 port map( G => N640, D => N645, Q => 
                           CACHE_mem_3_1_port);
   CACHE_mem_reg_3_0_inst : DLH_X1 port map( G => N640, D => N644, Q => 
                           CACHE_mem_3_0_port);
   CACHE_mem_reg_4_1_inst : DLH_X1 port map( G => N639, D => N645, Q => 
                           CACHE_mem_4_1_port);
   CACHE_mem_reg_4_0_inst : DLH_X1 port map( G => N639, D => N644, Q => 
                           CACHE_mem_4_0_port);
   CACHE_mem_reg_5_1_inst : DLH_X1 port map( G => N638, D => N645, Q => 
                           CACHE_mem_5_1_port);
   CACHE_mem_reg_5_0_inst : DLH_X1 port map( G => N638, D => N644, Q => 
                           CACHE_mem_5_0_port);
   CACHE_mem_reg_6_1_inst : DLH_X1 port map( G => N637, D => N645, Q => 
                           CACHE_mem_6_1_port);
   CACHE_mem_reg_6_0_inst : DLH_X1 port map( G => N637, D => N644, Q => 
                           CACHE_mem_6_0_port);
   CACHE_mem_reg_7_1_inst : DLH_X1 port map( G => N636, D => N645, Q => 
                           CACHE_mem_7_1_port);
   CACHE_mem_reg_7_0_inst : DLH_X1 port map( G => N636, D => N644, Q => 
                           CACHE_mem_7_0_port);
   CACHE_mem_reg_8_1_inst : DLH_X1 port map( G => N635, D => N645, Q => 
                           CACHE_mem_8_1_port);
   CACHE_mem_reg_8_0_inst : DLH_X1 port map( G => N635, D => N644, Q => 
                           CACHE_mem_8_0_port);
   CACHE_mem_reg_9_1_inst : DLH_X1 port map( G => N634, D => N645, Q => 
                           CACHE_mem_9_1_port);
   CACHE_mem_reg_9_0_inst : DLH_X1 port map( G => N634, D => N644, Q => 
                           CACHE_mem_9_0_port);
   CACHE_mem_reg_10_1_inst : DLH_X1 port map( G => N633, D => N645, Q => 
                           CACHE_mem_10_1_port);
   CACHE_mem_reg_10_0_inst : DLH_X1 port map( G => N633, D => N644, Q => 
                           CACHE_mem_10_0_port);
   CACHE_mem_reg_11_1_inst : DLH_X1 port map( G => N632, D => N645, Q => 
                           CACHE_mem_11_1_port);
   CACHE_mem_reg_11_0_inst : DLH_X1 port map( G => N632, D => N644, Q => 
                           CACHE_mem_11_0_port);
   CACHE_mem_reg_12_1_inst : DLH_X1 port map( G => N631, D => N645, Q => 
                           CACHE_mem_12_1_port);
   CACHE_mem_reg_12_0_inst : DLH_X1 port map( G => N631, D => N644, Q => 
                           CACHE_mem_12_0_port);
   CACHE_mem_reg_13_1_inst : DLH_X1 port map( G => N630, D => N645, Q => 
                           CACHE_mem_13_1_port);
   CACHE_mem_reg_13_0_inst : DLH_X1 port map( G => N630, D => N644, Q => 
                           CACHE_mem_13_0_port);
   CACHE_mem_reg_14_1_inst : DLH_X1 port map( G => N629, D => N645, Q => 
                           CACHE_mem_14_1_port);
   CACHE_mem_reg_14_0_inst : DLH_X1 port map( G => N629, D => N644, Q => 
                           CACHE_mem_14_0_port);
   CACHE_mem_reg_15_1_inst : DLH_X1 port map( G => N628, D => N645, Q => 
                           CACHE_mem_15_1_port);
   CACHE_mem_reg_15_0_inst : DLH_X1 port map( G => N628, D => N644, Q => 
                           CACHE_mem_15_0_port);
   CACHE_mem_reg_16_1_inst : DLH_X1 port map( G => N627, D => N645, Q => 
                           CACHE_mem_16_1_port);
   CACHE_mem_reg_16_0_inst : DLH_X1 port map( G => N627, D => N644, Q => 
                           CACHE_mem_16_0_port);
   CACHE_mem_reg_17_1_inst : DLH_X1 port map( G => N626, D => N645, Q => 
                           CACHE_mem_17_1_port);
   CACHE_mem_reg_17_0_inst : DLH_X1 port map( G => N626, D => N644, Q => 
                           CACHE_mem_17_0_port);
   CACHE_mem_reg_18_1_inst : DLH_X1 port map( G => N625, D => N645, Q => 
                           CACHE_mem_18_1_port);
   CACHE_mem_reg_18_0_inst : DLH_X1 port map( G => N625, D => N644, Q => 
                           CACHE_mem_18_0_port);
   CACHE_mem_reg_19_1_inst : DLH_X1 port map( G => N624, D => N645, Q => 
                           CACHE_mem_19_1_port);
   CACHE_mem_reg_19_0_inst : DLH_X1 port map( G => N624, D => N644, Q => 
                           CACHE_mem_19_0_port);
   CACHE_mem_reg_20_1_inst : DLH_X1 port map( G => N623, D => N645, Q => 
                           CACHE_mem_20_1_port);
   CACHE_mem_reg_20_0_inst : DLH_X1 port map( G => N623, D => N644, Q => 
                           CACHE_mem_20_0_port);
   CACHE_mem_reg_21_1_inst : DLH_X1 port map( G => N622, D => N645, Q => 
                           CACHE_mem_21_1_port);
   CACHE_mem_reg_21_0_inst : DLH_X1 port map( G => N622, D => N644, Q => 
                           CACHE_mem_21_0_port);
   CACHE_mem_reg_22_1_inst : DLH_X1 port map( G => N621, D => N645, Q => 
                           CACHE_mem_22_1_port);
   CACHE_mem_reg_22_0_inst : DLH_X1 port map( G => N621, D => N644, Q => 
                           CACHE_mem_22_0_port);
   CACHE_mem_reg_23_1_inst : DLH_X1 port map( G => N620, D => N645, Q => 
                           CACHE_mem_23_1_port);
   CACHE_mem_reg_23_0_inst : DLH_X1 port map( G => N620, D => N644, Q => 
                           CACHE_mem_23_0_port);
   CACHE_mem_reg_24_1_inst : DLH_X1 port map( G => N619, D => N645, Q => 
                           CACHE_mem_24_1_port);
   CACHE_mem_reg_24_0_inst : DLH_X1 port map( G => N619, D => N644, Q => 
                           CACHE_mem_24_0_port);
   CACHE_mem_reg_25_1_inst : DLH_X1 port map( G => N618, D => N645, Q => 
                           CACHE_mem_25_1_port);
   CACHE_mem_reg_25_0_inst : DLH_X1 port map( G => N618, D => N644, Q => 
                           CACHE_mem_25_0_port);
   CACHE_mem_reg_26_1_inst : DLH_X1 port map( G => N617, D => N645, Q => 
                           CACHE_mem_26_1_port);
   CACHE_mem_reg_26_0_inst : DLH_X1 port map( G => N617, D => N644, Q => 
                           CACHE_mem_26_0_port);
   CACHE_mem_reg_27_1_inst : DLH_X1 port map( G => N616, D => N645, Q => 
                           CACHE_mem_27_1_port);
   CACHE_mem_reg_27_0_inst : DLH_X1 port map( G => N616, D => N644, Q => 
                           CACHE_mem_27_0_port);
   CACHE_mem_reg_28_1_inst : DLH_X1 port map( G => N615, D => N645, Q => 
                           CACHE_mem_28_1_port);
   CACHE_mem_reg_28_0_inst : DLH_X1 port map( G => N615, D => N644, Q => 
                           CACHE_mem_28_0_port);
   CACHE_mem_reg_29_1_inst : DLH_X1 port map( G => N614, D => N645, Q => 
                           CACHE_mem_29_1_port);
   CACHE_mem_reg_29_0_inst : DLH_X1 port map( G => N614, D => N644, Q => 
                           CACHE_mem_29_0_port);
   CACHE_mem_reg_30_1_inst : DLH_X1 port map( G => N613, D => N645, Q => 
                           CACHE_mem_30_1_port);
   CACHE_mem_reg_30_0_inst : DLH_X1 port map( G => N613, D => N644, Q => 
                           CACHE_mem_30_0_port);
   CACHE_mem_reg_31_1_inst : DLH_X1 port map( G => N612, D => N645, Q => 
                           CACHE_mem_31_1_port);
   CACHE_mem_reg_31_0_inst : DLH_X1 port map( G => N612, D => N644, Q => 
                           CACHE_mem_31_0_port);
   add_65_U1_1 : FA_X1 port map( A => PC_IN(1), B => IR_IN(1), CI => add_59_n1,
                           CO => add_65_carry_2_port, S => N220);
   add_65_U1_2 : FA_X1 port map( A => PC_IN(2), B => IR_IN(2), CI => 
                           add_65_carry_2_port, CO => add_65_carry_3_port, S =>
                           N221);
   add_65_U1_3 : FA_X1 port map( A => PC_IN(3), B => IR_IN(3), CI => 
                           add_65_carry_3_port, CO => add_65_carry_4_port, S =>
                           N222);
   add_65_U1_4 : FA_X1 port map( A => PC_IN(4), B => IR_IN(4), CI => 
                           add_65_carry_4_port, CO => add_65_carry_5_port, S =>
                           N223);
   add_65_U1_5 : FA_X1 port map( A => PC_IN(5), B => IR_IN(5), CI => 
                           add_65_carry_5_port, CO => add_65_carry_6_port, S =>
                           N224);
   add_65_U1_6 : FA_X1 port map( A => PC_IN(6), B => IR_IN(6), CI => 
                           add_65_carry_6_port, CO => add_65_carry_7_port, S =>
                           N225);
   add_65_U1_7 : FA_X1 port map( A => PC_IN(7), B => IR_IN(7), CI => 
                           add_65_carry_7_port, CO => add_65_carry_8_port, S =>
                           N226);
   add_65_U1_8 : FA_X1 port map( A => PC_IN(8), B => IR_IN(8), CI => 
                           add_65_carry_8_port, CO => add_65_carry_9_port, S =>
                           N227);
   add_65_U1_9 : FA_X1 port map( A => PC_IN(9), B => IR_IN(9), CI => 
                           add_65_carry_9_port, CO => add_65_carry_10_port, S 
                           => N228);
   add_65_U1_10 : FA_X1 port map( A => PC_IN(10), B => IR_IN(10), CI => 
                           add_65_carry_10_port, CO => add_65_carry_11_port, S 
                           => N229);
   add_65_U1_11 : FA_X1 port map( A => PC_IN(11), B => IR_IN(11), CI => 
                           add_65_carry_11_port, CO => add_65_carry_12_port, S 
                           => N230);
   add_65_U1_12 : FA_X1 port map( A => PC_IN(12), B => IR_IN(12), CI => 
                           add_65_carry_12_port, CO => add_65_carry_13_port, S 
                           => N231);
   add_65_U1_13 : FA_X1 port map( A => PC_IN(13), B => IR_IN(13), CI => 
                           add_65_carry_13_port, CO => add_65_carry_14_port, S 
                           => N232);
   add_65_U1_14 : FA_X1 port map( A => PC_IN(14), B => IR_IN(14), CI => 
                           add_65_carry_14_port, CO => add_65_carry_15_port, S 
                           => N233);
   add_65_U1_15 : FA_X1 port map( A => PC_IN(15), B => IR_IN(15), CI => 
                           add_65_carry_15_port, CO => add_65_carry_16_port, S 
                           => N234);
   add_65_U1_16 : FA_X1 port map( A => PC_IN(16), B => IR_IN(15), CI => 
                           add_65_carry_16_port, CO => add_65_carry_17_port, S 
                           => N235);
   add_65_U1_17 : FA_X1 port map( A => PC_IN(17), B => IR_IN(15), CI => 
                           add_65_carry_17_port, CO => add_65_carry_18_port, S 
                           => N236);
   add_65_U1_18 : FA_X1 port map( A => PC_IN(18), B => IR_IN(15), CI => 
                           add_65_carry_18_port, CO => add_65_carry_19_port, S 
                           => N237);
   add_65_U1_19 : FA_X1 port map( A => PC_IN(19), B => IR_IN(15), CI => 
                           add_65_carry_19_port, CO => add_65_carry_20_port, S 
                           => N238);
   add_65_U1_20 : FA_X1 port map( A => PC_IN(20), B => IR_IN(15), CI => 
                           add_65_carry_20_port, CO => add_65_carry_21_port, S 
                           => N239);
   add_65_U1_21 : FA_X1 port map( A => PC_IN(21), B => IR_IN(15), CI => 
                           add_65_carry_21_port, CO => add_65_carry_22_port, S 
                           => N240);
   add_65_U1_22 : FA_X1 port map( A => PC_IN(22), B => IR_IN(15), CI => 
                           add_65_carry_22_port, CO => add_65_carry_23_port, S 
                           => N241);
   add_65_U1_23 : FA_X1 port map( A => PC_IN(23), B => IR_IN(15), CI => 
                           add_65_carry_23_port, CO => add_65_carry_24_port, S 
                           => N242);
   add_65_U1_24 : FA_X1 port map( A => PC_IN(24), B => IR_IN(15), CI => 
                           add_65_carry_24_port, CO => add_65_carry_25_port, S 
                           => N243);
   add_65_U1_25 : FA_X1 port map( A => PC_IN(25), B => IR_IN(15), CI => 
                           add_65_carry_25_port, CO => add_65_carry_26_port, S 
                           => N244);
   add_65_U1_26 : FA_X1 port map( A => PC_IN(26), B => IR_IN(15), CI => 
                           add_65_carry_26_port, CO => add_65_carry_27_port, S 
                           => N245);
   add_65_U1_27 : FA_X1 port map( A => PC_IN(27), B => IR_IN(15), CI => 
                           add_65_carry_27_port, CO => add_65_carry_28_port, S 
                           => N246);
   add_65_U1_28 : FA_X1 port map( A => PC_IN(28), B => IR_IN(15), CI => 
                           add_65_carry_28_port, CO => add_65_carry_29_port, S 
                           => N247);
   add_65_U1_29 : FA_X1 port map( A => PC_IN(29), B => IR_IN(15), CI => 
                           add_65_carry_29_port, CO => add_65_carry_30_port, S 
                           => N248);
   add_65_U1_30 : FA_X1 port map( A => PC_IN(30), B => IR_IN(15), CI => 
                           add_65_carry_30_port, CO => add_65_carry_31_port, S 
                           => N249);
   add_65_U1_31 : FA_X1 port map( A => PC_IN(31), B => IR_IN(15), CI => 
                           add_65_carry_31_port, CO => n_1001, S => N250);
   add_59_U1_1 : FA_X1 port map( A => PC_IN(1), B => IR_IN(1), CI => add_59_n1,
                           CO => add_59_carry_2_port, S => N82);
   add_59_U1_2 : FA_X1 port map( A => PC_IN(2), B => IR_IN(2), CI => 
                           add_59_carry_2_port, CO => add_59_carry_3_port, S =>
                           N83);
   add_59_U1_3 : FA_X1 port map( A => PC_IN(3), B => IR_IN(3), CI => 
                           add_59_carry_3_port, CO => add_59_carry_4_port, S =>
                           N84);
   add_59_U1_4 : FA_X1 port map( A => PC_IN(4), B => IR_IN(4), CI => 
                           add_59_carry_4_port, CO => add_59_carry_5_port, S =>
                           N85);
   add_59_U1_5 : FA_X1 port map( A => PC_IN(5), B => IR_IN(5), CI => 
                           add_59_carry_5_port, CO => add_59_carry_6_port, S =>
                           N86);
   add_59_U1_6 : FA_X1 port map( A => PC_IN(6), B => IR_IN(6), CI => 
                           add_59_carry_6_port, CO => add_59_carry_7_port, S =>
                           N87);
   add_59_U1_7 : FA_X1 port map( A => PC_IN(7), B => IR_IN(7), CI => 
                           add_59_carry_7_port, CO => add_59_carry_8_port, S =>
                           N88);
   add_59_U1_8 : FA_X1 port map( A => PC_IN(8), B => IR_IN(8), CI => 
                           add_59_carry_8_port, CO => add_59_carry_9_port, S =>
                           N89);
   add_59_U1_9 : FA_X1 port map( A => PC_IN(9), B => IR_IN(9), CI => 
                           add_59_carry_9_port, CO => add_59_carry_10_port, S 
                           => N90);
   add_59_U1_10 : FA_X1 port map( A => PC_IN(10), B => IR_IN(10), CI => 
                           add_59_carry_10_port, CO => add_59_carry_11_port, S 
                           => N91);
   add_59_U1_11 : FA_X1 port map( A => PC_IN(11), B => IR_IN(11), CI => 
                           add_59_carry_11_port, CO => add_59_carry_12_port, S 
                           => N92);
   add_59_U1_12 : FA_X1 port map( A => PC_IN(12), B => IR_IN(12), CI => 
                           add_59_carry_12_port, CO => add_59_carry_13_port, S 
                           => N93);
   add_59_U1_13 : FA_X1 port map( A => PC_IN(13), B => IR_IN(13), CI => 
                           add_59_carry_13_port, CO => add_59_carry_14_port, S 
                           => N94);
   add_59_U1_14 : FA_X1 port map( A => PC_IN(14), B => IR_IN(14), CI => 
                           add_59_carry_14_port, CO => add_59_carry_15_port, S 
                           => N95);
   add_59_U1_15 : FA_X1 port map( A => PC_IN(15), B => IR_IN(15), CI => 
                           add_59_carry_15_port, CO => add_59_carry_16_port, S 
                           => N96);
   add_59_U1_16 : FA_X1 port map( A => PC_IN(16), B => IR_IN(16), CI => 
                           add_59_carry_16_port, CO => add_59_carry_17_port, S 
                           => N97);
   add_59_U1_17 : FA_X1 port map( A => PC_IN(17), B => IR_IN(17), CI => 
                           add_59_carry_17_port, CO => add_59_carry_18_port, S 
                           => N98);
   add_59_U1_18 : FA_X1 port map( A => PC_IN(18), B => IR_IN(18), CI => 
                           add_59_carry_18_port, CO => add_59_carry_19_port, S 
                           => N99);
   add_59_U1_19 : FA_X1 port map( A => PC_IN(19), B => IR_IN(19), CI => 
                           add_59_carry_19_port, CO => add_59_carry_20_port, S 
                           => N100);
   add_59_U1_20 : FA_X1 port map( A => PC_IN(20), B => IR_IN(20), CI => 
                           add_59_carry_20_port, CO => add_59_carry_21_port, S 
                           => N101);
   add_59_U1_21 : FA_X1 port map( A => PC_IN(21), B => IR_IN(21), CI => 
                           add_59_carry_21_port, CO => add_59_carry_22_port, S 
                           => N102);
   add_59_U1_22 : FA_X1 port map( A => PC_IN(22), B => IR_IN(22), CI => 
                           add_59_carry_22_port, CO => add_59_carry_23_port, S 
                           => N103);
   add_59_U1_23 : FA_X1 port map( A => PC_IN(23), B => IR_IN(23), CI => 
                           add_59_carry_23_port, CO => add_59_carry_24_port, S 
                           => N104);
   add_59_U1_24 : FA_X1 port map( A => PC_IN(24), B => IR_IN(24), CI => 
                           add_59_carry_24_port, CO => add_59_carry_25_port, S 
                           => N105);
   add_59_U1_25 : FA_X1 port map( A => PC_IN(25), B => IR_IN(25), CI => 
                           add_59_carry_25_port, CO => add_59_carry_26_port, S 
                           => N106);
   add_59_U1_26 : FA_X1 port map( A => PC_IN(26), B => IR_IN(25), CI => 
                           add_59_carry_26_port, CO => add_59_carry_27_port, S 
                           => N107);
   add_59_U1_27 : FA_X1 port map( A => PC_IN(27), B => IR_IN(25), CI => 
                           add_59_carry_27_port, CO => add_59_carry_28_port, S 
                           => N108);
   add_59_U1_28 : FA_X1 port map( A => PC_IN(28), B => IR_IN(25), CI => 
                           add_59_carry_28_port, CO => add_59_carry_29_port, S 
                           => N109);
   add_59_U1_29 : FA_X1 port map( A => PC_IN(29), B => IR_IN(25), CI => 
                           add_59_carry_29_port, CO => add_59_carry_30_port, S 
                           => N110);
   add_59_U1_30 : FA_X1 port map( A => PC_IN(30), B => IR_IN(25), CI => 
                           add_59_carry_30_port, CO => add_59_carry_31_port, S 
                           => N111);
   add_59_U1_31 : FA_X1 port map( A => PC_IN(31), B => IR_IN(25), CI => 
                           add_59_carry_31_port, CO => n_1002, S => N112);
   add_53_aco_U1_1 : FA_X1 port map( A => PC_FAIL(1), B => n6, CI => 
                           add_53_aco_n2, CO => add_53_aco_carry_2_port, S => 
                           N47);
   add_53_aco_U1_2 : FA_X1 port map( A => PC_FAIL(2), B => n8, CI => 
                           add_53_aco_carry_2_port, CO => 
                           add_53_aco_carry_3_port, S => N48);
   add_53_aco_U1_3 : FA_X1 port map( A => PC_FAIL(3), B => n9, CI => 
                           add_53_aco_carry_3_port, CO => 
                           add_53_aco_carry_4_port, S => N49);
   add_53_aco_U1_4 : FA_X1 port map( A => PC_FAIL(4), B => n10, CI => 
                           add_53_aco_carry_4_port, CO => 
                           add_53_aco_carry_5_port, S => N50);
   add_53_aco_U1_5 : FA_X1 port map( A => PC_FAIL(5), B => n7, CI => 
                           add_53_aco_carry_5_port, CO => 
                           add_53_aco_carry_6_port, S => N51);
   add_53_aco_U1_6 : FA_X1 port map( A => PC_FAIL(6), B => n11, CI => 
                           add_53_aco_carry_6_port, CO => 
                           add_53_aco_carry_7_port, S => N52);
   add_53_aco_U1_7 : FA_X1 port map( A => PC_FAIL(7), B => n12, CI => 
                           add_53_aco_carry_7_port, CO => 
                           add_53_aco_carry_8_port, S => N53);
   add_53_aco_U1_8 : FA_X1 port map( A => PC_FAIL(8), B => n13, CI => 
                           add_53_aco_carry_8_port, CO => 
                           add_53_aco_carry_9_port, S => N54);
   add_53_aco_U1_9 : FA_X1 port map( A => PC_FAIL(9), B => n14, CI => 
                           add_53_aco_carry_9_port, CO => 
                           add_53_aco_carry_10_port, S => N55);
   add_53_aco_U1_10 : FA_X1 port map( A => PC_FAIL(10), B => n15, CI => 
                           add_53_aco_carry_10_port, CO => 
                           add_53_aco_carry_11_port, S => N56);
   add_53_aco_U1_11 : FA_X1 port map( A => PC_FAIL(11), B => n16, CI => 
                           add_53_aco_carry_11_port, CO => 
                           add_53_aco_carry_12_port, S => N57);
   add_53_aco_U1_12 : FA_X1 port map( A => PC_FAIL(12), B => n17, CI => 
                           add_53_aco_carry_12_port, CO => 
                           add_53_aco_carry_13_port, S => N58);
   add_53_aco_U1_13 : FA_X1 port map( A => PC_FAIL(13), B => n18, CI => 
                           add_53_aco_carry_13_port, CO => 
                           add_53_aco_carry_14_port, S => N59);
   add_53_aco_U1_14 : FA_X1 port map( A => PC_FAIL(14), B => n19, CI => 
                           add_53_aco_carry_14_port, CO => 
                           add_53_aco_carry_15_port, S => N60);
   add_53_aco_U1_15 : FA_X1 port map( A => PC_FAIL(15), B => n5, CI => 
                           add_53_aco_carry_15_port, CO => 
                           add_53_aco_carry_16_port, S => N61);
   add_53_aco_U1_16 : FA_X1 port map( A => PC_FAIL(16), B => n5, CI => 
                           add_53_aco_carry_16_port, CO => 
                           add_53_aco_carry_17_port, S => N62);
   add_53_aco_U1_17 : FA_X1 port map( A => PC_FAIL(17), B => n5, CI => 
                           add_53_aco_carry_17_port, CO => 
                           add_53_aco_carry_18_port, S => N63);
   add_53_aco_U1_18 : FA_X1 port map( A => PC_FAIL(18), B => n5, CI => 
                           add_53_aco_carry_18_port, CO => 
                           add_53_aco_carry_19_port, S => N64);
   add_53_aco_U1_19 : FA_X1 port map( A => PC_FAIL(19), B => n5, CI => 
                           add_53_aco_carry_19_port, CO => 
                           add_53_aco_carry_20_port, S => N65);
   add_53_aco_U1_20 : FA_X1 port map( A => PC_FAIL(20), B => n5, CI => 
                           add_53_aco_carry_20_port, CO => 
                           add_53_aco_carry_21_port, S => N66);
   add_53_aco_U1_21 : FA_X1 port map( A => PC_FAIL(21), B => n5, CI => 
                           add_53_aco_carry_21_port, CO => 
                           add_53_aco_carry_22_port, S => N67);
   add_53_aco_U1_22 : FA_X1 port map( A => PC_FAIL(22), B => n5, CI => 
                           add_53_aco_carry_22_port, CO => 
                           add_53_aco_carry_23_port, S => N68);
   add_53_aco_U1_23 : FA_X1 port map( A => PC_FAIL(23), B => n5, CI => 
                           add_53_aco_carry_23_port, CO => 
                           add_53_aco_carry_24_port, S => N69);
   add_53_aco_U1_24 : FA_X1 port map( A => PC_FAIL(24), B => n5, CI => 
                           add_53_aco_carry_24_port, CO => 
                           add_53_aco_carry_25_port, S => N70);
   add_53_aco_U1_25 : FA_X1 port map( A => PC_FAIL(25), B => n5, CI => 
                           add_53_aco_carry_25_port, CO => 
                           add_53_aco_carry_26_port, S => N71);
   add_53_aco_U1_26 : FA_X1 port map( A => PC_FAIL(26), B => n5, CI => 
                           add_53_aco_carry_26_port, CO => 
                           add_53_aco_carry_27_port, S => N72);
   add_53_aco_U1_27 : FA_X1 port map( A => PC_FAIL(27), B => n5, CI => 
                           add_53_aco_carry_27_port, CO => 
                           add_53_aco_carry_28_port, S => N73);
   add_53_aco_U1_28 : FA_X1 port map( A => PC_FAIL(28), B => n5, CI => 
                           add_53_aco_carry_28_port, CO => 
                           add_53_aco_carry_29_port, S => N74);
   add_53_aco_U1_29 : FA_X1 port map( A => PC_FAIL(29), B => n5, CI => 
                           add_53_aco_carry_29_port, CO => 
                           add_53_aco_carry_30_port, S => N75);
   add_53_aco_U1_30 : FA_X1 port map( A => PC_FAIL(30), B => n5, CI => 
                           add_53_aco_carry_30_port, CO => 
                           add_53_aco_carry_31_port, S => N76);
   add_53_aco_U1_31 : FA_X1 port map( A => PC_FAIL(31), B => n5, CI => 
                           add_53_aco_carry_31_port, CO => n_1003, S => N77);
   U3 : NAND2_X1 port map( A1 => n5317, A2 => n5225, ZN => N323);
   U4 : INV_X2 port map( A => n5224, ZN => n5317);
   U5 : NOR2_X2 port map( A1 => n5222, A2 => n5090, ZN => N644);
   U6 : INV_X2 port map( A => n5090, ZN => n5089);
   U7 : NOR3_X2 port map( A1 => PC_FAIL(4), A2 => n5143, A3 => n5145, ZN => 
                           n5205);
   U8 : AOI211_X1 port map( C1 => n5202, C2 => CACHE_mem_26_1_port, A => n5192,
                           B => n5191, ZN => n5216);
   U9 : NOR3_X2 port map( A1 => PC_FAIL(2), A2 => PC_FAIL(4), A3 => n5145, ZN 
                           => n5202);
   U10 : NOR3_X2 port map( A1 => PC_FAIL(4), A2 => PC_FAIL(3), A3 => n5143, ZN 
                           => n5203);
   U11 : NOR3_X2 port map( A1 => PC_FAIL(2), A2 => PC_FAIL(4), A3 => PC_FAIL(3)
                           , ZN => n5207);
   U12 : AOI211_X4 port map( C1 => n5218, C2 => n5217, A => n5216, B => n5215, 
                           ZN => n5236);
   U13 : INV_X1 port map( A => n5202, ZN => n5178);
   U14 : INV_X1 port map( A => n5203, ZN => n5179);
   U15 : INV_X1 port map( A => n5207, ZN => n5181);
   U16 : BUF_X1 port map( A => N356, Z => n5092);
   U17 : OAI221_X1 port map( B1 => n5093, B2 => n5284, C1 => n5093, C2 => n5225
                           , A => n5090, ZN => SEL);
   U18 : INV_X1 port map( A => RST, ZN => n5093);
   U19 : BUF_X1 port map( A => n5316, Z => n5091);
   U20 : NOR2_X1 port map( A1 => n5285, A2 => n5284, ZN => n5316);
   U21 : OR2_X1 port map( A1 => n5094, A2 => n5219, ZN => n5090);
   U22 : AND2_X1 port map( A1 => RST, A2 => n5223, ZN => N645);
   U23 : INV_X1 port map( A => n5205, ZN => n5187);
   U24 : INV_X1 port map( A => PC_FAIL(5), ZN => n5199);
   U25 : INV_X1 port map( A => RST, ZN => n5094);
   U26 : INV_X1 port map( A => IR_IN(28), ZN => n5095);
   U27 : INV_X1 port map( A => PC_IN(6), ZN => n5229);
   U28 : INV_X1 port map( A => PC_IN(3), ZN => n5233);
   U29 : AND2_X2 port map( A1 => n5236, A2 => IR_FAIL(15), ZN => n5);
   U30 : INV_X1 port map( A => PC_FAIL(6), ZN => n5200);
   U31 : NOR2_X1 port map( A1 => PC_FAIL(2), A2 => n5144, ZN => n5206);
   U32 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(30), A3 => IR_IN(31), 
                           ZN => n5135);
   U33 : NAND3_X1 port map( A1 => n5135, A2 => IR_IN(27), A3 => n5095, ZN => 
                           n5284);
   U34 : INV_X1 port map( A => WRONG_PRE, ZN => n5219);
   U35 : NAND2_X1 port map( A1 => RST, A2 => n5219, ZN => n5285);
   U36 : INV_X1 port map( A => n5285, ZN => n5096);
   U37 : NAND2_X1 port map( A1 => n5284, A2 => n5096, ZN => n5224);
   U38 : INV_X1 port map( A => PC_IN(2), ZN => n5232);
   U39 : NOR2_X1 port map( A1 => n5233, A2 => n5232, ZN => n5231);
   U40 : INV_X1 port map( A => PC_IN(5), ZN => n5138);
   U41 : INV_X1 port map( A => PC_IN(4), ZN => n5226);
   U42 : NOR2_X1 port map( A1 => n5138, A2 => n5226, ZN => n5121);
   U43 : NAND2_X1 port map( A1 => n5231, A2 => n5121, ZN => n5230);
   U44 : NOR2_X1 port map( A1 => n5230, A2 => n5229, ZN => n5228);
   U45 : AOI21_X1 port map( B1 => CACHE_mem_31_1_port, B2 => n5228, A => 
                           IR_IN(27), ZN => n5134);
   U46 : NAND2_X1 port map( A1 => PC_IN(5), A2 => n5226, ZN => n5123);
   U47 : INV_X1 port map( A => CACHE_mem_27_1_port, ZN => n5186);
   U48 : NOR2_X1 port map( A1 => PC_IN(5), A2 => PC_IN(4), ZN => n5126);
   U49 : NOR2_X1 port map( A1 => PC_IN(5), A2 => n5226, ZN => n5120);
   U50 : AOI22_X1 port map( A1 => CACHE_mem_19_1_port, A2 => n5126, B1 => 
                           CACHE_mem_23_1_port, B2 => n5120, ZN => n5097);
   U51 : OAI211_X1 port map( C1 => n5123, C2 => n5186, A => PC_IN(6), B => 
                           n5097, ZN => n5132);
   U52 : INV_X1 port map( A => n5231, ZN => n5227);
   U53 : INV_X1 port map( A => CACHE_mem_11_1_port, ZN => n5099);
   U54 : AOI22_X1 port map( A1 => CACHE_mem_3_1_port, A2 => n5126, B1 => 
                           CACHE_mem_7_1_port, B2 => n5120, ZN => n5098);
   U55 : OAI211_X1 port map( C1 => n5099, C2 => n5123, A => n5098, B => n5229, 
                           ZN => n5100);
   U56 : AOI21_X1 port map( B1 => CACHE_mem_15_1_port, B2 => n5121, A => n5100,
                           ZN => n5101);
   U57 : NOR2_X1 port map( A1 => n5227, A2 => n5101, ZN => n5131);
   U58 : AOI22_X1 port map( A1 => n5121, A2 => CACHE_mem_30_1_port, B1 => 
                           CACHE_mem_22_1_port, B2 => n5120, ZN => n5103);
   U59 : INV_X1 port map( A => n5123, ZN => n5110);
   U60 : AOI22_X1 port map( A1 => CACHE_mem_26_1_port, A2 => n5110, B1 => 
                           CACHE_mem_18_1_port, B2 => n5126, ZN => n5102);
   U61 : AOI21_X1 port map( B1 => n5103, B2 => n5102, A => n5233, ZN => n5107);
   U62 : AOI22_X1 port map( A1 => n5121, A2 => CACHE_mem_28_1_port, B1 => 
                           CACHE_mem_20_1_port, B2 => n5120, ZN => n5105);
   U63 : AOI22_X1 port map( A1 => CACHE_mem_24_1_port, A2 => n5110, B1 => 
                           CACHE_mem_16_1_port, B2 => n5126, ZN => n5104);
   U64 : AOI21_X1 port map( B1 => n5105, B2 => n5104, A => PC_IN(3), ZN => 
                           n5106);
   U65 : OAI21_X1 port map( B1 => n5107, B2 => n5106, A => PC_IN(6), ZN => 
                           n5116);
   U66 : AOI22_X1 port map( A1 => n5121, A2 => CACHE_mem_14_1_port, B1 => 
                           CACHE_mem_6_1_port, B2 => n5120, ZN => n5109);
   U67 : AOI22_X1 port map( A1 => CACHE_mem_10_1_port, A2 => n5110, B1 => 
                           CACHE_mem_2_1_port, B2 => n5126, ZN => n5108);
   U68 : AOI21_X1 port map( B1 => n5109, B2 => n5108, A => n5233, ZN => n5114);
   U69 : AOI22_X1 port map( A1 => n5121, A2 => CACHE_mem_12_1_port, B1 => 
                           CACHE_mem_4_1_port, B2 => n5120, ZN => n5112);
   U70 : AOI22_X1 port map( A1 => CACHE_mem_8_1_port, A2 => n5110, B1 => 
                           CACHE_mem_0_1_port, B2 => n5126, ZN => n5111);
   U71 : AOI21_X1 port map( B1 => n5112, B2 => n5111, A => PC_IN(3), ZN => 
                           n5113);
   U72 : OAI21_X1 port map( B1 => n5114, B2 => n5113, A => n5229, ZN => n5115);
   U73 : AOI21_X1 port map( B1 => n5116, B2 => n5115, A => PC_IN(2), ZN => 
                           n5130);
   U74 : INV_X1 port map( A => CACHE_mem_25_1_port, ZN => n5118);
   U75 : AOI22_X1 port map( A1 => n5121, A2 => CACHE_mem_29_1_port, B1 => 
                           CACHE_mem_21_1_port, B2 => n5120, ZN => n5117);
   U76 : OAI211_X1 port map( C1 => n5123, C2 => n5118, A => PC_IN(6), B => 
                           n5117, ZN => n5119);
   U77 : AOI21_X1 port map( B1 => CACHE_mem_17_1_port, B2 => n5126, A => n5119,
                           ZN => n5128);
   U78 : INV_X1 port map( A => CACHE_mem_9_1_port, ZN => n5124);
   U79 : AOI22_X1 port map( A1 => n5121, A2 => CACHE_mem_13_1_port, B1 => 
                           CACHE_mem_5_1_port, B2 => n5120, ZN => n5122);
   U80 : OAI211_X1 port map( C1 => n5124, C2 => n5123, A => n5122, B => n5229, 
                           ZN => n5125);
   U81 : AOI21_X1 port map( B1 => CACHE_mem_1_1_port, B2 => n5126, A => n5125, 
                           ZN => n5127);
   U82 : NOR4_X1 port map( A1 => PC_IN(3), A2 => n5128, A3 => n5127, A4 => 
                           n5232, ZN => n5129);
   U83 : AOI211_X1 port map( C1 => n5132, C2 => n5131, A => n5130, B => n5129, 
                           ZN => n5133);
   U84 : NAND4_X1 port map( A1 => n5135, A2 => IR_IN(28), A3 => n5134, A4 => 
                           n5133, ZN => n5225);
   U85 : OAI21_X1 port map( B1 => WRONG_PRE, B2 => n5284, A => RST, ZN => N356)
                           ;
   U86 : AND2_X1 port map( A1 => RST, A2 => PC_IN(0), ZN => N357);
   U87 : AND2_X1 port map( A1 => RST, A2 => PC_IN(1), ZN => N358);
   U88 : NAND2_X1 port map( A1 => n5231, A2 => PC_IN(4), ZN => n5137);
   U89 : INV_X1 port map( A => n5230, ZN => n5136);
   U90 : AOI211_X1 port map( C1 => n5138, C2 => n5137, A => n5136, B => n5094, 
                           ZN => N362);
   U91 : INV_X1 port map( A => n5228, ZN => n5250);
   U92 : INV_X1 port map( A => PC_IN(7), ZN => n5249);
   U93 : NOR2_X1 port map( A1 => n5250, A2 => n5249, ZN => n5248);
   U94 : NAND2_X1 port map( A1 => n5248, A2 => PC_IN(8), ZN => n5253);
   U95 : INV_X1 port map( A => PC_IN(9), ZN => n5252);
   U96 : NOR2_X1 port map( A1 => n5253, A2 => n5252, ZN => n5251);
   U97 : NAND2_X1 port map( A1 => n5251, A2 => PC_IN(10), ZN => n5256);
   U98 : INV_X1 port map( A => PC_IN(11), ZN => n5255);
   U99 : NOR2_X1 port map( A1 => n5256, A2 => n5255, ZN => n5254);
   U100 : NAND2_X1 port map( A1 => n5254, A2 => PC_IN(12), ZN => n5259);
   U101 : INV_X1 port map( A => PC_IN(13), ZN => n5258);
   U102 : NOR2_X1 port map( A1 => n5259, A2 => n5258, ZN => n5257);
   U103 : NAND2_X1 port map( A1 => n5257, A2 => PC_IN(14), ZN => n5262);
   U104 : INV_X1 port map( A => PC_IN(15), ZN => n5261);
   U105 : NOR2_X1 port map( A1 => n5262, A2 => n5261, ZN => n5260);
   U106 : NAND2_X1 port map( A1 => n5260, A2 => PC_IN(16), ZN => n5265);
   U107 : INV_X1 port map( A => PC_IN(17), ZN => n5264);
   U108 : NOR2_X1 port map( A1 => n5265, A2 => n5264, ZN => n5263);
   U109 : NAND2_X1 port map( A1 => n5263, A2 => PC_IN(18), ZN => n5268);
   U110 : INV_X1 port map( A => PC_IN(19), ZN => n5267);
   U111 : NOR2_X1 port map( A1 => n5268, A2 => n5267, ZN => n5266);
   U112 : NAND2_X1 port map( A1 => n5266, A2 => PC_IN(20), ZN => n5271);
   U113 : INV_X1 port map( A => PC_IN(21), ZN => n5270);
   U114 : NOR2_X1 port map( A1 => n5271, A2 => n5270, ZN => n5269);
   U115 : NAND2_X1 port map( A1 => n5269, A2 => PC_IN(22), ZN => n5274);
   U116 : INV_X1 port map( A => PC_IN(23), ZN => n5273);
   U117 : NOR2_X1 port map( A1 => n5274, A2 => n5273, ZN => n5272);
   U118 : NAND2_X1 port map( A1 => n5272, A2 => PC_IN(24), ZN => n5277);
   U119 : INV_X1 port map( A => PC_IN(25), ZN => n5276);
   U120 : NOR2_X1 port map( A1 => n5277, A2 => n5276, ZN => n5275);
   U121 : NAND2_X1 port map( A1 => n5275, A2 => PC_IN(26), ZN => n5280);
   U122 : INV_X1 port map( A => PC_IN(27), ZN => n5279);
   U123 : NOR2_X1 port map( A1 => n5280, A2 => n5279, ZN => n5278);
   U124 : NAND2_X1 port map( A1 => n5278, A2 => PC_IN(28), ZN => n5283);
   U125 : INV_X1 port map( A => PC_IN(29), ZN => n5282);
   U126 : NOR2_X1 port map( A1 => n5283, A2 => n5282, ZN => n5281);
   U127 : INV_X1 port map( A => n5281, ZN => n5140);
   U128 : INV_X1 port map( A => PC_IN(30), ZN => n5139);
   U129 : NOR2_X1 port map( A1 => n5140, A2 => n5139, ZN => n5142);
   U130 : AOI211_X1 port map( C1 => n5140, C2 => n5139, A => n5142, B => n5093,
                           ZN => N387);
   U131 : OAI21_X1 port map( B1 => PC_IN(31), B2 => n5142, A => RST, ZN => 
                           n5141);
   U132 : AOI21_X1 port map( B1 => PC_IN(31), B2 => n5142, A => n5141, ZN => 
                           N388);
   U133 : NAND3_X1 port map( A1 => PC_FAIL(2), A2 => PC_FAIL(4), A3 => 
                           PC_FAIL(3), ZN => n5174);
   U134 : INV_X1 port map( A => PC_FAIL(2), ZN => n5143);
   U135 : INV_X1 port map( A => PC_FAIL(3), ZN => n5145);
   U136 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_9_0_port, B1 => n5202
                           , B2 => CACHE_mem_10_0_port, ZN => n5155);
   U137 : NAND3_X1 port map( A1 => n5143, A2 => n5145, A3 => PC_FAIL(4), ZN => 
                           n5177);
   U138 : INV_X1 port map( A => n5177, ZN => n5204);
   U139 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_11_0_port, B1 => 
                           n5204, B2 => CACHE_mem_12_0_port, ZN => n5148);
   U140 : NAND2_X1 port map( A1 => PC_FAIL(4), A2 => PC_FAIL(3), ZN => n5144);
   U141 : AOI22_X1 port map( A1 => n5207, A2 => CACHE_mem_8_0_port, B1 => n5206
                           , B2 => CACHE_mem_14_0_port, ZN => n5147);
   U142 : INV_X1 port map( A => n5174, ZN => n5198);
   U143 : NAND3_X1 port map( A1 => n5145, A2 => PC_FAIL(4), A3 => PC_FAIL(2), 
                           ZN => n5176);
   U144 : INV_X1 port map( A => n5176, ZN => n5197);
   U145 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_15_0_port, B1 => 
                           n5197, B2 => CACHE_mem_13_0_port, ZN => n5146);
   U146 : AND4_X1 port map( A1 => PC_FAIL(5), A2 => n5148, A3 => n5147, A4 => 
                           n5146, ZN => n5154);
   U147 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_1_0_port, B1 => n5202
                           , B2 => CACHE_mem_2_0_port, ZN => n5153);
   U148 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_3_0_port, B1 => n5204
                           , B2 => CACHE_mem_4_0_port, ZN => n5151);
   U149 : AOI22_X1 port map( A1 => n5207, A2 => CACHE_mem_0_0_port, B1 => n5206
                           , B2 => CACHE_mem_6_0_port, ZN => n5150);
   U150 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_7_0_port, B1 => n5197
                           , B2 => CACHE_mem_5_0_port, ZN => n5149);
   U151 : AND4_X1 port map( A1 => n5151, A2 => n5150, A3 => n5149, A4 => n5199,
                           ZN => n5152);
   U152 : AOI22_X1 port map( A1 => n5155, A2 => n5154, B1 => n5153, B2 => n5152
                           , ZN => n5167);
   U153 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_25_0_port, B1 => 
                           n5202, B2 => CACHE_mem_26_0_port, ZN => n5165);
   U154 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_27_0_port, B1 => 
                           n5204, B2 => CACHE_mem_28_0_port, ZN => n5158);
   U155 : AOI22_X1 port map( A1 => n5207, A2 => CACHE_mem_24_0_port, B1 => 
                           n5206, B2 => CACHE_mem_30_0_port, ZN => n5157);
   U156 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_31_0_port, B1 => 
                           n5197, B2 => CACHE_mem_29_0_port, ZN => n5156);
   U157 : AND4_X1 port map( A1 => PC_FAIL(5), A2 => n5158, A3 => n5157, A4 => 
                           n5156, ZN => n5164);
   U158 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_17_0_port, B1 => 
                           n5202, B2 => CACHE_mem_18_0_port, ZN => n5163);
   U159 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_19_0_port, B1 => 
                           n5204, B2 => CACHE_mem_20_0_port, ZN => n5161);
   U160 : AOI22_X1 port map( A1 => n5207, A2 => CACHE_mem_16_0_port, B1 => 
                           n5206, B2 => CACHE_mem_22_0_port, ZN => n5160);
   U161 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_23_0_port, B1 => 
                           n5197, B2 => CACHE_mem_21_0_port, ZN => n5159);
   U162 : AND4_X1 port map( A1 => n5161, A2 => n5160, A3 => n5159, A4 => n5199,
                           ZN => n5162);
   U163 : AOI22_X1 port map( A1 => n5165, A2 => n5164, B1 => n5163, B2 => n5162
                           , ZN => n5166);
   U164 : MUX2_X1 port map( A => n5167, B => n5166, S => PC_FAIL(6), Z => n5222
                           );
   U165 : AOI21_X1 port map( B1 => n5222, B2 => RIGHT_PRE, A => n5089, ZN => 
                           n5169);
   U166 : NOR2_X1 port map( A1 => n5169, A2 => n5199, ZN => n5171);
   U167 : NAND2_X1 port map( A1 => PC_FAIL(6), A2 => n5171, ZN => n5168);
   U168 : OAI21_X1 port map( B1 => n5174, B2 => n5168, A => RST, ZN => N612);
   U169 : INV_X1 port map( A => n5206, ZN => n5175);
   U170 : OAI21_X1 port map( B1 => n5175, B2 => n5168, A => RST, ZN => N613);
   U171 : OAI21_X1 port map( B1 => n5176, B2 => n5168, A => RST, ZN => N614);
   U172 : OAI21_X1 port map( B1 => n5177, B2 => n5168, A => RST, ZN => N615);
   U173 : OAI21_X1 port map( B1 => n5187, B2 => n5168, A => RST, ZN => N616);
   U174 : OAI21_X1 port map( B1 => n5178, B2 => n5168, A => RST, ZN => N617);
   U175 : OAI21_X1 port map( B1 => n5179, B2 => n5168, A => RST, ZN => N618);
   U176 : OAI21_X1 port map( B1 => n5181, B2 => n5168, A => RST, ZN => N619);
   U177 : NOR2_X1 port map( A1 => PC_FAIL(5), A2 => n5169, ZN => n5173);
   U178 : NAND2_X1 port map( A1 => PC_FAIL(6), A2 => n5173, ZN => n5170);
   U179 : OAI21_X1 port map( B1 => n5174, B2 => n5170, A => RST, ZN => N620);
   U180 : OAI21_X1 port map( B1 => n5175, B2 => n5170, A => RST, ZN => N621);
   U181 : OAI21_X1 port map( B1 => n5176, B2 => n5170, A => RST, ZN => N622);
   U182 : OAI21_X1 port map( B1 => n5177, B2 => n5170, A => RST, ZN => N623);
   U183 : OAI21_X1 port map( B1 => n5187, B2 => n5170, A => RST, ZN => N624);
   U184 : OAI21_X1 port map( B1 => n5178, B2 => n5170, A => RST, ZN => N625);
   U185 : OAI21_X1 port map( B1 => n5179, B2 => n5170, A => RST, ZN => N626);
   U186 : OAI21_X1 port map( B1 => n5181, B2 => n5170, A => RST, ZN => N627);
   U187 : NAND2_X1 port map( A1 => n5171, A2 => n5200, ZN => n5172);
   U188 : OAI21_X1 port map( B1 => n5174, B2 => n5172, A => RST, ZN => N628);
   U189 : OAI21_X1 port map( B1 => n5175, B2 => n5172, A => RST, ZN => N629);
   U190 : OAI21_X1 port map( B1 => n5176, B2 => n5172, A => RST, ZN => N630);
   U191 : OAI21_X1 port map( B1 => n5177, B2 => n5172, A => RST, ZN => N631);
   U192 : OAI21_X1 port map( B1 => n5187, B2 => n5172, A => RST, ZN => N632);
   U193 : OAI21_X1 port map( B1 => n5178, B2 => n5172, A => RST, ZN => N633);
   U194 : OAI21_X1 port map( B1 => n5179, B2 => n5172, A => RST, ZN => N634);
   U195 : OAI21_X1 port map( B1 => n5181, B2 => n5172, A => RST, ZN => N635);
   U196 : NAND2_X1 port map( A1 => n5173, A2 => n5200, ZN => n5180);
   U197 : OAI21_X1 port map( B1 => n5174, B2 => n5180, A => RST, ZN => N636);
   U198 : OAI21_X1 port map( B1 => n5175, B2 => n5180, A => RST, ZN => N637);
   U199 : OAI21_X1 port map( B1 => n5176, B2 => n5180, A => RST, ZN => N638);
   U200 : OAI21_X1 port map( B1 => n5177, B2 => n5180, A => RST, ZN => N639);
   U201 : OAI21_X1 port map( B1 => n5187, B2 => n5180, A => RST, ZN => N640);
   U202 : OAI21_X1 port map( B1 => n5178, B2 => n5180, A => RST, ZN => N641);
   U203 : OAI21_X1 port map( B1 => n5179, B2 => n5180, A => RST, ZN => N642);
   U204 : OAI21_X1 port map( B1 => n5181, B2 => n5180, A => RST, ZN => N643);
   U205 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_9_1_port, B1 => n5202
                           , B2 => CACHE_mem_10_1_port, ZN => n5218);
   U206 : NOR2_X1 port map( A1 => PC_FAIL(6), A2 => n5199, ZN => n5185);
   U207 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_11_1_port, B1 => 
                           n5206, B2 => CACHE_mem_14_1_port, ZN => n5184);
   U208 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_15_1_port, B1 => 
                           n5207, B2 => CACHE_mem_8_1_port, ZN => n5183);
   U209 : AOI22_X1 port map( A1 => n5204, A2 => CACHE_mem_12_1_port, B1 => 
                           n5197, B2 => CACHE_mem_13_1_port, ZN => n5182);
   U210 : AND4_X1 port map( A1 => n5185, A2 => n5184, A3 => n5183, A4 => n5182,
                           ZN => n5217);
   U211 : OAI211_X1 port map( C1 => n5187, C2 => n5186, A => PC_FAIL(5), B => 
                           PC_FAIL(6), ZN => n5192);
   U212 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_25_1_port, B1 => 
                           n5207, B2 => CACHE_mem_24_1_port, ZN => n5190);
   U213 : AOI22_X1 port map( A1 => n5204, A2 => CACHE_mem_28_1_port, B1 => 
                           n5206, B2 => CACHE_mem_30_1_port, ZN => n5189);
   U214 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_31_1_port, B1 => 
                           n5197, B2 => CACHE_mem_29_1_port, ZN => n5188);
   U215 : NAND3_X1 port map( A1 => n5190, A2 => n5189, A3 => n5188, ZN => n5191
                           );
   U216 : AOI22_X1 port map( A1 => n5202, A2 => CACHE_mem_18_1_port, B1 => 
                           n5207, B2 => CACHE_mem_16_1_port, ZN => n5193);
   U217 : NAND3_X1 port map( A1 => PC_FAIL(6), A2 => n5193, A3 => n5199, ZN => 
                           n5214);
   U218 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_17_1_port, B1 => 
                           n5197, B2 => CACHE_mem_21_1_port, ZN => n5196);
   U219 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_19_1_port, B1 => 
                           n5204, B2 => CACHE_mem_20_1_port, ZN => n5195);
   U220 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_23_1_port, B1 => 
                           n5206, B2 => CACHE_mem_22_1_port, ZN => n5194);
   U221 : NAND3_X1 port map( A1 => n5196, A2 => n5195, A3 => n5194, ZN => n5213
                           );
   U222 : AOI22_X1 port map( A1 => n5198, A2 => CACHE_mem_7_1_port, B1 => n5197
                           , B2 => CACHE_mem_5_1_port, ZN => n5201);
   U223 : NAND3_X1 port map( A1 => n5201, A2 => n5200, A3 => n5199, ZN => n5212
                           );
   U224 : AOI22_X1 port map( A1 => n5203, A2 => CACHE_mem_1_1_port, B1 => n5202
                           , B2 => CACHE_mem_2_1_port, ZN => n5210);
   U225 : AOI22_X1 port map( A1 => n5205, A2 => CACHE_mem_3_1_port, B1 => n5204
                           , B2 => CACHE_mem_4_1_port, ZN => n5209);
   U226 : AOI22_X1 port map( A1 => n5207, A2 => CACHE_mem_0_1_port, B1 => n5206
                           , B2 => CACHE_mem_6_1_port, ZN => n5208);
   U227 : NAND3_X1 port map( A1 => n5210, A2 => n5209, A3 => n5208, ZN => n5211
                           );
   U228 : OAI22_X1 port map( A1 => n5214, A2 => n5213, B1 => n5212, B2 => n5211
                           , ZN => n5215);
   U229 : NOR2_X1 port map( A1 => n5236, A2 => n5219, ZN => n5221);
   U230 : AOI22_X1 port map( A1 => n5236, A2 => n5219, B1 => n5222, B2 => n5221
                           , ZN => n5220);
   U231 : OAI21_X1 port map( B1 => n5222, B2 => n5221, A => n5220, ZN => n5223)
                           ;
   U232 : NOR2_X1 port map( A1 => n5225, A2 => n5224, ZN => TAKEN);
   U233 : AND3_X1 port map( A1 => n5236, A2 => IR_FAIL(0), A3 => PC_FAIL(0), ZN
                           => add_53_aco_n2);
   U234 : AND2_X1 port map( A1 => PC_IN(0), A2 => IR_IN(0), ZN => add_59_n1);
   U235 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(4), ZN => n10);
   U236 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(6), ZN => n11);
   U237 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(7), ZN => n12);
   U238 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(8), ZN => n13);
   U239 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(9), ZN => n14);
   U240 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(10), ZN => n15);
   U241 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(11), ZN => n16);
   U242 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(12), ZN => n17);
   U243 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(13), ZN => n18);
   U244 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(14), ZN => n19);
   U245 : AOI221_X1 port map( B1 => n5231, B2 => PC_IN(4), C1 => n5227, C2 => 
                           n5226, A => n5094, ZN => n286);
   U246 : AOI211_X1 port map( C1 => n5230, C2 => n5229, A => n5228, B => n5093,
                           ZN => n291);
   U247 : AOI211_X1 port map( C1 => n5233, C2 => n5232, A => n5231, B => n5093,
                           ZN => n59_port);
   U248 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(1), ZN => n6);
   U249 : NOR2_X1 port map( A1 => PC_IN(0), A2 => IR_IN(0), ZN => n5235);
   U250 : AOI21_X1 port map( B1 => IR_FAIL(0), B2 => n5236, A => PC_FAIL(0), ZN
                           => n5234);
   U251 : OAI33_X1 port map( A1 => n5285, A2 => add_59_n1, A3 => n5235, B1 => 
                           n5090, B2 => n5234, B3 => add_53_aco_n2, ZN => 
                           n60_port);
   U252 : NOR2_X1 port map( A1 => PC_IN(2), A2 => n5093, ZN => n62_port);
   U253 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(5), ZN => n7);
   U254 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(2), ZN => n8);
   U255 : AND2_X1 port map( A1 => n5236, A2 => IR_FAIL(3), ZN => n9);
   U256 : OAI211_X1 port map( C1 => n5272, C2 => PC_IN(24), A => n5277, B => 
                           RST, ZN => n5237);
   U257 : INV_X1 port map( A => n5237, ZN => n293);
   U258 : OAI211_X1 port map( C1 => n5254, C2 => PC_IN(12), A => n5259, B => 
                           RST, ZN => n5238);
   U259 : INV_X1 port map( A => n5238, ZN => n292);
   U260 : OAI211_X1 port map( C1 => n5269, C2 => PC_IN(22), A => n5274, B => 
                           RST, ZN => n5239);
   U261 : INV_X1 port map( A => n5239, ZN => n290);
   U262 : OAI211_X1 port map( C1 => n5266, C2 => PC_IN(20), A => n5271, B => 
                           RST, ZN => n5240);
   U263 : INV_X1 port map( A => n5240, ZN => n289);
   U264 : OAI211_X1 port map( C1 => n5263, C2 => PC_IN(18), A => n5268, B => 
                           RST, ZN => n5241);
   U265 : INV_X1 port map( A => n5241, ZN => n288);
   U266 : OAI211_X1 port map( C1 => n5278, C2 => PC_IN(28), A => n5283, B => 
                           RST, ZN => n5242);
   U267 : INV_X1 port map( A => n5242, ZN => n287);
   U268 : OAI211_X1 port map( C1 => n5260, C2 => PC_IN(16), A => n5265, B => 
                           RST, ZN => n5243);
   U269 : INV_X1 port map( A => n5243, ZN => n285);
   U270 : OAI211_X1 port map( C1 => n5257, C2 => PC_IN(14), A => n5262, B => 
                           RST, ZN => n5244);
   U271 : INV_X1 port map( A => n5244, ZN => n284);
   U272 : OAI211_X1 port map( C1 => n5275, C2 => PC_IN(26), A => n5280, B => 
                           RST, ZN => n5245);
   U273 : INV_X1 port map( A => n5245, ZN => n283);
   U274 : OAI211_X1 port map( C1 => n5248, C2 => PC_IN(8), A => n5253, B => RST
                           , ZN => n5246);
   U275 : INV_X1 port map( A => n5246, ZN => n282);
   U276 : OAI211_X1 port map( C1 => n5251, C2 => PC_IN(10), A => n5256, B => 
                           RST, ZN => n5247);
   U277 : INV_X1 port map( A => n5247, ZN => n281);
   U278 : AOI211_X1 port map( C1 => n5250, C2 => n5249, A => n5248, B => n5093,
                           ZN => n61_port);
   U279 : AOI211_X1 port map( C1 => n5253, C2 => n5252, A => n5251, B => n5093,
                           ZN => n58_port);
   U280 : AOI211_X1 port map( C1 => n5256, C2 => n5255, A => n5254, B => n5093,
                           ZN => n57_port);
   U281 : AOI211_X1 port map( C1 => n5259, C2 => n5258, A => n5257, B => n5093,
                           ZN => n56_port);
   U282 : AOI211_X1 port map( C1 => n5262, C2 => n5261, A => n5260, B => n5093,
                           ZN => n55_port);
   U283 : AOI211_X1 port map( C1 => n5265, C2 => n5264, A => n5263, B => n5094,
                           ZN => n54_port);
   U284 : AOI211_X1 port map( C1 => n5268, C2 => n5267, A => n5266, B => n5094,
                           ZN => n53_port);
   U285 : AOI211_X1 port map( C1 => n5271, C2 => n5270, A => n5269, B => n5094,
                           ZN => n52_port);
   U286 : AOI211_X1 port map( C1 => n5274, C2 => n5273, A => n5272, B => n5094,
                           ZN => n51_port);
   U287 : AOI211_X1 port map( C1 => n5277, C2 => n5276, A => n5275, B => n5094,
                           ZN => n50_port);
   U288 : AOI211_X1 port map( C1 => n5280, C2 => n5279, A => n5278, B => n5094,
                           ZN => n49_port);
   U289 : AOI211_X1 port map( C1 => n5283, C2 => n5282, A => n5281, B => n5093,
                           ZN => n48_port);
   U290 : AOI222_X1 port map( A1 => n5089, A2 => N47, B1 => n5317, B2 => N220, 
                           C1 => n5316, C2 => N82, ZN => n5286);
   U291 : INV_X1 port map( A => n5286, ZN => n46);
   U292 : AOI222_X1 port map( A1 => n5089, A2 => N48, B1 => n5317, B2 => N221, 
                           C1 => n5091, C2 => N83, ZN => n5287);
   U293 : INV_X1 port map( A => n5287, ZN => n45);
   U294 : AOI222_X1 port map( A1 => n5089, A2 => N49, B1 => n5317, B2 => N222, 
                           C1 => n5316, C2 => N84, ZN => n5288);
   U295 : INV_X1 port map( A => n5288, ZN => n44);
   U296 : AOI222_X1 port map( A1 => n5089, A2 => N50, B1 => n5317, B2 => N223, 
                           C1 => n5091, C2 => N85, ZN => n5289);
   U297 : INV_X1 port map( A => n5289, ZN => n43);
   U298 : AOI222_X1 port map( A1 => n5089, A2 => N51, B1 => n5317, B2 => N224, 
                           C1 => n5316, C2 => N86, ZN => n5290);
   U299 : INV_X1 port map( A => n5290, ZN => n42);
   U300 : AOI222_X1 port map( A1 => n5089, A2 => N52, B1 => n5317, B2 => N225, 
                           C1 => n5091, C2 => N87, ZN => n5291);
   U301 : INV_X1 port map( A => n5291, ZN => n41);
   U302 : AOI222_X1 port map( A1 => n5089, A2 => N53, B1 => n5317, B2 => N226, 
                           C1 => n5316, C2 => N88, ZN => n5292);
   U303 : INV_X1 port map( A => n5292, ZN => n40);
   U304 : AOI222_X1 port map( A1 => n5089, A2 => N54, B1 => n5317, B2 => N227, 
                           C1 => n5316, C2 => N89, ZN => n5293);
   U305 : INV_X1 port map( A => n5293, ZN => n39);
   U306 : AOI222_X1 port map( A1 => n5089, A2 => N55, B1 => n5317, B2 => N228, 
                           C1 => n5316, C2 => N90, ZN => n5294);
   U307 : INV_X1 port map( A => n5294, ZN => n38);
   U308 : AOI222_X1 port map( A1 => n5089, A2 => N56, B1 => n5317, B2 => N229, 
                           C1 => n5316, C2 => N91, ZN => n5295);
   U309 : INV_X1 port map( A => n5295, ZN => n37);
   U310 : AOI222_X1 port map( A1 => n5089, A2 => N57, B1 => n5317, B2 => N230, 
                           C1 => n5316, C2 => N92, ZN => n5296);
   U311 : INV_X1 port map( A => n5296, ZN => n36);
   U312 : AOI222_X1 port map( A1 => n5089, A2 => N58, B1 => n5317, B2 => N231, 
                           C1 => n5316, C2 => N93, ZN => n5297);
   U313 : INV_X1 port map( A => n5297, ZN => n35);
   U314 : AOI222_X1 port map( A1 => n5089, A2 => N59, B1 => n5317, B2 => N232, 
                           C1 => n5091, C2 => N94, ZN => n5298);
   U315 : INV_X1 port map( A => n5298, ZN => n34);
   U316 : AOI222_X1 port map( A1 => n5089, A2 => N60, B1 => n5317, B2 => N233, 
                           C1 => n5091, C2 => N95, ZN => n5299);
   U317 : INV_X1 port map( A => n5299, ZN => n33);
   U318 : AOI222_X1 port map( A1 => n5089, A2 => N61, B1 => n5317, B2 => N234, 
                           C1 => n5091, C2 => N96, ZN => n5300);
   U319 : INV_X1 port map( A => n5300, ZN => n32);
   U320 : AOI222_X1 port map( A1 => n5089, A2 => N62, B1 => n5317, B2 => N235, 
                           C1 => n5091, C2 => N97, ZN => n5301);
   U321 : INV_X1 port map( A => n5301, ZN => n31);
   U322 : AOI222_X1 port map( A1 => n5089, A2 => N63, B1 => n5317, B2 => N236, 
                           C1 => n5091, C2 => N98, ZN => n5302);
   U323 : INV_X1 port map( A => n5302, ZN => n30);
   U324 : AOI222_X1 port map( A1 => n5089, A2 => N64, B1 => n5317, B2 => N237, 
                           C1 => n5091, C2 => N99, ZN => n5303);
   U325 : INV_X1 port map( A => n5303, ZN => n29);
   U326 : AOI222_X1 port map( A1 => n5089, A2 => N65, B1 => n5317, B2 => N238, 
                           C1 => n5091, C2 => N100, ZN => n5304);
   U327 : INV_X1 port map( A => n5304, ZN => n28);
   U328 : AOI222_X1 port map( A1 => n5089, A2 => N66, B1 => n5317, B2 => N239, 
                           C1 => n5316, C2 => N101, ZN => n5305);
   U329 : INV_X1 port map( A => n5305, ZN => n27);
   U330 : AOI222_X1 port map( A1 => n5089, A2 => N67, B1 => n5317, B2 => N240, 
                           C1 => n5091, C2 => N102, ZN => n5306);
   U331 : INV_X1 port map( A => n5306, ZN => n26);
   U332 : AOI222_X1 port map( A1 => n5089, A2 => N68, B1 => n5317, B2 => N241, 
                           C1 => n5316, C2 => N103, ZN => n5307);
   U333 : INV_X1 port map( A => n5307, ZN => n25);
   U334 : AOI222_X1 port map( A1 => n5089, A2 => N69, B1 => n5317, B2 => N242, 
                           C1 => n5091, C2 => N104, ZN => n5308);
   U335 : INV_X1 port map( A => n5308, ZN => n24);
   U336 : AOI222_X1 port map( A1 => n5089, A2 => N70, B1 => n5317, B2 => N243, 
                           C1 => n5316, C2 => N105, ZN => n5309);
   U337 : INV_X1 port map( A => n5309, ZN => n23);
   U338 : AOI222_X1 port map( A1 => n5089, A2 => N71, B1 => n5317, B2 => N244, 
                           C1 => n5091, C2 => N106, ZN => n5310);
   U339 : INV_X1 port map( A => n5310, ZN => n22);
   U340 : AOI222_X1 port map( A1 => n5089, A2 => N72, B1 => n5317, B2 => N245, 
                           C1 => n5091, C2 => N107, ZN => n5311);
   U341 : INV_X1 port map( A => n5311, ZN => n21);
   U342 : AOI222_X1 port map( A1 => n5089, A2 => N73, B1 => n5317, B2 => N246, 
                           C1 => n5091, C2 => N108, ZN => n5312);
   U343 : INV_X1 port map( A => n5312, ZN => n20);
   U344 : AOI222_X1 port map( A1 => n5089, A2 => N74, B1 => n5317, B2 => N247, 
                           C1 => n5091, C2 => N109, ZN => n5313);
   U345 : INV_X1 port map( A => n5313, ZN => n4);
   U346 : AOI222_X1 port map( A1 => n5089, A2 => N75, B1 => n5317, B2 => N248, 
                           C1 => n5091, C2 => N110, ZN => n5314);
   U347 : INV_X1 port map( A => n5314, ZN => n3);
   U348 : AOI222_X1 port map( A1 => n5089, A2 => N76, B1 => n5317, B2 => N249, 
                           C1 => n5091, C2 => N111, ZN => n5315);
   U349 : INV_X1 port map( A => n5315, ZN => n2);
   U350 : AOI222_X1 port map( A1 => n5089, A2 => N77, B1 => n5317, B2 => N250, 
                           C1 => n5091, C2 => N112, ZN => n5318);
   U351 : INV_X1 port map( A => n5318, ZN => n1);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity register_file_N32_addBit5 is

   port( RESET, RE, WE : in std_logic;  ADD_WR, ADD_RDA, ADD_RDB : in 
         std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUTA, OUTB : out std_logic_vector (31 downto 0));

end register_file_N32_addBit5;

architecture SYN_A of register_file_N32_addBit5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_1_31_port, REGISTERS_1_30_port, REGISTERS_1_29_port, 
      REGISTERS_1_28_port, REGISTERS_1_27_port, REGISTERS_1_26_port, 
      REGISTERS_1_25_port, REGISTERS_1_24_port, REGISTERS_1_23_port, 
      REGISTERS_1_22_port, REGISTERS_1_21_port, REGISTERS_1_20_port, 
      REGISTERS_1_19_port, REGISTERS_1_18_port, REGISTERS_1_17_port, 
      REGISTERS_1_16_port, REGISTERS_1_15_port, REGISTERS_1_14_port, 
      REGISTERS_1_13_port, REGISTERS_1_12_port, REGISTERS_1_11_port, 
      REGISTERS_1_10_port, REGISTERS_1_9_port, REGISTERS_1_8_port, 
      REGISTERS_1_7_port, REGISTERS_1_6_port, REGISTERS_1_5_port, 
      REGISTERS_1_4_port, REGISTERS_1_3_port, REGISTERS_1_2_port, 
      REGISTERS_1_1_port, REGISTERS_1_0_port, REGISTERS_2_31_port, 
      REGISTERS_2_30_port, REGISTERS_2_29_port, REGISTERS_2_28_port, 
      REGISTERS_2_27_port, REGISTERS_2_26_port, REGISTERS_2_25_port, 
      REGISTERS_2_24_port, REGISTERS_2_23_port, REGISTERS_2_22_port, 
      REGISTERS_2_21_port, REGISTERS_2_20_port, REGISTERS_2_19_port, 
      REGISTERS_2_18_port, REGISTERS_2_17_port, REGISTERS_2_16_port, 
      REGISTERS_2_15_port, REGISTERS_2_14_port, REGISTERS_2_13_port, 
      REGISTERS_2_12_port, REGISTERS_2_11_port, REGISTERS_2_10_port, 
      REGISTERS_2_9_port, REGISTERS_2_8_port, REGISTERS_2_7_port, 
      REGISTERS_2_6_port, REGISTERS_2_5_port, REGISTERS_2_4_port, 
      REGISTERS_2_3_port, REGISTERS_2_2_port, REGISTERS_2_1_port, 
      REGISTERS_2_0_port, REGISTERS_3_31_port, REGISTERS_3_30_port, 
      REGISTERS_3_29_port, REGISTERS_3_28_port, REGISTERS_3_27_port, 
      REGISTERS_3_26_port, REGISTERS_3_25_port, REGISTERS_3_24_port, 
      REGISTERS_3_23_port, REGISTERS_3_22_port, REGISTERS_3_21_port, 
      REGISTERS_3_20_port, REGISTERS_3_19_port, REGISTERS_3_18_port, 
      REGISTERS_3_17_port, REGISTERS_3_16_port, REGISTERS_3_15_port, 
      REGISTERS_3_14_port, REGISTERS_3_13_port, REGISTERS_3_12_port, 
      REGISTERS_3_11_port, REGISTERS_3_10_port, REGISTERS_3_9_port, 
      REGISTERS_3_8_port, REGISTERS_3_7_port, REGISTERS_3_6_port, 
      REGISTERS_3_5_port, REGISTERS_3_4_port, REGISTERS_3_3_port, 
      REGISTERS_3_2_port, REGISTERS_3_1_port, REGISTERS_3_0_port, 
      REGISTERS_4_31_port, REGISTERS_4_30_port, REGISTERS_4_29_port, 
      REGISTERS_4_28_port, REGISTERS_4_27_port, REGISTERS_4_26_port, 
      REGISTERS_4_25_port, REGISTERS_4_24_port, REGISTERS_4_23_port, 
      REGISTERS_4_22_port, REGISTERS_4_21_port, REGISTERS_4_20_port, 
      REGISTERS_4_19_port, REGISTERS_4_18_port, REGISTERS_4_17_port, 
      REGISTERS_4_16_port, REGISTERS_4_15_port, REGISTERS_4_14_port, 
      REGISTERS_4_13_port, REGISTERS_4_12_port, REGISTERS_4_11_port, 
      REGISTERS_4_10_port, REGISTERS_4_9_port, REGISTERS_4_8_port, 
      REGISTERS_4_7_port, REGISTERS_4_6_port, REGISTERS_4_5_port, 
      REGISTERS_4_4_port, REGISTERS_4_3_port, REGISTERS_4_2_port, 
      REGISTERS_4_1_port, REGISTERS_4_0_port, REGISTERS_5_31_port, 
      REGISTERS_5_30_port, REGISTERS_5_29_port, REGISTERS_5_28_port, 
      REGISTERS_5_27_port, REGISTERS_5_26_port, REGISTERS_5_25_port, 
      REGISTERS_5_24_port, REGISTERS_5_23_port, REGISTERS_5_22_port, 
      REGISTERS_5_21_port, REGISTERS_5_20_port, REGISTERS_5_19_port, 
      REGISTERS_5_18_port, REGISTERS_5_17_port, REGISTERS_5_16_port, 
      REGISTERS_5_15_port, REGISTERS_5_14_port, REGISTERS_5_13_port, 
      REGISTERS_5_12_port, REGISTERS_5_11_port, REGISTERS_5_10_port, 
      REGISTERS_5_9_port, REGISTERS_5_8_port, REGISTERS_5_7_port, 
      REGISTERS_5_6_port, REGISTERS_5_5_port, REGISTERS_5_4_port, 
      REGISTERS_5_3_port, REGISTERS_5_2_port, REGISTERS_5_1_port, 
      REGISTERS_5_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_8_31_port, 
      REGISTERS_8_30_port, REGISTERS_8_29_port, REGISTERS_8_28_port, 
      REGISTERS_8_27_port, REGISTERS_8_26_port, REGISTERS_8_25_port, 
      REGISTERS_8_24_port, REGISTERS_8_23_port, REGISTERS_8_22_port, 
      REGISTERS_8_21_port, REGISTERS_8_20_port, REGISTERS_8_19_port, 
      REGISTERS_8_18_port, REGISTERS_8_17_port, REGISTERS_8_16_port, 
      REGISTERS_8_15_port, REGISTERS_8_14_port, REGISTERS_8_13_port, 
      REGISTERS_8_12_port, REGISTERS_8_11_port, REGISTERS_8_10_port, 
      REGISTERS_8_9_port, REGISTERS_8_8_port, REGISTERS_8_7_port, 
      REGISTERS_8_6_port, REGISTERS_8_5_port, REGISTERS_8_4_port, 
      REGISTERS_8_3_port, REGISTERS_8_2_port, REGISTERS_8_1_port, 
      REGISTERS_8_0_port, REGISTERS_9_31_port, REGISTERS_9_30_port, 
      REGISTERS_9_29_port, REGISTERS_9_28_port, REGISTERS_9_27_port, 
      REGISTERS_9_26_port, REGISTERS_9_25_port, REGISTERS_9_24_port, 
      REGISTERS_9_23_port, REGISTERS_9_22_port, REGISTERS_9_21_port, 
      REGISTERS_9_20_port, REGISTERS_9_19_port, REGISTERS_9_18_port, 
      REGISTERS_9_17_port, REGISTERS_9_16_port, REGISTERS_9_15_port, 
      REGISTERS_9_14_port, REGISTERS_9_13_port, REGISTERS_9_12_port, 
      REGISTERS_9_11_port, REGISTERS_9_10_port, REGISTERS_9_9_port, 
      REGISTERS_9_8_port, REGISTERS_9_7_port, REGISTERS_9_6_port, 
      REGISTERS_9_5_port, REGISTERS_9_4_port, REGISTERS_9_3_port, 
      REGISTERS_9_2_port, REGISTERS_9_1_port, REGISTERS_9_0_port, 
      REGISTERS_10_31_port, REGISTERS_10_30_port, REGISTERS_10_29_port, 
      REGISTERS_10_28_port, REGISTERS_10_27_port, REGISTERS_10_26_port, 
      REGISTERS_10_25_port, REGISTERS_10_24_port, REGISTERS_10_23_port, 
      REGISTERS_10_22_port, REGISTERS_10_21_port, REGISTERS_10_20_port, 
      REGISTERS_10_19_port, REGISTERS_10_18_port, REGISTERS_10_17_port, 
      REGISTERS_10_16_port, REGISTERS_10_15_port, REGISTERS_10_14_port, 
      REGISTERS_10_13_port, REGISTERS_10_12_port, REGISTERS_10_11_port, 
      REGISTERS_10_10_port, REGISTERS_10_9_port, REGISTERS_10_8_port, 
      REGISTERS_10_7_port, REGISTERS_10_6_port, REGISTERS_10_5_port, 
      REGISTERS_10_4_port, REGISTERS_10_3_port, REGISTERS_10_2_port, 
      REGISTERS_10_1_port, REGISTERS_10_0_port, REGISTERS_11_31_port, 
      REGISTERS_11_30_port, REGISTERS_11_29_port, REGISTERS_11_28_port, 
      REGISTERS_11_27_port, REGISTERS_11_26_port, REGISTERS_11_25_port, 
      REGISTERS_11_24_port, REGISTERS_11_23_port, REGISTERS_11_22_port, 
      REGISTERS_11_21_port, REGISTERS_11_20_port, REGISTERS_11_19_port, 
      REGISTERS_11_18_port, REGISTERS_11_17_port, REGISTERS_11_16_port, 
      REGISTERS_11_15_port, REGISTERS_11_14_port, REGISTERS_11_13_port, 
      REGISTERS_11_12_port, REGISTERS_11_11_port, REGISTERS_11_10_port, 
      REGISTERS_11_9_port, REGISTERS_11_8_port, REGISTERS_11_7_port, 
      REGISTERS_11_6_port, REGISTERS_11_5_port, REGISTERS_11_4_port, 
      REGISTERS_11_3_port, REGISTERS_11_2_port, REGISTERS_11_1_port, 
      REGISTERS_11_0_port, REGISTERS_12_31_port, REGISTERS_12_30_port, 
      REGISTERS_12_29_port, REGISTERS_12_28_port, REGISTERS_12_27_port, 
      REGISTERS_12_26_port, REGISTERS_12_25_port, REGISTERS_12_24_port, 
      REGISTERS_12_23_port, REGISTERS_12_22_port, REGISTERS_12_21_port, 
      REGISTERS_12_20_port, REGISTERS_12_19_port, REGISTERS_12_18_port, 
      REGISTERS_12_17_port, REGISTERS_12_16_port, REGISTERS_12_15_port, 
      REGISTERS_12_14_port, REGISTERS_12_13_port, REGISTERS_12_12_port, 
      REGISTERS_12_11_port, REGISTERS_12_10_port, REGISTERS_12_9_port, 
      REGISTERS_12_8_port, REGISTERS_12_7_port, REGISTERS_12_6_port, 
      REGISTERS_12_5_port, REGISTERS_12_4_port, REGISTERS_12_3_port, 
      REGISTERS_12_2_port, REGISTERS_12_1_port, REGISTERS_12_0_port, 
      REGISTERS_13_31_port, REGISTERS_13_30_port, REGISTERS_13_29_port, 
      REGISTERS_13_28_port, REGISTERS_13_27_port, REGISTERS_13_26_port, 
      REGISTERS_13_25_port, REGISTERS_13_24_port, REGISTERS_13_23_port, 
      REGISTERS_13_22_port, REGISTERS_13_21_port, REGISTERS_13_20_port, 
      REGISTERS_13_19_port, REGISTERS_13_18_port, REGISTERS_13_17_port, 
      REGISTERS_13_16_port, REGISTERS_13_15_port, REGISTERS_13_14_port, 
      REGISTERS_13_13_port, REGISTERS_13_12_port, REGISTERS_13_11_port, 
      REGISTERS_13_10_port, REGISTERS_13_9_port, REGISTERS_13_8_port, 
      REGISTERS_13_7_port, REGISTERS_13_6_port, REGISTERS_13_5_port, 
      REGISTERS_13_4_port, REGISTERS_13_3_port, REGISTERS_13_2_port, 
      REGISTERS_13_1_port, REGISTERS_13_0_port, REGISTERS_14_31_port, 
      REGISTERS_14_30_port, REGISTERS_14_29_port, REGISTERS_14_28_port, 
      REGISTERS_14_27_port, REGISTERS_14_26_port, REGISTERS_14_25_port, 
      REGISTERS_14_24_port, REGISTERS_14_23_port, REGISTERS_14_22_port, 
      REGISTERS_14_21_port, REGISTERS_14_20_port, REGISTERS_14_19_port, 
      REGISTERS_14_18_port, REGISTERS_14_17_port, REGISTERS_14_16_port, 
      REGISTERS_14_15_port, REGISTERS_14_14_port, REGISTERS_14_13_port, 
      REGISTERS_14_12_port, REGISTERS_14_11_port, REGISTERS_14_10_port, 
      REGISTERS_14_9_port, REGISTERS_14_8_port, REGISTERS_14_7_port, 
      REGISTERS_14_6_port, REGISTERS_14_5_port, REGISTERS_14_4_port, 
      REGISTERS_14_3_port, REGISTERS_14_2_port, REGISTERS_14_1_port, 
      REGISTERS_14_0_port, REGISTERS_15_31_port, REGISTERS_15_30_port, 
      REGISTERS_15_29_port, REGISTERS_15_28_port, REGISTERS_15_27_port, 
      REGISTERS_15_26_port, REGISTERS_15_25_port, REGISTERS_15_24_port, 
      REGISTERS_15_23_port, REGISTERS_15_22_port, REGISTERS_15_21_port, 
      REGISTERS_15_20_port, REGISTERS_15_19_port, REGISTERS_15_18_port, 
      REGISTERS_15_17_port, REGISTERS_15_16_port, REGISTERS_15_15_port, 
      REGISTERS_15_14_port, REGISTERS_15_13_port, REGISTERS_15_12_port, 
      REGISTERS_15_11_port, REGISTERS_15_10_port, REGISTERS_15_9_port, 
      REGISTERS_15_8_port, REGISTERS_15_7_port, REGISTERS_15_6_port, 
      REGISTERS_15_5_port, REGISTERS_15_4_port, REGISTERS_15_3_port, 
      REGISTERS_15_2_port, REGISTERS_15_1_port, REGISTERS_15_0_port, 
      REGISTERS_16_31_port, REGISTERS_16_30_port, REGISTERS_16_29_port, 
      REGISTERS_16_28_port, REGISTERS_16_27_port, REGISTERS_16_26_port, 
      REGISTERS_16_25_port, REGISTERS_16_24_port, REGISTERS_16_23_port, 
      REGISTERS_16_22_port, REGISTERS_16_21_port, REGISTERS_16_20_port, 
      REGISTERS_16_19_port, REGISTERS_16_18_port, REGISTERS_16_17_port, 
      REGISTERS_16_16_port, REGISTERS_16_15_port, REGISTERS_16_14_port, 
      REGISTERS_16_13_port, REGISTERS_16_12_port, REGISTERS_16_11_port, 
      REGISTERS_16_10_port, REGISTERS_16_9_port, REGISTERS_16_8_port, 
      REGISTERS_16_7_port, REGISTERS_16_6_port, REGISTERS_16_5_port, 
      REGISTERS_16_4_port, REGISTERS_16_3_port, REGISTERS_16_2_port, 
      REGISTERS_16_1_port, REGISTERS_16_0_port, REGISTERS_17_31_port, 
      REGISTERS_17_30_port, REGISTERS_17_29_port, REGISTERS_17_28_port, 
      REGISTERS_17_27_port, REGISTERS_17_26_port, REGISTERS_17_25_port, 
      REGISTERS_17_24_port, REGISTERS_17_23_port, REGISTERS_17_22_port, 
      REGISTERS_17_21_port, REGISTERS_17_20_port, REGISTERS_17_19_port, 
      REGISTERS_17_18_port, REGISTERS_17_17_port, REGISTERS_17_16_port, 
      REGISTERS_17_15_port, REGISTERS_17_14_port, REGISTERS_17_13_port, 
      REGISTERS_17_12_port, REGISTERS_17_11_port, REGISTERS_17_10_port, 
      REGISTERS_17_9_port, REGISTERS_17_8_port, REGISTERS_17_7_port, 
      REGISTERS_17_6_port, REGISTERS_17_5_port, REGISTERS_17_4_port, 
      REGISTERS_17_3_port, REGISTERS_17_2_port, REGISTERS_17_1_port, 
      REGISTERS_17_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_20_31_port, 
      REGISTERS_20_30_port, REGISTERS_20_29_port, REGISTERS_20_28_port, 
      REGISTERS_20_27_port, REGISTERS_20_26_port, REGISTERS_20_25_port, 
      REGISTERS_20_24_port, REGISTERS_20_23_port, REGISTERS_20_22_port, 
      REGISTERS_20_21_port, REGISTERS_20_20_port, REGISTERS_20_19_port, 
      REGISTERS_20_18_port, REGISTERS_20_17_port, REGISTERS_20_16_port, 
      REGISTERS_20_15_port, REGISTERS_20_14_port, REGISTERS_20_13_port, 
      REGISTERS_20_12_port, REGISTERS_20_11_port, REGISTERS_20_10_port, 
      REGISTERS_20_9_port, REGISTERS_20_8_port, REGISTERS_20_7_port, 
      REGISTERS_20_6_port, REGISTERS_20_5_port, REGISTERS_20_4_port, 
      REGISTERS_20_3_port, REGISTERS_20_2_port, REGISTERS_20_1_port, 
      REGISTERS_20_0_port, REGISTERS_21_31_port, REGISTERS_21_30_port, 
      REGISTERS_21_29_port, REGISTERS_21_28_port, REGISTERS_21_27_port, 
      REGISTERS_21_26_port, REGISTERS_21_25_port, REGISTERS_21_24_port, 
      REGISTERS_21_23_port, REGISTERS_21_22_port, REGISTERS_21_21_port, 
      REGISTERS_21_20_port, REGISTERS_21_19_port, REGISTERS_21_18_port, 
      REGISTERS_21_17_port, REGISTERS_21_16_port, REGISTERS_21_15_port, 
      REGISTERS_21_14_port, REGISTERS_21_13_port, REGISTERS_21_12_port, 
      REGISTERS_21_11_port, REGISTERS_21_10_port, REGISTERS_21_9_port, 
      REGISTERS_21_8_port, REGISTERS_21_7_port, REGISTERS_21_6_port, 
      REGISTERS_21_5_port, REGISTERS_21_4_port, REGISTERS_21_3_port, 
      REGISTERS_21_2_port, REGISTERS_21_1_port, REGISTERS_21_0_port, 
      REGISTERS_22_31_port, REGISTERS_22_30_port, REGISTERS_22_29_port, 
      REGISTERS_22_28_port, REGISTERS_22_27_port, REGISTERS_22_26_port, 
      REGISTERS_22_25_port, REGISTERS_22_24_port, REGISTERS_22_23_port, 
      REGISTERS_22_22_port, REGISTERS_22_21_port, REGISTERS_22_20_port, 
      REGISTERS_22_19_port, REGISTERS_22_18_port, REGISTERS_22_17_port, 
      REGISTERS_22_16_port, REGISTERS_22_15_port, REGISTERS_22_14_port, 
      REGISTERS_22_13_port, REGISTERS_22_12_port, REGISTERS_22_11_port, 
      REGISTERS_22_10_port, REGISTERS_22_9_port, REGISTERS_22_8_port, 
      REGISTERS_22_7_port, REGISTERS_22_6_port, REGISTERS_22_5_port, 
      REGISTERS_22_4_port, REGISTERS_22_3_port, REGISTERS_22_2_port, 
      REGISTERS_22_1_port, REGISTERS_22_0_port, REGISTERS_23_31_port, 
      REGISTERS_23_30_port, REGISTERS_23_29_port, REGISTERS_23_28_port, 
      REGISTERS_23_27_port, REGISTERS_23_26_port, REGISTERS_23_25_port, 
      REGISTERS_23_24_port, REGISTERS_23_23_port, REGISTERS_23_22_port, 
      REGISTERS_23_21_port, REGISTERS_23_20_port, REGISTERS_23_19_port, 
      REGISTERS_23_18_port, REGISTERS_23_17_port, REGISTERS_23_16_port, 
      REGISTERS_23_15_port, REGISTERS_23_14_port, REGISTERS_23_13_port, 
      REGISTERS_23_12_port, REGISTERS_23_11_port, REGISTERS_23_10_port, 
      REGISTERS_23_9_port, REGISTERS_23_8_port, REGISTERS_23_7_port, 
      REGISTERS_23_6_port, REGISTERS_23_5_port, REGISTERS_23_4_port, 
      REGISTERS_23_3_port, REGISTERS_23_2_port, REGISTERS_23_1_port, 
      REGISTERS_23_0_port, REGISTERS_24_31_port, REGISTERS_24_30_port, 
      REGISTERS_24_29_port, REGISTERS_24_28_port, REGISTERS_24_27_port, 
      REGISTERS_24_26_port, REGISTERS_24_25_port, REGISTERS_24_24_port, 
      REGISTERS_24_23_port, REGISTERS_24_22_port, REGISTERS_24_21_port, 
      REGISTERS_24_20_port, REGISTERS_24_19_port, REGISTERS_24_18_port, 
      REGISTERS_24_17_port, REGISTERS_24_16_port, REGISTERS_24_15_port, 
      REGISTERS_24_14_port, REGISTERS_24_13_port, REGISTERS_24_12_port, 
      REGISTERS_24_11_port, REGISTERS_24_10_port, REGISTERS_24_9_port, 
      REGISTERS_24_8_port, REGISTERS_24_7_port, REGISTERS_24_6_port, 
      REGISTERS_24_5_port, REGISTERS_24_4_port, REGISTERS_24_3_port, 
      REGISTERS_24_2_port, REGISTERS_24_1_port, REGISTERS_24_0_port, 
      REGISTERS_25_31_port, REGISTERS_25_30_port, REGISTERS_25_29_port, 
      REGISTERS_25_28_port, REGISTERS_25_27_port, REGISTERS_25_26_port, 
      REGISTERS_25_25_port, REGISTERS_25_24_port, REGISTERS_25_23_port, 
      REGISTERS_25_22_port, REGISTERS_25_21_port, REGISTERS_25_20_port, 
      REGISTERS_25_19_port, REGISTERS_25_18_port, REGISTERS_25_17_port, 
      REGISTERS_25_16_port, REGISTERS_25_15_port, REGISTERS_25_14_port, 
      REGISTERS_25_13_port, REGISTERS_25_12_port, REGISTERS_25_11_port, 
      REGISTERS_25_10_port, REGISTERS_25_9_port, REGISTERS_25_8_port, 
      REGISTERS_25_7_port, REGISTERS_25_6_port, REGISTERS_25_5_port, 
      REGISTERS_25_4_port, REGISTERS_25_3_port, REGISTERS_25_2_port, 
      REGISTERS_25_1_port, REGISTERS_25_0_port, REGISTERS_26_31_port, 
      REGISTERS_26_30_port, REGISTERS_26_29_port, REGISTERS_26_28_port, 
      REGISTERS_26_27_port, REGISTERS_26_26_port, REGISTERS_26_25_port, 
      REGISTERS_26_24_port, REGISTERS_26_23_port, REGISTERS_26_22_port, 
      REGISTERS_26_21_port, REGISTERS_26_20_port, REGISTERS_26_19_port, 
      REGISTERS_26_18_port, REGISTERS_26_17_port, REGISTERS_26_16_port, 
      REGISTERS_26_15_port, REGISTERS_26_14_port, REGISTERS_26_13_port, 
      REGISTERS_26_12_port, REGISTERS_26_11_port, REGISTERS_26_10_port, 
      REGISTERS_26_9_port, REGISTERS_26_8_port, REGISTERS_26_7_port, 
      REGISTERS_26_6_port, REGISTERS_26_5_port, REGISTERS_26_4_port, 
      REGISTERS_26_3_port, REGISTERS_26_2_port, REGISTERS_26_1_port, 
      REGISTERS_26_0_port, REGISTERS_27_31_port, REGISTERS_27_30_port, 
      REGISTERS_27_29_port, REGISTERS_27_28_port, REGISTERS_27_27_port, 
      REGISTERS_27_26_port, REGISTERS_27_25_port, REGISTERS_27_24_port, 
      REGISTERS_27_23_port, REGISTERS_27_22_port, REGISTERS_27_21_port, 
      REGISTERS_27_20_port, REGISTERS_27_19_port, REGISTERS_27_18_port, 
      REGISTERS_27_17_port, REGISTERS_27_16_port, REGISTERS_27_15_port, 
      REGISTERS_27_14_port, REGISTERS_27_13_port, REGISTERS_27_12_port, 
      REGISTERS_27_11_port, REGISTERS_27_10_port, REGISTERS_27_9_port, 
      REGISTERS_27_8_port, REGISTERS_27_7_port, REGISTERS_27_6_port, 
      REGISTERS_27_5_port, REGISTERS_27_4_port, REGISTERS_27_3_port, 
      REGISTERS_27_2_port, REGISTERS_27_1_port, REGISTERS_27_0_port, 
      REGISTERS_28_31_port, REGISTERS_28_30_port, REGISTERS_28_29_port, 
      REGISTERS_28_28_port, REGISTERS_28_27_port, REGISTERS_28_26_port, 
      REGISTERS_28_25_port, REGISTERS_28_24_port, REGISTERS_28_23_port, 
      REGISTERS_28_22_port, REGISTERS_28_21_port, REGISTERS_28_20_port, 
      REGISTERS_28_19_port, REGISTERS_28_18_port, REGISTERS_28_17_port, 
      REGISTERS_28_16_port, REGISTERS_28_15_port, REGISTERS_28_14_port, 
      REGISTERS_28_13_port, REGISTERS_28_12_port, REGISTERS_28_11_port, 
      REGISTERS_28_10_port, REGISTERS_28_9_port, REGISTERS_28_8_port, 
      REGISTERS_28_7_port, REGISTERS_28_6_port, REGISTERS_28_5_port, 
      REGISTERS_28_4_port, REGISTERS_28_3_port, REGISTERS_28_2_port, 
      REGISTERS_28_1_port, REGISTERS_28_0_port, REGISTERS_29_31_port, 
      REGISTERS_29_30_port, REGISTERS_29_29_port, REGISTERS_29_28_port, 
      REGISTERS_29_27_port, REGISTERS_29_26_port, REGISTERS_29_25_port, 
      REGISTERS_29_24_port, REGISTERS_29_23_port, REGISTERS_29_22_port, 
      REGISTERS_29_21_port, REGISTERS_29_20_port, REGISTERS_29_19_port, 
      REGISTERS_29_18_port, REGISTERS_29_17_port, REGISTERS_29_16_port, 
      REGISTERS_29_15_port, REGISTERS_29_14_port, REGISTERS_29_13_port, 
      REGISTERS_29_12_port, REGISTERS_29_11_port, REGISTERS_29_10_port, 
      REGISTERS_29_9_port, REGISTERS_29_8_port, REGISTERS_29_7_port, 
      REGISTERS_29_6_port, REGISTERS_29_5_port, REGISTERS_29_4_port, 
      REGISTERS_29_3_port, REGISTERS_29_2_port, REGISTERS_29_1_port, 
      REGISTERS_29_0_port, REGISTERS_30_31_port, REGISTERS_30_30_port, 
      REGISTERS_30_29_port, REGISTERS_30_28_port, REGISTERS_30_27_port, 
      REGISTERS_30_26_port, REGISTERS_30_25_port, REGISTERS_30_24_port, 
      REGISTERS_30_23_port, REGISTERS_30_22_port, REGISTERS_30_21_port, 
      REGISTERS_30_20_port, REGISTERS_30_19_port, REGISTERS_30_18_port, 
      REGISTERS_30_17_port, REGISTERS_30_16_port, REGISTERS_30_15_port, 
      REGISTERS_30_14_port, REGISTERS_30_13_port, REGISTERS_30_12_port, 
      REGISTERS_30_11_port, REGISTERS_30_10_port, REGISTERS_30_9_port, 
      REGISTERS_30_8_port, REGISTERS_30_7_port, REGISTERS_30_6_port, 
      REGISTERS_30_5_port, REGISTERS_30_4_port, REGISTERS_30_3_port, 
      REGISTERS_30_2_port, REGISTERS_30_1_port, REGISTERS_30_0_port, 
      REGISTERS_31_31_port, REGISTERS_31_30_port, REGISTERS_31_29_port, 
      REGISTERS_31_28_port, REGISTERS_31_27_port, REGISTERS_31_26_port, 
      REGISTERS_31_25_port, REGISTERS_31_24_port, REGISTERS_31_23_port, 
      REGISTERS_31_22_port, REGISTERS_31_21_port, REGISTERS_31_20_port, 
      REGISTERS_31_19_port, REGISTERS_31_18_port, REGISTERS_31_17_port, 
      REGISTERS_31_16_port, REGISTERS_31_15_port, REGISTERS_31_14_port, 
      REGISTERS_31_13_port, REGISTERS_31_12_port, REGISTERS_31_11_port, 
      REGISTERS_31_10_port, REGISTERS_31_9_port, REGISTERS_31_8_port, 
      REGISTERS_31_7_port, REGISTERS_31_6_port, REGISTERS_31_5_port, 
      REGISTERS_31_4_port, REGISTERS_31_3_port, REGISTERS_31_2_port, 
      REGISTERS_31_1_port, REGISTERS_31_0_port, N243, N244, N245, N246, N247, 
      N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, 
      N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, n35412, 
      n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, 
      n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, 
      n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, 
      n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, 
      n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, 
      n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, 
      n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, 
      n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, 
      n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, 
      n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, 
      n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, 
      n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, 
      n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, 
      n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, 
      n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, 
      n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, 
      n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, 
      n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, 
      n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, 
      n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, 
      n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, 
      n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, 
      n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, 
      n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, 
      n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, 
      n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, 
      n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, 
      n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, 
      n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, 
      n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, 
      n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, 
      n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, 
      n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, 
      n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, 
      n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, 
      n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, 
      n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, 
      n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, 
      n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, 
      n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, 
      n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, 
      n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, 
      n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, 
      n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, 
      n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, 
      n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, 
      n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, 
      n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, 
      n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, 
      n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, 
      n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, 
      n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, 
      n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, 
      n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, 
      n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, 
      n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, 
      n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, 
      n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, 
      n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, 
      n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, 
      n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, 
      n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, 
      n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, 
      n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, 
      n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, 
      n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, 
      n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, 
      n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, 
      n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, 
      n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, 
      n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, 
      n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, 
      n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, 
      n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, 
      n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, 
      n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, 
      n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, 
      n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, 
      n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, 
      n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, 
      n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, 
      n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, 
      n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, 
      n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, 
      n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, 
      n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, 
      n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, 
      n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, 
      n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, 
      n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, 
      n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, 
      n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, 
      n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, 
      n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, 
      n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, 
      n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, 
      n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, 
      n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, 
      n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, 
      n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, 
      n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, 
      n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, 
      n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, 
      n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, 
      n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, 
      n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, 
      n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, 
      n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, 
      n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, 
      n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, 
      n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, 
      n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, 
      n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, 
      n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, 
      n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, 
      n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, 
      n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, 
      n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, 
      n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, 
      n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, 
      n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, 
      n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, 
      n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, 
      n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, 
      n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, 
      n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, 
      n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, 
      n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, 
      n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, 
      n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, 
      n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, 
      n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, 
      n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, 
      n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, 
      n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, 
      n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, 
      n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, 
      n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, 
      n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, 
      n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, 
      n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, 
      n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, 
      n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, 
      n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, 
      n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, 
      n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, 
      n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, 
      n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, 
      n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, 
      n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, 
      n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, 
      n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, 
      n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, 
      n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, 
      n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, 
      n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, 
      n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, 
      n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, 
      n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, 
      n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, 
      n36853, n36854, n36855, n36856, n36857, n36858 : std_logic;

begin
   
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => N305, D => N275, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => N305, D => N274, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => N305, D => N273, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => n36299, D => N272, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => N305, D => N271, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N305, D => N270, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => N305, D => N269, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => N305, D => N268, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => N305, D => N267, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => N305, D => N266, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => n36299, D => N265, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => n36299, D => N264, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => n36299, D => N263, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => n36299, D => N262, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => n36299, D => N261, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => N305, D => N260, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N305, D => N259, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => n36299, D => N258, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N305, D => N257, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N305, D => N256, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => n36299, D => N255, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => n36299, D => N254, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => n36299, D => N253, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => n36299, D => N252, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => n36299, D => N251, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => N305, D => N250, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => n36299, D => N249, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => n36299, D => N248, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => n36299, D => N247, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => n36299, D => N246, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => N305, D => N245, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => n36299, D => N244, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => N304, D => N275, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => N304, D => N274, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => N304, D => N273, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => N304, D => N272, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => N304, D => N271, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => N304, D => N270, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => n36300, D => N269, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => n36300, D => N268, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => n36300, D => N267, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => n36300, D => N266, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => N304, D => N265, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => N304, D => N264, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => n36300, D => N263, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => n36300, D => N262, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => n36300, D => N261, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N304, D => N260, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => N304, D => N259, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N304, D => N258, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N304, D => N257, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N304, D => N256, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => n36300, D => N255, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => n36300, D => N254, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => n36300, D => N253, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => n36300, D => N252, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => n36300, D => N251, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => N304, D => N250, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => n36300, D => N249, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => n36300, D => N248, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => n36300, D => N247, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => n36300, D => N246, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => N304, D => N245, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => n36300, D => N244, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => N303, D => N275, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => N303, D => N274, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => N303, D => N273, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => N303, D => N272, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => N303, D => N271, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => N303, D => N270, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => n36301, D => N269, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => n36301, D => N268, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => n36301, D => N267, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => n36301, D => N266, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => N303, D => N265, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => N303, D => N264, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => n36301, D => N263, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => n36301, D => N262, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => n36301, D => N261, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N303, D => N260, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => N303, D => N259, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N303, D => N258, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N303, D => N257, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N303, D => N256, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => n36301, D => N255, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => n36301, D => N254, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => n36301, D => N253, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => n36301, D => N252, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => n36301, D => N251, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => N303, D => N250, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => n36301, D => N249, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => n36301, D => N248, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => n36301, D => N247, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => n36301, D => N246, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => N303, D => N245, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => n36301, D => N244, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => N302, D => N275, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => N302, D => N274, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => N302, D => N273, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => N302, D => N272, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => N302, D => N271, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => N302, D => N270, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => n36302, D => N269, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => n36302, D => N268, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => n36302, D => N267, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => n36302, D => N266, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => N302, D => N265, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => N302, D => N264, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => n36302, D => N263, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => n36302, D => N262, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => n36302, D => N261, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N302, D => N260, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => N302, D => N259, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N302, D => N258, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N302, D => N257, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N302, D => N256, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => n36302, D => N255, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => n36302, D => N254, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => n36302, D => N253, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => n36302, D => N252, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => n36302, D => N251, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => N302, D => N250, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => n36302, D => N249, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => n36302, D => N248, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => n36302, D => N247, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => n36302, D => N246, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => N302, D => N245, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => n36302, D => N244, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => N301, D => N275, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => N301, D => N274, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => N301, D => N273, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => N301, D => N272, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => N301, D => N271, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => N301, D => N270, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => n36303, D => N269, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => n36303, D => N268, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => n36303, D => N267, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => n36303, D => N266, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => N301, D => N265, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => N301, D => N264, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => n36303, D => N263, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => n36303, D => N262, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => n36303, D => N261, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N301, D => N260, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => N301, D => N259, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N301, D => N258, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N301, D => N257, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N301, D => N256, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => n36303, D => N255, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => n36303, D => N254, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => n36303, D => N253, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => n36303, D => N252, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => n36303, D => N251, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => N301, D => N250, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => n36303, D => N249, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => n36303, D => N248, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => n36303, D => N247, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => n36303, D => N246, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => N301, D => N245, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => n36303, D => N244, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => N300, D => N275, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => N300, D => N274, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => N300, D => N273, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => N300, D => N272, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => N300, D => N271, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => N300, D => N270, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => n36304, D => N269, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => n36304, D => N268, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => n36304, D => N267, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => n36304, D => N266, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => N300, D => N265, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => N300, D => N264, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => n36304, D => N263, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => n36304, D => N262, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => n36304, D => N261, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N300, D => N260, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => N300, D => N259, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N300, D => N258, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N300, D => N257, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N300, D => N256, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => n36304, D => N255, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => n36304, D => N254, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => n36304, D => N253, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => n36304, D => N252, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => n36304, D => N251, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => N300, D => N250, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => n36304, D => N249, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => n36304, D => N248, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => n36304, D => N247, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => n36304, D => N246, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => N300, D => N245, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => n36304, D => N244, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => N299, D => N275, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => N299, D => N274, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => N299, D => N273, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => N299, D => N272, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => N299, D => N271, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => N299, D => N270, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => n36305, D => N269, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => n36305, D => N268, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => n36305, D => N267, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => n36305, D => N266, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => N299, D => N265, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => N299, D => N264, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => n36305, D => N263, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => n36305, D => N262, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => n36305, D => N261, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N299, D => N260, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => N299, D => N259, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N299, D => N258, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N299, D => N257, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N299, D => N256, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => n36305, D => N255, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => n36305, D => N254, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => n36305, D => N253, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => n36305, D => N252, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => n36305, D => N251, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => N299, D => N250, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => n36305, D => N249, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => n36305, D => N248, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => n36305, D => N247, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => n36305, D => N246, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => N299, D => N245, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => n36305, D => N244, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => N298, D => N275, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => N298, D => N274, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => N298, D => N273, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => N298, D => N272, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => N298, D => N271, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => N298, D => N270, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => n36306, D => N269, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => n36306, D => N268, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => n36306, D => N267, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => n36306, D => N266, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => N298, D => N265, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => N298, D => N264, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => n36306, D => N263, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => n36306, D => N262, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => n36306, D => N261, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => n36306, D => N260, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => N298, D => N259, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N298, D => N258, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N298, D => N257, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N298, D => N256, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => n36306, D => N255, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => n36306, D => N254, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => n36306, D => N253, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => n36306, D => N252, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => n36306, D => N251, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => N298, D => N250, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => n36306, D => N249, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => n36306, D => N248, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => n36306, D => N247, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => n36306, D => N246, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => N298, D => N245, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N298, D => N244, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => N297, D => N275, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => N297, D => N274, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => N297, D => N273, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => N297, D => N272, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => N297, D => N271, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => N297, D => N270, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => n36307, D => N269, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => n36307, D => N268, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => n36307, D => N267, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => n36307, D => N266, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => N297, D => N265, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => N297, D => N264, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => n36307, D => N263, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => n36307, D => N262, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => n36307, D => N261, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N297, D => N260, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => N297, D => N259, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N297, D => N258, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N297, D => N257, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N297, D => N256, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => n36307, D => N255, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => n36307, D => N254, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => n36307, D => N253, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => n36307, D => N252, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => n36307, D => N251, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => N297, D => N250, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => n36307, D => N249, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => n36307, D => N248, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => n36307, D => N247, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => n36307, D => N246, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => N297, D => N245, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => n36307, D => N244, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => N296, D => N275, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => N296, D => N274, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => N296, D => N273, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => N296, D => N272, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => N296, D => N271, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => N296, D => N270, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => n36308, D => N269, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => n36308, D => N268, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => n36308, D => N267, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => n36308, D => N266, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => N296, D => N265, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => N296, D => N264, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => n36308, D => N263, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => n36308, D => N262, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N296, D => N261, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => n36308, D => N260, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N296, D => N259, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => N296, D => N258, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => n36308, D => N257, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N296, D => N256, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => n36308, D => N255, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => n36308, D => N254, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => n36308, D => N253, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => n36308, D => N252, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => n36308, D => N251, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => N296, D => N250, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => n36308, D => N249, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => n36308, D => N248, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => n36308, D => N247, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => n36308, D => N246, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => N296, D => N245, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N296, D => N244, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => N295, D => N275, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => N295, D => N274, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => N295, D => N273, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => N295, D => N272, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => N295, D => N271, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => N295, D => N270, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => n36309, D => N269, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => n36309, D => N268, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => n36309, D => N267, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => n36309, D => N266, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => N295, D => N265, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => N295, D => N264, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => n36309, D => N263, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => n36309, D => N262, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => n36309, D => N261, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N295, D => N260, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => N295, D => N259, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N295, D => N258, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N295, D => N257, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N295, D => N256, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => n36309, D => N255, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => n36309, D => N254, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => n36309, D => N253, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => n36309, D => N252, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => n36309, D => N251, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => N295, D => N250, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => n36309, D => N249, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => n36309, D => N248, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => n36309, D => N247, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => n36309, D => N246, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => N295, D => N245, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => n36309, D => N244, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => N294, D => N275, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => N294, D => N274, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => N294, D => N273, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => N294, D => N272, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => N294, D => N271, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => N294, D => N270, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => n36310, D => N269, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => n36310, D => N268, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => n36310, D => N267, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => n36310, D => N266, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => N294, D => N265, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => N294, D => N264, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => n36310, D => N263, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => n36310, D => N262, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => n36310, D => N261, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N294, D => N260, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => N294, D => N259, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N294, D => N258, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N294, D => N257, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N294, D => N256, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => n36310, D => N255, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => n36310, D => N254, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => n36310, D => N253, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => n36310, D => N252, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => n36310, D => N251, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => N294, D => N250, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => n36310, D => N249, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => n36310, D => N248, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => n36310, D => N247, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => n36310, D => N246, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => N294, D => N245, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => n36310, D => N244, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => N293, D => N275, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => N293, D => N274, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => N293, D => N273, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => N293, D => N272, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => N293, D => N271, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => N293, D => N270, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => n36311, D => N269, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => n36311, D => N268, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => n36311, D => N267, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => n36311, D => N266, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => N293, D => N265, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => N293, D => N264, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => n36311, D => N263, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => n36311, D => N262, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => n36311, D => N261, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N293, D => N260, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => N293, D => N259, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N293, D => N258, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N293, D => N257, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N293, D => N256, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => n36311, D => N255, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => n36311, D => N254, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => n36311, D => N253, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => n36311, D => N252, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => n36311, D => N251, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => N293, D => N250, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => n36311, D => N249, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => n36311, D => N248, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => n36311, D => N247, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => n36311, D => N246, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => N293, D => N245, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => n36311, D => N244, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => N292, D => N275, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => N292, D => N274, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => N292, D => N273, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => N292, D => N272, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => N292, D => N271, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => N292, D => N270, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => n36312, D => N269, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => n36312, D => N268, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => n36312, D => N267, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => n36312, D => N266, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => N292, D => N265, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => N292, D => N264, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => n36312, D => N263, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => n36312, D => N262, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => n36312, D => N261, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N292, D => N260, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => N292, D => N259, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N292, D => N258, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N292, D => N257, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N292, D => N256, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => n36312, D => N255, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => n36312, D => N254, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => n36312, D => N253, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => n36312, D => N252, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => n36312, D => N251, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => N292, D => N250, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => n36312, D => N249, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => n36312, D => N248, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => n36312, D => N247, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => n36312, D => N246, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => N292, D => N245, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => n36312, D => N244, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => N291, D => N275, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => N291, D => N274, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => N291, D => N273, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => N291, D => N272, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => N291, D => N271, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => N291, D => N270, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => n36313, D => N269, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => n36313, D => N268, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => n36313, D => N267, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => n36313, D => N266, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => N291, D => N265, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => N291, D => N264, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => n36313, D => N263, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => n36313, D => N262, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => n36313, D => N261, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N291, D => N260, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => N291, D => N259, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N291, D => N258, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N291, D => N257, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N291, D => N256, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => n36313, D => N255, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => n36313, D => N254, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => n36313, D => N253, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => n36313, D => N252, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => n36313, D => N251, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => N291, D => N250, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => n36313, D => N249, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => n36313, D => N248, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => n36313, D => N247, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => n36313, D => N246, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => N291, D => N245, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => n36313, D => N244, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => N290, D => N275, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => N290, D => N274, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => N290, D => N273, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => N290, D => N272, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => N290, D => N271, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => N290, D => N270, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => n36314, D => N269, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => n36314, D => N268, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => n36314, D => N267, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => n36314, D => N266, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => N290, D => N265, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => N290, D => N264, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => n36314, D => N263, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => n36314, D => N262, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => n36314, D => N261, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N290, D => N260, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => N290, D => N259, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N290, D => N258, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N290, D => N257, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N290, D => N256, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => n36314, D => N255, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => n36314, D => N254, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => n36314, D => N253, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => n36314, D => N252, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => n36314, D => N251, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => N290, D => N250, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => n36314, D => N249, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => n36314, D => N248, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => n36314, D => N247, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => n36314, D => N246, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => N290, D => N245, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => n36314, D => N244, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => N289, D => N275, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => N289, D => N274, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => N289, D => N273, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => N289, D => N272, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => N289, D => N271, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => N289, D => N270, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => n36315, D => N269, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => n36315, D => N268, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => n36315, D => N267, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => n36315, D => N266, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => N289, D => N265, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => N289, D => N264, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => n36315, D => N263, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => n36315, D => N262, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => n36315, D => N261, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N289, D => N260, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => N289, D => N259, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N289, D => N258, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N289, D => N257, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N289, D => N256, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => n36315, D => N255, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => n36315, D => N254, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => n36315, D => N253, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => n36315, D => N252, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => n36315, D => N251, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => N289, D => N250, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => n36315, D => N249, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => n36315, D => N248, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => n36315, D => N247, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => n36315, D => N246, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => N289, D => N245, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => n36315, D => N244, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => N288, D => N275, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => N288, D => N274, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => N288, D => N273, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => N288, D => N272, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => N288, D => N271, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => N288, D => N270, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => n36316, D => N269, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => n36316, D => N268, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => n36316, D => N267, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => n36316, D => N266, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => N288, D => N265, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => N288, D => N264, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => n36316, D => N263, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => n36316, D => N262, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => n36316, D => N261, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N288, D => N260, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => N288, D => N259, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N288, D => N258, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N288, D => N257, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N288, D => N256, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => n36316, D => N255, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => n36316, D => N254, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => n36316, D => N253, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => n36316, D => N252, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => n36316, D => N251, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => N288, D => N250, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => n36316, D => N249, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => n36316, D => N248, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => n36316, D => N247, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => n36316, D => N246, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => N288, D => N245, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => n36316, D => N244, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => N287, D => N275, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => N287, D => N274, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => N287, D => N273, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => N287, D => N272, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => N287, D => N271, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => N287, D => N270, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => n36317, D => N269, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => n36317, D => N268, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => n36317, D => N267, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => n36317, D => N266, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => N287, D => N265, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => N287, D => N264, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => n36317, D => N263, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => n36317, D => N262, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => n36317, D => N261, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N287, D => N260, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => N287, D => N259, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N287, D => N258, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N287, D => N257, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N287, D => N256, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => n36317, D => N255, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => n36317, D => N254, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => n36317, D => N253, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => n36317, D => N252, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => n36317, D => N251, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => N287, D => N250, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => n36317, D => N249, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => n36317, D => N248, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => n36317, D => N247, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => n36317, D => N246, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => N287, D => N245, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => n36317, D => N244, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => N286, D => N275, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => N286, D => N274, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => N286, D => N273, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => N286, D => N272, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => N286, D => N271, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => N286, D => N270, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => n36318, D => N269, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => n36318, D => N268, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => n36318, D => N267, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => n36318, D => N266, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => N286, D => N265, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => N286, D => N264, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => n36318, D => N263, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => n36318, D => N262, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => n36318, D => N261, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N286, D => N260, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => N286, D => N259, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N286, D => N258, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N286, D => N257, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N286, D => N256, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => n36318, D => N255, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => n36318, D => N254, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => n36318, D => N253, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => n36318, D => N252, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => n36318, D => N251, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => N286, D => N250, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => n36318, D => N249, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => n36318, D => N248, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => n36318, D => N247, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => n36318, D => N246, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => N286, D => N245, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => n36318, D => N244, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => N285, D => N275, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => N285, D => N274, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => N285, D => N273, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => N285, D => N272, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => N285, D => N271, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => N285, D => N270, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => n36319, D => N269, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => n36319, D => N268, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => n36319, D => N267, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => n36319, D => N266, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => N285, D => N265, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => N285, D => N264, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => n36319, D => N263, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => n36319, D => N262, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => n36319, D => N261, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N285, D => N260, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => N285, D => N259, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N285, D => N258, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N285, D => N257, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N285, D => N256, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => n36319, D => N255, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => n36319, D => N254, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => n36319, D => N253, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => n36319, D => N252, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => n36319, D => N251, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => N285, D => N250, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => n36319, D => N249, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => n36319, D => N248, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => n36319, D => N247, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => n36319, D => N246, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => N285, D => N245, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => n36319, D => N244, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => N284, D => N275, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => N284, D => N274, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => N284, D => N273, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => N284, D => N272, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => N284, D => N271, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => N284, D => N270, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => n36320, D => N269, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => n36320, D => N268, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => n36320, D => N267, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => n36320, D => N266, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => N284, D => N265, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => N284, D => N264, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => n36320, D => N263, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => n36320, D => N262, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => n36320, D => N261, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N284, D => N260, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => N284, D => N259, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N284, D => N258, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N284, D => N257, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N284, D => N256, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => n36320, D => N255, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => n36320, D => N254, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => n36320, D => N253, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => n36320, D => N252, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => n36320, D => N251, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => N284, D => N250, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => n36320, D => N249, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => n36320, D => N248, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => n36320, D => N247, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => n36320, D => N246, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => N284, D => N245, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => n36320, D => N244, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => N283, D => N275, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => N283, D => N274, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => N283, D => N273, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => N283, D => N272, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => N283, D => N271, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => N283, D => N270, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => n36321, D => N269, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => n36321, D => N268, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => n36321, D => N267, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => n36321, D => N266, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => N283, D => N265, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => N283, D => N264, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => n36321, D => N263, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => n36321, D => N262, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => n36321, D => N261, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N283, D => N260, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => N283, D => N259, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N283, D => N258, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N283, D => N257, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N283, D => N256, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => n36321, D => N255, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => n36321, D => N254, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => n36321, D => N253, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => n36321, D => N252, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => n36321, D => N251, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => N283, D => N250, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => n36321, D => N249, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => n36321, D => N248, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => n36321, D => N247, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => n36321, D => N246, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => N283, D => N245, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => n36321, D => N244, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => N282, D => N275, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => N282, D => N274, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => N282, D => N273, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => N282, D => N272, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => N282, D => N271, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => N282, D => N270, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => N282, D => N269, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => n36322, D => N268, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => n36322, D => N267, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => n36322, D => N266, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => n36322, D => N265, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => n36322, D => N264, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => N282, D => N263, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => n36322, D => N262, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N282, D => N261, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N282, D => N260, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => n36322, D => N259, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N282, D => N258, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N282, D => N257, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => n36322, D => N256, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => N282, D => N255, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => N282, D => N254, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => n36322, D => N253, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => n36322, D => N252, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => N282, D => N251, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => n36322, D => N250, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => n36322, D => N249, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => n36322, D => N248, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => n36322, D => N247, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => n36322, D => N246, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => n36322, D => N245, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => n36322, D => N244, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => N281, D => N275, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => N281, D => N274, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => N281, D => N273, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => N281, D => N272, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => N281, D => N271, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => N281, D => N270, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => n36323, D => N269, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => n36323, D => N268, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => n36323, D => N267, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => n36323, D => N266, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => N281, D => N265, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => N281, D => N264, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => n36323, D => N263, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => n36323, D => N262, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => n36323, D => N261, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N281, D => N260, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => N281, D => N259, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N281, D => N258, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N281, D => N257, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N281, D => N256, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => n36323, D => N255, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => n36323, D => N254, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => n36323, D => N253, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => n36323, D => N252, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => n36323, D => N251, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => N281, D => N250, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => n36323, D => N249, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => n36323, D => N248, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => n36323, D => N247, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => n36323, D => N246, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => N281, D => N245, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => n36323, D => N244, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => N280, D => N275, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => N280, D => N274, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => N280, D => N273, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => N280, D => N272, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => N280, D => N271, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => N280, D => N270, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => n36324, D => N269, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => n36324, D => N268, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => n36324, D => N267, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => n36324, D => N266, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => N280, D => N265, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => N280, D => N264, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => n36324, D => N263, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => n36324, D => N262, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => n36324, D => N261, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N280, D => N260, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => N280, D => N259, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N280, D => N258, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N280, D => N257, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N280, D => N256, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => n36324, D => N255, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => n36324, D => N254, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => n36324, D => N253, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => n36324, D => N252, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => n36324, D => N251, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => N280, D => N250, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => n36324, D => N249, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => n36324, D => N248, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => n36324, D => N247, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => n36324, D => N246, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => N280, D => N245, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => n36324, D => N244, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => N279, D => N275, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => N279, D => N274, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => N279, D => N273, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => N279, D => N272, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => N279, D => N271, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => N279, D => N270, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => n36325, D => N269, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => n36325, D => N268, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => n36325, D => N267, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => n36325, D => N266, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => N279, D => N265, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => N279, D => N264, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => n36325, D => N263, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => n36325, D => N262, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => n36325, D => N261, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N279, D => N260, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => N279, D => N259, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N279, D => N258, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N279, D => N257, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N279, D => N256, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => n36325, D => N255, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => n36325, D => N254, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => n36325, D => N253, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => n36325, D => N252, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => n36325, D => N251, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => N279, D => N250, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => n36325, D => N249, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => n36325, D => N248, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => n36325, D => N247, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => n36325, D => N246, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => N279, D => N245, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => n36325, D => N244, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => N278, D => N275, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => N278, D => N274, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => N278, D => N273, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => N278, D => N272, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => N278, D => N271, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => N278, D => N270, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => n36326, D => N269, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => n36326, D => N268, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => n36326, D => N267, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => n36326, D => N266, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => N278, D => N265, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => N278, D => N264, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => n36326, D => N263, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => n36326, D => N262, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => n36326, D => N261, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N278, D => N260, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => N278, D => N259, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N278, D => N258, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N278, D => N257, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N278, D => N256, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => n36326, D => N255, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => n36326, D => N254, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => n36326, D => N253, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => n36326, D => N252, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => n36326, D => N251, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => N278, D => N250, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => n36326, D => N249, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => n36326, D => N248, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => n36326, D => N247, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => n36326, D => N246, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => N278, D => N245, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => n36326, D => N244, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => N277, D => N275, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => N277, D => N274, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => N277, D => N273, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => N277, D => N272, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => N277, D => N271, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => N277, D => N270, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => n36327, D => N269, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => n36327, D => N268, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => n36327, D => N267, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => n36327, D => N266, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => N277, D => N265, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => N277, D => N264, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => n36327, D => N263, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => n36327, D => N262, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => n36327, D => N261, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N277, D => N260, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => N277, D => N259, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N277, D => N258, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N277, D => N257, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N277, D => N256, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => n36327, D => N255, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => n36327, D => N254, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => n36327, D => N253, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => n36327, D => N252, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => n36327, D => N251, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => N277, D => N250, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => n36327, D => N249, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => n36327, D => N248, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => n36327, D => N247, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => n36327, D => N246, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => N277, D => N245, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => n36327, D => N244, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => N276, D => N275, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => N276, D => N274, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => N276, D => N273, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => N276, D => N272, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => N276, D => N271, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => N276, D => N270, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => n36328, D => N269, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => n36328, D => N268, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => n36328, D => N267, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => n36328, D => N266, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => N276, D => N265, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => N276, D => N264, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => n36328, D => N263, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => n36328, D => N262, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => n36328, D => N261, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N276, D => N260, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => N276, D => N259, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N276, D => N258, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N276, D => N257, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N276, D => N256, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => n36328, D => N255, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => n36328, D => N254, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => n36328, D => N253, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => n36328, D => N252, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => n36328, D => N251, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => N276, D => N250, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => n36328, D => N249, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => n36328, D => N248, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => n36328, D => N247, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => n36328, D => N246, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => N276, D => N245, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => n36328, D => N244, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => N243, D => N275, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => N243, D => N274, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => N243, D => N273, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => N243, D => N272, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => N243, D => N271, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => N243, D => N270, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => N243, D => N269, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => N243, D => N268, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => N243, D => N267, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => N243, D => N266, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => n36329, D => N265, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => n36329, D => N264, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => n36329, D => N263, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => n36329, D => N262, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => n36329, D => N261, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N243, D => N260, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => N243, D => N259, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N243, D => N258, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N243, D => N257, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N243, D => N256, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => n36329, D => N255, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => n36329, D => N254, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => n36329, D => N253, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => n36329, D => N252, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => n36329, D => N251, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => n36329, D => N250, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => n36329, D => N249, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => n36329, D => N248, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => n36329, D => N247, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => n36329, D => N246, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => n36329, D => N245, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => n36329, D => N244, Q => 
                           REGISTERS_31_0_port);
   U3 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n36283, B1 => 
                           REGISTERS_10_16_port, B2 => n36284, ZN => n35412);
   U4 : AOI22_X1 port map( A1 => REGISTERS_18_16_port, A2 => n36285, B1 => 
                           REGISTERS_2_16_port, B2 => n36286, ZN => n35413);
   U5 : AOI22_X1 port map( A1 => REGISTERS_31_16_port, A2 => n36287, B1 => 
                           REGISTERS_3_16_port, B2 => n36288, ZN => n35414);
   U6 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n36289, B1 => 
                           REGISTERS_30_16_port, B2 => n36290, ZN => n35415);
   U7 : NAND4_X1 port map( A1 => n35412, A2 => n35413, A3 => n35414, A4 => 
                           n35415, ZN => n35416);
   U8 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n36291, B1 => 
                           REGISTERS_11_16_port, B2 => n36292, ZN => n35417);
   U9 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n36293, B1 => 
                           REGISTERS_1_16_port, B2 => n36294, ZN => n35418);
   U10 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n36295, B1 => 
                           REGISTERS_12_16_port, B2 => n36296, ZN => n35419);
   U11 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n36297, B1 => 
                           REGISTERS_20_16_port, B2 => n36298, ZN => n35420);
   U12 : NAND4_X1 port map( A1 => n35417, A2 => n35418, A3 => n35419, A4 => 
                           n35420, ZN => n35421);
   U13 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n36268, B1 => 
                           REGISTERS_5_16_port, B2 => n36269, ZN => n35422);
   U14 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n36270, B1 => 
                           REGISTERS_25_16_port, B2 => n36271, ZN => n35423);
   U15 : AOI222_X1 port map( A1 => REGISTERS_23_16_port, A2 => n36272, B1 => 
                           REGISTERS_17_16_port, B2 => n36273, C1 => 
                           REGISTERS_19_16_port, C2 => n36274, ZN => n35424);
   U16 : NAND3_X1 port map( A1 => n35422, A2 => n35423, A3 => n35424, ZN => 
                           n35425);
   U17 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n36275, B1 => 
                           REGISTERS_14_16_port, B2 => n36276, ZN => n35426);
   U18 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n36279, B1 => 
                           REGISTERS_6_16_port, B2 => n36280, ZN => n35427);
   U19 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n36281, B1 => 
                           REGISTERS_26_16_port, B2 => n36282, ZN => n35428);
   U20 : NAND4_X1 port map( A1 => n35426, A2 => n36488, A3 => n35427, A4 => 
                           n35428, ZN => n35429);
   U21 : OR4_X1 port map( A1 => n35416, A2 => n35421, A3 => n35425, A4 => 
                           n35429, ZN => OUTA(16));
   U22 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n36283, B1 => 
                           REGISTERS_10_17_port, B2 => n36284, ZN => n35430);
   U23 : AOI22_X1 port map( A1 => REGISTERS_18_17_port, A2 => n36285, B1 => 
                           REGISTERS_2_17_port, B2 => n36286, ZN => n35431);
   U24 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n36287, B1 => 
                           REGISTERS_3_17_port, B2 => n36288, ZN => n35432);
   U25 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n36289, B1 => 
                           REGISTERS_30_17_port, B2 => n36290, ZN => n35433);
   U26 : NAND4_X1 port map( A1 => n35430, A2 => n35431, A3 => n35432, A4 => 
                           n35433, ZN => n35434);
   U27 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n36291, B1 => 
                           REGISTERS_11_17_port, B2 => n36292, ZN => n35435);
   U28 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n36293, B1 => 
                           REGISTERS_1_17_port, B2 => n36294, ZN => n35436);
   U29 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n36295, B1 => 
                           REGISTERS_12_17_port, B2 => n36296, ZN => n35437);
   U30 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n36297, B1 => 
                           REGISTERS_20_17_port, B2 => n36298, ZN => n35438);
   U31 : NAND4_X1 port map( A1 => n35435, A2 => n35436, A3 => n35437, A4 => 
                           n35438, ZN => n35439);
   U32 : AOI22_X1 port map( A1 => REGISTERS_22_17_port, A2 => n36268, B1 => 
                           REGISTERS_5_17_port, B2 => n36269, ZN => n35440);
   U33 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n36270, B1 => 
                           REGISTERS_25_17_port, B2 => n36271, ZN => n35441);
   U34 : AOI222_X1 port map( A1 => REGISTERS_23_17_port, A2 => n36272, B1 => 
                           REGISTERS_17_17_port, B2 => n36273, C1 => 
                           REGISTERS_19_17_port, C2 => n36274, ZN => n35442);
   U35 : NAND3_X1 port map( A1 => n35440, A2 => n35441, A3 => n35442, ZN => 
                           n35443);
   U36 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n36275, B1 => 
                           REGISTERS_14_17_port, B2 => n36276, ZN => n35444);
   U37 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n36279, B1 => 
                           REGISTERS_6_17_port, B2 => n36280, ZN => n35445);
   U38 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n36281, B1 => 
                           REGISTERS_26_17_port, B2 => n36282, ZN => n35446);
   U39 : NAND4_X1 port map( A1 => n35444, A2 => n36489, A3 => n35445, A4 => 
                           n35446, ZN => n35447);
   U40 : OR4_X1 port map( A1 => n35434, A2 => n35439, A3 => n35443, A4 => 
                           n35447, ZN => OUTA(17));
   U41 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n36283, B1 => 
                           REGISTERS_10_18_port, B2 => n36284, ZN => n35448);
   U42 : AOI22_X1 port map( A1 => REGISTERS_18_18_port, A2 => n36285, B1 => 
                           REGISTERS_2_18_port, B2 => n36286, ZN => n35449);
   U43 : AOI22_X1 port map( A1 => REGISTERS_31_18_port, A2 => n36287, B1 => 
                           REGISTERS_3_18_port, B2 => n36288, ZN => n35450);
   U44 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n36289, B1 => 
                           REGISTERS_30_18_port, B2 => n36290, ZN => n35451);
   U45 : NAND4_X1 port map( A1 => n35448, A2 => n35449, A3 => n35450, A4 => 
                           n35451, ZN => n35452);
   U46 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n36291, B1 => 
                           REGISTERS_11_18_port, B2 => n36292, ZN => n35453);
   U47 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n36293, B1 => 
                           REGISTERS_1_18_port, B2 => n36294, ZN => n35454);
   U48 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n36295, B1 => 
                           REGISTERS_12_18_port, B2 => n36296, ZN => n35455);
   U49 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n36297, B1 => 
                           REGISTERS_20_18_port, B2 => n36298, ZN => n35456);
   U50 : NAND4_X1 port map( A1 => n35453, A2 => n35454, A3 => n35455, A4 => 
                           n35456, ZN => n35457);
   U51 : AOI22_X1 port map( A1 => REGISTERS_22_18_port, A2 => n36268, B1 => 
                           REGISTERS_5_18_port, B2 => n36269, ZN => n35458);
   U52 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n36270, B1 => 
                           REGISTERS_25_18_port, B2 => n36271, ZN => n35459);
   U53 : AOI222_X1 port map( A1 => REGISTERS_23_18_port, A2 => n36272, B1 => 
                           REGISTERS_17_18_port, B2 => n36273, C1 => 
                           REGISTERS_19_18_port, C2 => n36274, ZN => n35460);
   U54 : NAND3_X1 port map( A1 => n35458, A2 => n35459, A3 => n35460, ZN => 
                           n35461);
   U55 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n36275, B1 => 
                           REGISTERS_14_18_port, B2 => n36276, ZN => n35462);
   U56 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n36279, B1 => 
                           REGISTERS_6_18_port, B2 => n36280, ZN => n35463);
   U57 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n36281, B1 => 
                           REGISTERS_26_18_port, B2 => n36282, ZN => n35464);
   U58 : NAND4_X1 port map( A1 => n35462, A2 => n36490, A3 => n35463, A4 => 
                           n35464, ZN => n35465);
   U59 : OR4_X1 port map( A1 => n35452, A2 => n35457, A3 => n35461, A4 => 
                           n35465, ZN => OUTA(18));
   U60 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n36283, B1 => 
                           REGISTERS_10_19_port, B2 => n36284, ZN => n35466);
   U61 : AOI22_X1 port map( A1 => REGISTERS_18_19_port, A2 => n36285, B1 => 
                           REGISTERS_2_19_port, B2 => n36286, ZN => n35467);
   U62 : AOI22_X1 port map( A1 => REGISTERS_31_19_port, A2 => n36287, B1 => 
                           REGISTERS_3_19_port, B2 => n36288, ZN => n35468);
   U63 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n36289, B1 => 
                           REGISTERS_30_19_port, B2 => n36290, ZN => n35469);
   U64 : NAND4_X1 port map( A1 => n35466, A2 => n35467, A3 => n35468, A4 => 
                           n35469, ZN => n35470);
   U65 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n36291, B1 => 
                           REGISTERS_11_19_port, B2 => n36292, ZN => n35471);
   U66 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n36293, B1 => 
                           REGISTERS_1_19_port, B2 => n36294, ZN => n35472);
   U67 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n36295, B1 => 
                           REGISTERS_12_19_port, B2 => n36296, ZN => n35473);
   U68 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n36297, B1 => 
                           REGISTERS_20_19_port, B2 => n36298, ZN => n35474);
   U69 : NAND4_X1 port map( A1 => n35471, A2 => n35472, A3 => n35473, A4 => 
                           n35474, ZN => n35475);
   U70 : AOI22_X1 port map( A1 => REGISTERS_22_19_port, A2 => n36268, B1 => 
                           REGISTERS_5_19_port, B2 => n36269, ZN => n35476);
   U71 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n36270, B1 => 
                           REGISTERS_25_19_port, B2 => n36271, ZN => n35477);
   U72 : AOI222_X1 port map( A1 => REGISTERS_23_19_port, A2 => n36272, B1 => 
                           REGISTERS_17_19_port, B2 => n36273, C1 => 
                           REGISTERS_19_19_port, C2 => n36274, ZN => n35478);
   U73 : NAND3_X1 port map( A1 => n35476, A2 => n35477, A3 => n35478, ZN => 
                           n35479);
   U74 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n36275, B1 => 
                           REGISTERS_14_19_port, B2 => n36276, ZN => n35480);
   U75 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n36279, B1 => 
                           REGISTERS_6_19_port, B2 => n36280, ZN => n35481);
   U76 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n36281, B1 => 
                           REGISTERS_26_19_port, B2 => n36282, ZN => n35482);
   U77 : NAND4_X1 port map( A1 => n35480, A2 => n36491, A3 => n35481, A4 => 
                           n35482, ZN => n35483);
   U78 : OR4_X1 port map( A1 => n35470, A2 => n35475, A3 => n35479, A4 => 
                           n35483, ZN => OUTA(19));
   U79 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n36283, B1 => 
                           REGISTERS_10_20_port, B2 => n36284, ZN => n35484);
   U80 : AOI22_X1 port map( A1 => REGISTERS_18_20_port, A2 => n36285, B1 => 
                           REGISTERS_2_20_port, B2 => n36784, ZN => n35485);
   U81 : AOI22_X1 port map( A1 => REGISTERS_31_20_port, A2 => n36287, B1 => 
                           REGISTERS_3_20_port, B2 => n36288, ZN => n35486);
   U82 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n36289, B1 => 
                           REGISTERS_30_20_port, B2 => n36290, ZN => n35487);
   U83 : NAND4_X1 port map( A1 => n35484, A2 => n35485, A3 => n35486, A4 => 
                           n35487, ZN => n35488);
   U84 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n36291, B1 => 
                           REGISTERS_11_20_port, B2 => n36292, ZN => n35489);
   U85 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n36293, B1 => 
                           REGISTERS_1_20_port, B2 => n36294, ZN => n35490);
   U86 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n36295, B1 => 
                           REGISTERS_12_20_port, B2 => n36296, ZN => n35491);
   U87 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n36297, B1 => 
                           REGISTERS_20_20_port, B2 => n36298, ZN => n35492);
   U88 : NAND4_X1 port map( A1 => n35489, A2 => n35490, A3 => n35491, A4 => 
                           n35492, ZN => n35493);
   U89 : AOI22_X1 port map( A1 => REGISTERS_22_20_port, A2 => n36268, B1 => 
                           REGISTERS_5_20_port, B2 => n36269, ZN => n35494);
   U90 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n36270, B1 => 
                           REGISTERS_25_20_port, B2 => n36271, ZN => n35495);
   U91 : AOI222_X1 port map( A1 => REGISTERS_23_20_port, A2 => n36272, B1 => 
                           REGISTERS_17_20_port, B2 => n36273, C1 => 
                           REGISTERS_19_20_port, C2 => n36274, ZN => n35496);
   U92 : NAND3_X1 port map( A1 => n35494, A2 => n35495, A3 => n35496, ZN => 
                           n35497);
   U93 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n36275, B1 => 
                           REGISTERS_14_20_port, B2 => n36276, ZN => n35498);
   U94 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n36279, B1 => 
                           REGISTERS_6_20_port, B2 => n36280, ZN => n35499);
   U95 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n36281, B1 => 
                           REGISTERS_26_20_port, B2 => n36282, ZN => n35500);
   U96 : NAND4_X1 port map( A1 => n35498, A2 => n36512, A3 => n35499, A4 => 
                           n35500, ZN => n35501);
   U97 : OR4_X1 port map( A1 => n35488, A2 => n35493, A3 => n35497, A4 => 
                           n35501, ZN => OUTA(20));
   U98 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n36283, B1 => 
                           REGISTERS_10_21_port, B2 => n36284, ZN => n35502);
   U99 : AOI22_X1 port map( A1 => REGISTERS_18_21_port, A2 => n36285, B1 => 
                           REGISTERS_2_21_port, B2 => n36286, ZN => n35503);
   U100 : AOI22_X1 port map( A1 => REGISTERS_31_21_port, A2 => n36287, B1 => 
                           REGISTERS_3_21_port, B2 => n36288, ZN => n35504);
   U101 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n36289, B1 => 
                           REGISTERS_30_21_port, B2 => n36290, ZN => n35505);
   U102 : NAND4_X1 port map( A1 => n35502, A2 => n35503, A3 => n35504, A4 => 
                           n35505, ZN => n35506);
   U103 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n36291, B1 => 
                           REGISTERS_11_21_port, B2 => n36292, ZN => n35507);
   U104 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n36293, B1 => 
                           REGISTERS_1_21_port, B2 => n36294, ZN => n35508);
   U105 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n36295, B1 => 
                           REGISTERS_12_21_port, B2 => n36296, ZN => n35509);
   U106 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n36297, B1 => 
                           REGISTERS_20_21_port, B2 => n36298, ZN => n35510);
   U107 : NAND4_X1 port map( A1 => n35507, A2 => n35508, A3 => n35509, A4 => 
                           n35510, ZN => n35511);
   U108 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n36268, B1 => 
                           REGISTERS_5_21_port, B2 => n36269, ZN => n35512);
   U109 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n36270, B1 => 
                           REGISTERS_25_21_port, B2 => n36271, ZN => n35513);
   U110 : AOI222_X1 port map( A1 => REGISTERS_23_21_port, A2 => n36272, B1 => 
                           REGISTERS_17_21_port, B2 => n36273, C1 => 
                           REGISTERS_19_21_port, C2 => n36274, ZN => n35514);
   U111 : NAND3_X1 port map( A1 => n35512, A2 => n35513, A3 => n35514, ZN => 
                           n35515);
   U112 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n36275, B1 => 
                           REGISTERS_14_21_port, B2 => n36276, ZN => n35516);
   U113 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n36279, B1 => 
                           REGISTERS_6_21_port, B2 => n36280, ZN => n35517);
   U114 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n36281, B1 => 
                           REGISTERS_26_21_port, B2 => n36282, ZN => n35518);
   U115 : NAND4_X1 port map( A1 => n35516, A2 => n36513, A3 => n35517, A4 => 
                           n35518, ZN => n35519);
   U116 : OR4_X1 port map( A1 => n35506, A2 => n35511, A3 => n35515, A4 => 
                           n35519, ZN => OUTA(21));
   U117 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n36283, B1 => 
                           REGISTERS_10_22_port, B2 => n36284, ZN => n35520);
   U118 : AOI22_X1 port map( A1 => REGISTERS_18_22_port, A2 => n36285, B1 => 
                           REGISTERS_2_22_port, B2 => n36286, ZN => n35521);
   U119 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n36287, B1 => 
                           REGISTERS_3_22_port, B2 => n36288, ZN => n35522);
   U120 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n36289, B1 => 
                           REGISTERS_30_22_port, B2 => n36290, ZN => n35523);
   U121 : NAND4_X1 port map( A1 => n35520, A2 => n35521, A3 => n35522, A4 => 
                           n35523, ZN => n35524);
   U122 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n36291, B1 => 
                           REGISTERS_11_22_port, B2 => n36292, ZN => n35525);
   U123 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n36293, B1 => 
                           REGISTERS_1_22_port, B2 => n36294, ZN => n35526);
   U124 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n36295, B1 => 
                           REGISTERS_12_22_port, B2 => n36296, ZN => n35527);
   U125 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n36297, B1 => 
                           REGISTERS_20_22_port, B2 => n36298, ZN => n35528);
   U126 : NAND4_X1 port map( A1 => n35525, A2 => n35526, A3 => n35527, A4 => 
                           n35528, ZN => n35529);
   U127 : AOI22_X1 port map( A1 => REGISTERS_22_22_port, A2 => n36268, B1 => 
                           REGISTERS_5_22_port, B2 => n36269, ZN => n35530);
   U128 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n36270, B1 => 
                           REGISTERS_25_22_port, B2 => n36271, ZN => n35531);
   U129 : AOI222_X1 port map( A1 => REGISTERS_23_22_port, A2 => n36272, B1 => 
                           REGISTERS_17_22_port, B2 => n36273, C1 => 
                           REGISTERS_19_22_port, C2 => n36274, ZN => n35532);
   U130 : NAND3_X1 port map( A1 => n35530, A2 => n35531, A3 => n35532, ZN => 
                           n35533);
   U131 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n36275, B1 => 
                           REGISTERS_14_22_port, B2 => n36276, ZN => n35534);
   U132 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n36279, B1 => 
                           REGISTERS_6_22_port, B2 => n36280, ZN => n35535);
   U133 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n36281, B1 => 
                           REGISTERS_26_22_port, B2 => n36282, ZN => n35536);
   U134 : NAND4_X1 port map( A1 => n35534, A2 => n36514, A3 => n35535, A4 => 
                           n35536, ZN => n35537);
   U135 : OR4_X1 port map( A1 => n35524, A2 => n35529, A3 => n35533, A4 => 
                           n35537, ZN => OUTA(22));
   U136 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n36283, B1 => 
                           REGISTERS_10_23_port, B2 => n36284, ZN => n35538);
   U137 : AOI22_X1 port map( A1 => REGISTERS_18_23_port, A2 => n36285, B1 => 
                           REGISTERS_2_23_port, B2 => n36286, ZN => n35539);
   U138 : AOI22_X1 port map( A1 => REGISTERS_31_23_port, A2 => n36287, B1 => 
                           REGISTERS_3_23_port, B2 => n36288, ZN => n35540);
   U139 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n36289, B1 => 
                           REGISTERS_30_23_port, B2 => n36290, ZN => n35541);
   U140 : NAND4_X1 port map( A1 => n35538, A2 => n35539, A3 => n35540, A4 => 
                           n35541, ZN => n35542);
   U141 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n36291, B1 => 
                           REGISTERS_11_23_port, B2 => n36292, ZN => n35543);
   U142 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n36293, B1 => 
                           REGISTERS_1_23_port, B2 => n36294, ZN => n35544);
   U143 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n36295, B1 => 
                           REGISTERS_12_23_port, B2 => n36296, ZN => n35545);
   U144 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n36297, B1 => 
                           REGISTERS_20_23_port, B2 => n36298, ZN => n35546);
   U145 : NAND4_X1 port map( A1 => n35543, A2 => n35544, A3 => n35545, A4 => 
                           n35546, ZN => n35547);
   U146 : AOI22_X1 port map( A1 => REGISTERS_22_23_port, A2 => n36268, B1 => 
                           REGISTERS_5_23_port, B2 => n36269, ZN => n35548);
   U147 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n36270, B1 => 
                           REGISTERS_25_23_port, B2 => n36271, ZN => n35549);
   U148 : AOI222_X1 port map( A1 => REGISTERS_23_23_port, A2 => n36272, B1 => 
                           REGISTERS_17_23_port, B2 => n36273, C1 => 
                           REGISTERS_19_23_port, C2 => n36274, ZN => n35550);
   U149 : NAND3_X1 port map( A1 => n35548, A2 => n35549, A3 => n35550, ZN => 
                           n35551);
   U150 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n36275, B1 => 
                           REGISTERS_14_23_port, B2 => n36276, ZN => n35552);
   U151 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n36279, B1 => 
                           REGISTERS_6_23_port, B2 => n36280, ZN => n35553);
   U152 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n36281, B1 => 
                           REGISTERS_26_23_port, B2 => n36282, ZN => n35554);
   U153 : NAND4_X1 port map( A1 => n35552, A2 => n36515, A3 => n35553, A4 => 
                           n35554, ZN => n35555);
   U154 : OR4_X1 port map( A1 => n35542, A2 => n35547, A3 => n35551, A4 => 
                           n35555, ZN => OUTA(23));
   U155 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n36283, B1 => 
                           REGISTERS_10_24_port, B2 => n36284, ZN => n35556);
   U156 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n36285, B1 => 
                           REGISTERS_2_24_port, B2 => n36286, ZN => n35557);
   U157 : AOI22_X1 port map( A1 => REGISTERS_31_24_port, A2 => n36287, B1 => 
                           REGISTERS_3_24_port, B2 => n36288, ZN => n35558);
   U158 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n36289, B1 => 
                           REGISTERS_30_24_port, B2 => n36290, ZN => n35559);
   U159 : NAND4_X1 port map( A1 => n35556, A2 => n35557, A3 => n35558, A4 => 
                           n35559, ZN => n35560);
   U160 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n36291, B1 => 
                           REGISTERS_11_24_port, B2 => n36292, ZN => n35561);
   U161 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n36293, B1 => 
                           REGISTERS_1_24_port, B2 => n36294, ZN => n35562);
   U162 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n36295, B1 => 
                           REGISTERS_12_24_port, B2 => n36296, ZN => n35563);
   U163 : AOI22_X1 port map( A1 => REGISTERS_15_24_port, A2 => n36297, B1 => 
                           REGISTERS_20_24_port, B2 => n36298, ZN => n35564);
   U164 : NAND4_X1 port map( A1 => n35561, A2 => n35562, A3 => n35563, A4 => 
                           n35564, ZN => n35565);
   U165 : AOI22_X1 port map( A1 => REGISTERS_22_24_port, A2 => n36268, B1 => 
                           REGISTERS_5_24_port, B2 => n36269, ZN => n35566);
   U166 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n36270, B1 => 
                           REGISTERS_25_24_port, B2 => n36271, ZN => n35567);
   U167 : AOI222_X1 port map( A1 => REGISTERS_23_24_port, A2 => n36272, B1 => 
                           REGISTERS_17_24_port, B2 => n36273, C1 => 
                           REGISTERS_19_24_port, C2 => n36274, ZN => n35568);
   U168 : NAND3_X1 port map( A1 => n35566, A2 => n35567, A3 => n35568, ZN => 
                           n35569);
   U169 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n36275, B1 => 
                           REGISTERS_14_24_port, B2 => n36276, ZN => n35570);
   U170 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n36279, B1 => 
                           REGISTERS_6_24_port, B2 => n36280, ZN => n35571);
   U171 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n36281, B1 => 
                           REGISTERS_26_24_port, B2 => n36282, ZN => n35572);
   U172 : NAND4_X1 port map( A1 => n35570, A2 => n36516, A3 => n35571, A4 => 
                           n35572, ZN => n35573);
   U173 : OR4_X1 port map( A1 => n35560, A2 => n35565, A3 => n35569, A4 => 
                           n35573, ZN => OUTA(24));
   U174 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n36283, B1 => 
                           REGISTERS_10_25_port, B2 => n36284, ZN => n35574);
   U175 : AOI22_X1 port map( A1 => REGISTERS_18_25_port, A2 => n36285, B1 => 
                           REGISTERS_2_25_port, B2 => n36286, ZN => n35575);
   U176 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n36287, B1 => 
                           REGISTERS_3_25_port, B2 => n36288, ZN => n35576);
   U177 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n36289, B1 => 
                           REGISTERS_30_25_port, B2 => n36290, ZN => n35577);
   U178 : NAND4_X1 port map( A1 => n35574, A2 => n35575, A3 => n35576, A4 => 
                           n35577, ZN => n35578);
   U179 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n36291, B1 => 
                           REGISTERS_11_25_port, B2 => n36292, ZN => n35579);
   U180 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n36293, B1 => 
                           REGISTERS_1_25_port, B2 => n36294, ZN => n35580);
   U181 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n36295, B1 => 
                           REGISTERS_12_25_port, B2 => n36296, ZN => n35581);
   U182 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n36297, B1 => 
                           REGISTERS_20_25_port, B2 => n36298, ZN => n35582);
   U183 : NAND4_X1 port map( A1 => n35579, A2 => n35580, A3 => n35581, A4 => 
                           n35582, ZN => n35583);
   U184 : AOI22_X1 port map( A1 => REGISTERS_22_25_port, A2 => n36268, B1 => 
                           REGISTERS_5_25_port, B2 => n36269, ZN => n35584);
   U185 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n36270, B1 => 
                           REGISTERS_25_25_port, B2 => n36271, ZN => n35585);
   U186 : AOI222_X1 port map( A1 => REGISTERS_23_25_port, A2 => n36272, B1 => 
                           REGISTERS_17_25_port, B2 => n36273, C1 => 
                           REGISTERS_19_25_port, C2 => n36274, ZN => n35586);
   U187 : NAND3_X1 port map( A1 => n35584, A2 => n35585, A3 => n35586, ZN => 
                           n35587);
   U188 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n36275, B1 => 
                           REGISTERS_14_25_port, B2 => n36276, ZN => n35588);
   U189 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n36279, B1 => 
                           REGISTERS_6_25_port, B2 => n36280, ZN => n35589);
   U190 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n36281, B1 => 
                           REGISTERS_26_25_port, B2 => n36282, ZN => n35590);
   U191 : NAND4_X1 port map( A1 => n35588, A2 => n36517, A3 => n35589, A4 => 
                           n35590, ZN => n35591);
   U192 : OR4_X1 port map( A1 => n35578, A2 => n35583, A3 => n35587, A4 => 
                           n35591, ZN => OUTA(25));
   U193 : AOI22_X1 port map( A1 => n36283, A2 => REGISTERS_9_0_port, B1 => 
                           n36284, B2 => REGISTERS_10_0_port, ZN => n35592);
   U194 : AOI22_X1 port map( A1 => n36285, A2 => REGISTERS_18_0_port, B1 => 
                           n36286, B2 => REGISTERS_2_0_port, ZN => n35593);
   U195 : AOI22_X1 port map( A1 => n36287, A2 => REGISTERS_31_0_port, B1 => 
                           n36288, B2 => REGISTERS_3_0_port, ZN => n35594);
   U196 : AOI22_X1 port map( A1 => n36289, A2 => REGISTERS_8_0_port, B1 => 
                           n36290, B2 => REGISTERS_30_0_port, ZN => n35595);
   U197 : NAND4_X1 port map( A1 => n35592, A2 => n35593, A3 => n35594, A4 => 
                           n35595, ZN => n35596);
   U198 : AOI22_X1 port map( A1 => n36291, A2 => REGISTERS_29_0_port, B1 => 
                           n36292, B2 => REGISTERS_11_0_port, ZN => n35597);
   U199 : AOI22_X1 port map( A1 => n36293, A2 => REGISTERS_16_0_port, B1 => 
                           n36294, B2 => REGISTERS_1_0_port, ZN => n35598);
   U200 : AOI22_X1 port map( A1 => n36295, A2 => REGISTERS_24_0_port, B1 => 
                           n36296, B2 => REGISTERS_12_0_port, ZN => n35599);
   U201 : AOI22_X1 port map( A1 => n36297, A2 => REGISTERS_15_0_port, B1 => 
                           n36298, B2 => REGISTERS_20_0_port, ZN => n35600);
   U202 : NAND4_X1 port map( A1 => n35597, A2 => n35598, A3 => n35599, A4 => 
                           n35600, ZN => n35601);
   U203 : AOI22_X1 port map( A1 => n36268, A2 => REGISTERS_22_0_port, B1 => 
                           n36269, B2 => REGISTERS_5_0_port, ZN => n35602);
   U204 : AOI22_X1 port map( A1 => n36270, A2 => REGISTERS_21_0_port, B1 => 
                           n36271, B2 => REGISTERS_25_0_port, ZN => n35603);
   U205 : AOI222_X1 port map( A1 => n36272, A2 => REGISTERS_23_0_port, B1 => 
                           n36273, B2 => REGISTERS_17_0_port, C1 => n36274, C2 
                           => REGISTERS_19_0_port, ZN => n35604);
   U206 : NAND3_X1 port map( A1 => n35602, A2 => n35603, A3 => n35604, ZN => 
                           n35605);
   U207 : AOI22_X1 port map( A1 => n36275, A2 => REGISTERS_13_0_port, B1 => 
                           n36276, B2 => REGISTERS_14_0_port, ZN => n35606);
   U208 : AOI22_X1 port map( A1 => n36279, A2 => REGISTERS_28_0_port, B1 => 
                           n36280, B2 => REGISTERS_6_0_port, ZN => n35607);
   U209 : AOI22_X1 port map( A1 => n36281, A2 => REGISTERS_7_0_port, B1 => 
                           n36282, B2 => REGISTERS_26_0_port, ZN => n35608);
   U210 : NAND4_X1 port map( A1 => n35606, A2 => n36355, A3 => n35607, A4 => 
                           n35608, ZN => n35609);
   U211 : OR4_X1 port map( A1 => n35596, A2 => n35601, A3 => n35605, A4 => 
                           n35609, ZN => OUTA(0));
   U212 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_31_port, B1 => 
                           n36237, B2 => REGISTERS_14_31_port, ZN => n35610);
   U213 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_31_port, B1 => 
                           n36242, B2 => REGISTERS_4_31_port, ZN => n35611);
   U214 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_31_port, B1 => 
                           n36245, B2 => REGISTERS_22_31_port, ZN => n35612);
   U215 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_31_port, B1 => 
                           n36258, B2 => REGISTERS_9_31_port, ZN => n35613);
   U216 : NAND4_X1 port map( A1 => n35610, A2 => n35611, A3 => n35612, A4 => 
                           n35613, ZN => n35614);
   U217 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_31_port, B1 => 
                           n36263, B2 => REGISTERS_25_31_port, ZN => n35615);
   U218 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_31_port, B1 => 
                           n36264, B2 => REGISTERS_2_31_port, ZN => n35616);
   U219 : AOI22_X1 port map( A1 => n36855, A2 => REGISTERS_31_31_port, B1 => 
                           n36261, B2 => REGISTERS_13_31_port, ZN => n35617);
   U220 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_31_port, B1 => 
                           n36259, B2 => REGISTERS_8_31_port, ZN => n35618);
   U221 : NAND4_X1 port map( A1 => n35615, A2 => n35616, A3 => n35617, A4 => 
                           n35618, ZN => n35619);
   U222 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_31_port, B1 => 
                           n36256, B2 => REGISTERS_21_31_port, ZN => n35620);
   U223 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_31_port, B1 => 
                           n36252, B2 => REGISTERS_7_31_port, ZN => n35621);
   U224 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_31_port, B1 => 
                           n36249, B2 => REGISTERS_5_31_port, C1 => n36247, C2 
                           => REGISTERS_18_31_port, ZN => n35622);
   U225 : NAND3_X1 port map( A1 => n35620, A2 => n35621, A3 => n35622, ZN => 
                           n35623);
   U226 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_31_port, B1 => 
                           n36246, B2 => REGISTERS_19_31_port, ZN => n35624);
   U227 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_31_port, B1 => 
                           n36257, B2 => REGISTERS_23_31_port, ZN => n35625);
   U228 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_31_port, B1 => 
                           n36241, B2 => REGISTERS_10_31_port, ZN => n35626);
   U229 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_31_port, B1 => 
                           n36266, B2 => REGISTERS_27_31_port, ZN => n35627);
   U230 : NAND4_X1 port map( A1 => n35624, A2 => n35625, A3 => n35626, A4 => 
                           n35627, ZN => n35628);
   U231 : OR4_X1 port map( A1 => n35614, A2 => n35619, A3 => n35623, A4 => 
                           n35628, ZN => OUTB(31));
   U232 : AOI22_X1 port map( A1 => n36781, A2 => REGISTERS_9_31_port, B1 => 
                           n36782, B2 => REGISTERS_10_31_port, ZN => n35629);
   U233 : AOI22_X1 port map( A1 => n36783, A2 => REGISTERS_18_31_port, B1 => 
                           n36784, B2 => REGISTERS_2_31_port, ZN => n35630);
   U234 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_31_port, B1 => 
                           n36785, B2 => REGISTERS_31_31_port, ZN => n35631);
   U235 : AOI22_X1 port map( A1 => n36787, A2 => REGISTERS_8_31_port, B1 => 
                           n36788, B2 => REGISTERS_30_31_port, ZN => n35632);
   U236 : NAND4_X1 port map( A1 => n35629, A2 => n35630, A3 => n35631, A4 => 
                           n35632, ZN => n35633);
   U237 : AOI22_X1 port map( A1 => n36793, A2 => REGISTERS_29_31_port, B1 => 
                           n36794, B2 => REGISTERS_11_31_port, ZN => n35634);
   U238 : AOI22_X1 port map( A1 => n36795, A2 => REGISTERS_16_31_port, B1 => 
                           n36796, B2 => REGISTERS_1_31_port, ZN => n35635);
   U239 : AOI22_X1 port map( A1 => n36797, A2 => REGISTERS_24_31_port, B1 => 
                           n36798, B2 => REGISTERS_12_31_port, ZN => n35636);
   U240 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_31_port, B1 => 
                           n36799, B2 => REGISTERS_15_31_port, ZN => n35637);
   U241 : NAND4_X1 port map( A1 => n35634, A2 => n35635, A3 => n35636, A4 => 
                           n35637, ZN => n35638);
   U242 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_31_port, B1 => 
                           n36758, B2 => REGISTERS_22_31_port, ZN => n35639);
   U243 : AOI22_X1 port map( A1 => n36760, A2 => REGISTERS_21_31_port, B1 => 
                           n36761, B2 => REGISTERS_25_31_port, ZN => n35640);
   U244 : AOI222_X1 port map( A1 => n36763, A2 => REGISTERS_17_31_port, B1 => 
                           n36762, B2 => REGISTERS_23_31_port, C1 => n36764, C2
                           => REGISTERS_19_31_port, ZN => n35641);
   U245 : NAND3_X1 port map( A1 => n35639, A2 => n35640, A3 => n35641, ZN => 
                           n35642);
   U246 : AOI22_X1 port map( A1 => n36769, A2 => REGISTERS_13_31_port, B1 => 
                           n36770, B2 => REGISTERS_14_31_port, ZN => n35643);
   U247 : AOI22_X1 port map( A1 => n36771, A2 => REGISTERS_4_31_port, B1 => 
                           n36772, B2 => REGISTERS_27_31_port, ZN => n35644);
   U248 : AOI22_X1 port map( A1 => n36773, A2 => REGISTERS_28_31_port, B1 => 
                           n36774, B2 => REGISTERS_6_31_port, ZN => n35645);
   U249 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_31_port, B1 => 
                           n36775, B2 => REGISTERS_7_31_port, ZN => n35646);
   U250 : NAND4_X1 port map( A1 => n35643, A2 => n35644, A3 => n35645, A4 => 
                           n35646, ZN => n35647);
   U251 : OR4_X1 port map( A1 => n35633, A2 => n35638, A3 => n35642, A4 => 
                           n35647, ZN => OUTA(31));
   U252 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_30_port, B1 => 
                           n36237, B2 => REGISTERS_14_30_port, ZN => n35648);
   U253 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_30_port, B1 => 
                           n36242, B2 => REGISTERS_4_30_port, ZN => n35649);
   U254 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_30_port, B1 => 
                           n36245, B2 => REGISTERS_22_30_port, ZN => n35650);
   U255 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_30_port, B1 => 
                           n36258, B2 => REGISTERS_9_30_port, ZN => n35651);
   U256 : NAND4_X1 port map( A1 => n35648, A2 => n35649, A3 => n35650, A4 => 
                           n35651, ZN => n35652);
   U257 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_30_port, B1 => 
                           n36263, B2 => REGISTERS_25_30_port, ZN => n35653);
   U258 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_30_port, B1 => 
                           n36264, B2 => REGISTERS_2_30_port, ZN => n35654);
   U259 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_30_port, B1 => 
                           n36261, B2 => REGISTERS_13_30_port, ZN => n35655);
   U260 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_30_port, B1 => 
                           n36259, B2 => REGISTERS_8_30_port, ZN => n35656);
   U261 : NAND4_X1 port map( A1 => n35653, A2 => n35654, A3 => n35655, A4 => 
                           n35656, ZN => n35657);
   U262 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_30_port, B1 => 
                           n36256, B2 => REGISTERS_21_30_port, ZN => n35658);
   U263 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_30_port, B1 => 
                           n36252, B2 => REGISTERS_7_30_port, ZN => n35659);
   U264 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_30_port, B1 => 
                           n36249, B2 => REGISTERS_5_30_port, C1 => n36247, C2 
                           => REGISTERS_18_30_port, ZN => n35660);
   U265 : NAND3_X1 port map( A1 => n35658, A2 => n35659, A3 => n35660, ZN => 
                           n35661);
   U266 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_30_port, B1 => 
                           n36246, B2 => REGISTERS_19_30_port, ZN => n35662);
   U267 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_30_port, B1 => 
                           n36257, B2 => REGISTERS_23_30_port, ZN => n35663);
   U268 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_30_port, B1 => 
                           n36241, B2 => REGISTERS_10_30_port, ZN => n35664);
   U269 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_30_port, B1 => 
                           n36266, B2 => REGISTERS_27_30_port, ZN => n35665);
   U270 : NAND4_X1 port map( A1 => n35662, A2 => n35663, A3 => n35664, A4 => 
                           n35665, ZN => n35666);
   U271 : OR4_X1 port map( A1 => n35652, A2 => n35657, A3 => n35661, A4 => 
                           n35666, ZN => OUTB(30));
   U272 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_29_port, B1 => 
                           n36237, B2 => REGISTERS_14_29_port, ZN => n35667);
   U273 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_29_port, B1 => 
                           n36242, B2 => REGISTERS_4_29_port, ZN => n35668);
   U274 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_29_port, B1 => 
                           n36245, B2 => REGISTERS_22_29_port, ZN => n35669);
   U275 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_29_port, B1 => 
                           n36258, B2 => REGISTERS_9_29_port, ZN => n35670);
   U276 : NAND4_X1 port map( A1 => n35667, A2 => n35668, A3 => n35669, A4 => 
                           n35670, ZN => n35671);
   U277 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_29_port, B1 => 
                           n36263, B2 => REGISTERS_25_29_port, ZN => n35672);
   U278 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_29_port, B1 => 
                           n36264, B2 => REGISTERS_2_29_port, ZN => n35673);
   U279 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_29_port, B1 => 
                           n36261, B2 => REGISTERS_13_29_port, ZN => n35674);
   U280 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_29_port, B1 => 
                           n36259, B2 => REGISTERS_8_29_port, ZN => n35675);
   U281 : NAND4_X1 port map( A1 => n35672, A2 => n35673, A3 => n35674, A4 => 
                           n35675, ZN => n35676);
   U282 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_29_port, B1 => 
                           n36256, B2 => REGISTERS_21_29_port, ZN => n35677);
   U283 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_29_port, B1 => 
                           n36252, B2 => REGISTERS_7_29_port, ZN => n35678);
   U284 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_29_port, B1 => 
                           n36249, B2 => REGISTERS_5_29_port, C1 => n36247, C2 
                           => REGISTERS_18_29_port, ZN => n35679);
   U285 : NAND3_X1 port map( A1 => n35677, A2 => n35678, A3 => n35679, ZN => 
                           n35680);
   U286 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_29_port, B1 => 
                           n36246, B2 => REGISTERS_19_29_port, ZN => n35681);
   U287 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_29_port, B1 => 
                           n36257, B2 => REGISTERS_23_29_port, ZN => n35682);
   U288 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_29_port, B1 => 
                           n36241, B2 => REGISTERS_10_29_port, ZN => n35683);
   U289 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_29_port, B1 => 
                           n36266, B2 => REGISTERS_27_29_port, ZN => n35684);
   U290 : NAND4_X1 port map( A1 => n35681, A2 => n35682, A3 => n35683, A4 => 
                           n35684, ZN => n35685);
   U291 : OR4_X1 port map( A1 => n35671, A2 => n35676, A3 => n35680, A4 => 
                           n35685, ZN => OUTB(29));
   U292 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_28_port, B1 => 
                           n36237, B2 => REGISTERS_14_28_port, ZN => n35686);
   U293 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_28_port, B1 => 
                           n36242, B2 => REGISTERS_4_28_port, ZN => n35687);
   U294 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_28_port, B1 => 
                           n36245, B2 => REGISTERS_22_28_port, ZN => n35688);
   U295 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_28_port, B1 => 
                           n36258, B2 => REGISTERS_9_28_port, ZN => n35689);
   U296 : NAND4_X1 port map( A1 => n35686, A2 => n35687, A3 => n35688, A4 => 
                           n35689, ZN => n35690);
   U297 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_28_port, B1 => 
                           n36263, B2 => REGISTERS_25_28_port, ZN => n35691);
   U298 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_28_port, B1 => 
                           n36264, B2 => REGISTERS_2_28_port, ZN => n35692);
   U299 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_28_port, B1 => 
                           n36261, B2 => REGISTERS_13_28_port, ZN => n35693);
   U300 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_28_port, B1 => 
                           n36259, B2 => REGISTERS_8_28_port, ZN => n35694);
   U301 : NAND4_X1 port map( A1 => n35691, A2 => n35692, A3 => n35693, A4 => 
                           n35694, ZN => n35695);
   U302 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_28_port, B1 => 
                           n36256, B2 => REGISTERS_21_28_port, ZN => n35696);
   U303 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_28_port, B1 => 
                           n36252, B2 => REGISTERS_7_28_port, ZN => n35697);
   U304 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_28_port, B1 => 
                           n36249, B2 => REGISTERS_5_28_port, C1 => n36247, C2 
                           => REGISTERS_18_28_port, ZN => n35698);
   U305 : NAND3_X1 port map( A1 => n35696, A2 => n35697, A3 => n35698, ZN => 
                           n35699);
   U306 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_28_port, B1 => 
                           n36246, B2 => REGISTERS_19_28_port, ZN => n35700);
   U307 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_28_port, B1 => 
                           n36257, B2 => REGISTERS_23_28_port, ZN => n35701);
   U308 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_28_port, B1 => 
                           n36241, B2 => REGISTERS_10_28_port, ZN => n35702);
   U309 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_28_port, B1 => 
                           n36266, B2 => REGISTERS_27_28_port, ZN => n35703);
   U310 : NAND4_X1 port map( A1 => n35700, A2 => n35701, A3 => n35702, A4 => 
                           n35703, ZN => n35704);
   U311 : OR4_X1 port map( A1 => n35690, A2 => n35695, A3 => n35699, A4 => 
                           n35704, ZN => OUTB(28));
   U312 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_27_port, B1 => 
                           n36237, B2 => REGISTERS_14_27_port, ZN => n35705);
   U313 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_27_port, B1 => 
                           n36242, B2 => REGISTERS_4_27_port, ZN => n35706);
   U314 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_27_port, B1 => 
                           n36245, B2 => REGISTERS_22_27_port, ZN => n35707);
   U315 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_27_port, B1 => 
                           n36258, B2 => REGISTERS_9_27_port, ZN => n35708);
   U316 : NAND4_X1 port map( A1 => n35705, A2 => n35706, A3 => n35707, A4 => 
                           n35708, ZN => n35709);
   U317 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_27_port, B1 => 
                           n36263, B2 => REGISTERS_25_27_port, ZN => n35710);
   U318 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_27_port, B1 => 
                           n36264, B2 => REGISTERS_2_27_port, ZN => n35711);
   U319 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_27_port, B1 => 
                           n36261, B2 => REGISTERS_13_27_port, ZN => n35712);
   U320 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_27_port, B1 => 
                           n36259, B2 => REGISTERS_8_27_port, ZN => n35713);
   U321 : NAND4_X1 port map( A1 => n35710, A2 => n35711, A3 => n35712, A4 => 
                           n35713, ZN => n35714);
   U322 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_27_port, B1 => 
                           n36256, B2 => REGISTERS_21_27_port, ZN => n35715);
   U323 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_27_port, B1 => 
                           n36252, B2 => REGISTERS_7_27_port, ZN => n35716);
   U324 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_27_port, B1 => 
                           n36249, B2 => REGISTERS_5_27_port, C1 => n36247, C2 
                           => REGISTERS_18_27_port, ZN => n35717);
   U325 : NAND3_X1 port map( A1 => n35715, A2 => n35716, A3 => n35717, ZN => 
                           n35718);
   U326 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_27_port, B1 => 
                           n36246, B2 => REGISTERS_19_27_port, ZN => n35719);
   U327 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_27_port, B1 => 
                           n36257, B2 => REGISTERS_23_27_port, ZN => n35720);
   U328 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_27_port, B1 => 
                           n36241, B2 => REGISTERS_10_27_port, ZN => n35721);
   U329 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_27_port, B1 => 
                           n36266, B2 => REGISTERS_27_27_port, ZN => n35722);
   U330 : NAND4_X1 port map( A1 => n35719, A2 => n35720, A3 => n35721, A4 => 
                           n35722, ZN => n35723);
   U331 : OR4_X1 port map( A1 => n35709, A2 => n35714, A3 => n35718, A4 => 
                           n35723, ZN => OUTB(27));
   U332 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_26_port, B1 => 
                           n36237, B2 => REGISTERS_14_26_port, ZN => n35724);
   U333 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_26_port, B1 => 
                           n36242, B2 => REGISTERS_4_26_port, ZN => n35725);
   U334 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_26_port, B1 => 
                           n36245, B2 => REGISTERS_22_26_port, ZN => n35726);
   U335 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_26_port, B1 => 
                           n36258, B2 => REGISTERS_9_26_port, ZN => n35727);
   U336 : NAND4_X1 port map( A1 => n35724, A2 => n35725, A3 => n35726, A4 => 
                           n35727, ZN => n35728);
   U337 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_26_port, B1 => 
                           n36263, B2 => REGISTERS_25_26_port, ZN => n35729);
   U338 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_26_port, B1 => 
                           n36264, B2 => REGISTERS_2_26_port, ZN => n35730);
   U339 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_26_port, B1 => 
                           n36261, B2 => REGISTERS_13_26_port, ZN => n35731);
   U340 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_26_port, B1 => 
                           n36259, B2 => REGISTERS_8_26_port, ZN => n35732);
   U341 : NAND4_X1 port map( A1 => n35729, A2 => n35730, A3 => n35731, A4 => 
                           n35732, ZN => n35733);
   U342 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_26_port, B1 => 
                           n36256, B2 => REGISTERS_21_26_port, ZN => n35734);
   U343 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_26_port, B1 => 
                           n36252, B2 => REGISTERS_7_26_port, ZN => n35735);
   U344 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_26_port, B1 => 
                           n36249, B2 => REGISTERS_5_26_port, C1 => n36247, C2 
                           => REGISTERS_18_26_port, ZN => n35736);
   U345 : NAND3_X1 port map( A1 => n35734, A2 => n35735, A3 => n35736, ZN => 
                           n35737);
   U346 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_26_port, B1 => 
                           n36246, B2 => REGISTERS_19_26_port, ZN => n35738);
   U347 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_26_port, B1 => 
                           n36257, B2 => REGISTERS_23_26_port, ZN => n35739);
   U348 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_26_port, B1 => 
                           n36241, B2 => REGISTERS_10_26_port, ZN => n35740);
   U349 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_26_port, B1 => 
                           n36266, B2 => REGISTERS_27_26_port, ZN => n35741);
   U350 : NAND4_X1 port map( A1 => n35738, A2 => n35739, A3 => n35740, A4 => 
                           n35741, ZN => n35742);
   U351 : OR4_X1 port map( A1 => n35728, A2 => n35733, A3 => n35737, A4 => 
                           n35742, ZN => OUTB(26));
   U352 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_25_port, B1 => 
                           n36237, B2 => REGISTERS_14_25_port, ZN => n35743);
   U353 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_25_port, B1 => 
                           n36242, B2 => REGISTERS_4_25_port, ZN => n35744);
   U354 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_25_port, B1 => 
                           n36245, B2 => REGISTERS_22_25_port, ZN => n35745);
   U355 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_25_port, B1 => 
                           n36258, B2 => REGISTERS_9_25_port, ZN => n35746);
   U356 : NAND4_X1 port map( A1 => n35743, A2 => n35744, A3 => n35745, A4 => 
                           n35746, ZN => n35747);
   U357 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_25_port, B1 => 
                           n36263, B2 => REGISTERS_25_25_port, ZN => n35748);
   U358 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_25_port, B1 => 
                           n36264, B2 => REGISTERS_2_25_port, ZN => n35749);
   U359 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_25_port, B1 => 
                           n36261, B2 => REGISTERS_13_25_port, ZN => n35750);
   U360 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_25_port, B1 => 
                           n36259, B2 => REGISTERS_8_25_port, ZN => n35751);
   U361 : NAND4_X1 port map( A1 => n35748, A2 => n35749, A3 => n35750, A4 => 
                           n35751, ZN => n35752);
   U362 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_25_port, B1 => 
                           n36256, B2 => REGISTERS_21_25_port, ZN => n35753);
   U363 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_25_port, B1 => 
                           n36252, B2 => REGISTERS_7_25_port, ZN => n35754);
   U364 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_25_port, B1 => 
                           n36249, B2 => REGISTERS_5_25_port, C1 => n36247, C2 
                           => REGISTERS_18_25_port, ZN => n35755);
   U365 : NAND3_X1 port map( A1 => n35753, A2 => n35754, A3 => n35755, ZN => 
                           n35756);
   U366 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_25_port, B1 => 
                           n36246, B2 => REGISTERS_19_25_port, ZN => n35757);
   U367 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_25_port, B1 => 
                           n36257, B2 => REGISTERS_23_25_port, ZN => n35758);
   U368 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_25_port, B1 => 
                           n36241, B2 => REGISTERS_10_25_port, ZN => n35759);
   U369 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_25_port, B1 => 
                           n36266, B2 => REGISTERS_27_25_port, ZN => n35760);
   U370 : NAND4_X1 port map( A1 => n35757, A2 => n35758, A3 => n35759, A4 => 
                           n35760, ZN => n35761);
   U371 : OR4_X1 port map( A1 => n35747, A2 => n35752, A3 => n35756, A4 => 
                           n35761, ZN => OUTB(25));
   U372 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_24_port, B1 => 
                           n36237, B2 => REGISTERS_14_24_port, ZN => n35762);
   U373 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_24_port, B1 => 
                           n36242, B2 => REGISTERS_4_24_port, ZN => n35763);
   U374 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_24_port, B1 => 
                           n36245, B2 => REGISTERS_22_24_port, ZN => n35764);
   U375 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_24_port, B1 => 
                           n36258, B2 => REGISTERS_9_24_port, ZN => n35765);
   U376 : NAND4_X1 port map( A1 => n35762, A2 => n35763, A3 => n35764, A4 => 
                           n35765, ZN => n35766);
   U377 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_24_port, B1 => 
                           n36263, B2 => REGISTERS_25_24_port, ZN => n35767);
   U378 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_24_port, B1 => 
                           n36264, B2 => REGISTERS_2_24_port, ZN => n35768);
   U379 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_24_port, B1 => 
                           n36261, B2 => REGISTERS_13_24_port, ZN => n35769);
   U380 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_24_port, B1 => 
                           n36259, B2 => REGISTERS_8_24_port, ZN => n35770);
   U381 : NAND4_X1 port map( A1 => n35767, A2 => n35768, A3 => n35769, A4 => 
                           n35770, ZN => n35771);
   U382 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_24_port, B1 => 
                           n36256, B2 => REGISTERS_21_24_port, ZN => n35772);
   U383 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_24_port, B1 => 
                           n36252, B2 => REGISTERS_7_24_port, ZN => n35773);
   U384 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_24_port, B1 => 
                           n36249, B2 => REGISTERS_5_24_port, C1 => n36247, C2 
                           => REGISTERS_18_24_port, ZN => n35774);
   U385 : NAND3_X1 port map( A1 => n35772, A2 => n35773, A3 => n35774, ZN => 
                           n35775);
   U386 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_24_port, B1 => 
                           n36246, B2 => REGISTERS_19_24_port, ZN => n35776);
   U387 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_24_port, B1 => 
                           n36257, B2 => REGISTERS_23_24_port, ZN => n35777);
   U388 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_24_port, B1 => 
                           n36241, B2 => REGISTERS_10_24_port, ZN => n35778);
   U389 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_24_port, B1 => 
                           n36266, B2 => REGISTERS_27_24_port, ZN => n35779);
   U390 : NAND4_X1 port map( A1 => n35776, A2 => n35777, A3 => n35778, A4 => 
                           n35779, ZN => n35780);
   U391 : OR4_X1 port map( A1 => n35766, A2 => n35771, A3 => n35775, A4 => 
                           n35780, ZN => OUTB(24));
   U392 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_23_port, B1 => 
                           n36237, B2 => REGISTERS_14_23_port, ZN => n35781);
   U393 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_23_port, B1 => 
                           n36242, B2 => REGISTERS_4_23_port, ZN => n35782);
   U394 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_23_port, B1 => 
                           n36245, B2 => REGISTERS_22_23_port, ZN => n35783);
   U395 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_23_port, B1 => 
                           n36258, B2 => REGISTERS_9_23_port, ZN => n35784);
   U396 : NAND4_X1 port map( A1 => n35781, A2 => n35782, A3 => n35783, A4 => 
                           n35784, ZN => n35785);
   U397 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_23_port, B1 => 
                           n36263, B2 => REGISTERS_25_23_port, ZN => n35786);
   U398 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_23_port, B1 => 
                           n36264, B2 => REGISTERS_2_23_port, ZN => n35787);
   U399 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_23_port, B1 => 
                           n36261, B2 => REGISTERS_13_23_port, ZN => n35788);
   U400 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_23_port, B1 => 
                           n36259, B2 => REGISTERS_8_23_port, ZN => n35789);
   U401 : NAND4_X1 port map( A1 => n35786, A2 => n35787, A3 => n35788, A4 => 
                           n35789, ZN => n35790);
   U402 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_23_port, B1 => 
                           n36256, B2 => REGISTERS_21_23_port, ZN => n35791);
   U403 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_23_port, B1 => 
                           n36252, B2 => REGISTERS_7_23_port, ZN => n35792);
   U404 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_23_port, B1 => 
                           n36249, B2 => REGISTERS_5_23_port, C1 => n36247, C2 
                           => REGISTERS_18_23_port, ZN => n35793);
   U405 : NAND3_X1 port map( A1 => n35791, A2 => n35792, A3 => n35793, ZN => 
                           n35794);
   U406 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_23_port, B1 => 
                           n36246, B2 => REGISTERS_19_23_port, ZN => n35795);
   U407 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_23_port, B1 => 
                           n36257, B2 => REGISTERS_23_23_port, ZN => n35796);
   U408 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_23_port, B1 => 
                           n36241, B2 => REGISTERS_10_23_port, ZN => n35797);
   U409 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_23_port, B1 => 
                           n36266, B2 => REGISTERS_27_23_port, ZN => n35798);
   U410 : NAND4_X1 port map( A1 => n35795, A2 => n35796, A3 => n35797, A4 => 
                           n35798, ZN => n35799);
   U411 : OR4_X1 port map( A1 => n35785, A2 => n35790, A3 => n35794, A4 => 
                           n35799, ZN => OUTB(23));
   U412 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_22_port, B1 => 
                           n36237, B2 => REGISTERS_14_22_port, ZN => n35800);
   U413 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_22_port, B1 => 
                           n36242, B2 => REGISTERS_4_22_port, ZN => n35801);
   U414 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_22_port, B1 => 
                           n36245, B2 => REGISTERS_22_22_port, ZN => n35802);
   U415 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_22_port, B1 => 
                           n36258, B2 => REGISTERS_9_22_port, ZN => n35803);
   U416 : NAND4_X1 port map( A1 => n35800, A2 => n35801, A3 => n35802, A4 => 
                           n35803, ZN => n35804);
   U417 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_22_port, B1 => 
                           n36263, B2 => REGISTERS_25_22_port, ZN => n35805);
   U418 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_22_port, B1 => 
                           n36264, B2 => REGISTERS_2_22_port, ZN => n35806);
   U419 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_22_port, B1 => 
                           n36261, B2 => REGISTERS_13_22_port, ZN => n35807);
   U420 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_22_port, B1 => 
                           n36259, B2 => REGISTERS_8_22_port, ZN => n35808);
   U421 : NAND4_X1 port map( A1 => n35805, A2 => n35806, A3 => n35807, A4 => 
                           n35808, ZN => n35809);
   U422 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_22_port, B1 => 
                           n36256, B2 => REGISTERS_21_22_port, ZN => n35810);
   U423 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_22_port, B1 => 
                           n36252, B2 => REGISTERS_7_22_port, ZN => n35811);
   U424 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_22_port, B1 => 
                           n36249, B2 => REGISTERS_5_22_port, C1 => n36247, C2 
                           => REGISTERS_18_22_port, ZN => n35812);
   U425 : NAND3_X1 port map( A1 => n35810, A2 => n35811, A3 => n35812, ZN => 
                           n35813);
   U426 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_22_port, B1 => 
                           n36246, B2 => REGISTERS_19_22_port, ZN => n35814);
   U427 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_22_port, B1 => 
                           n36257, B2 => REGISTERS_23_22_port, ZN => n35815);
   U428 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_22_port, B1 => 
                           n36241, B2 => REGISTERS_10_22_port, ZN => n35816);
   U429 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_22_port, B1 => 
                           n36266, B2 => REGISTERS_27_22_port, ZN => n35817);
   U430 : NAND4_X1 port map( A1 => n35814, A2 => n35815, A3 => n35816, A4 => 
                           n35817, ZN => n35818);
   U431 : OR4_X1 port map( A1 => n35804, A2 => n35809, A3 => n35813, A4 => 
                           n35818, ZN => OUTB(22));
   U432 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_21_port, B1 => 
                           n36237, B2 => REGISTERS_14_21_port, ZN => n35819);
   U433 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_21_port, B1 => 
                           n36242, B2 => REGISTERS_4_21_port, ZN => n35820);
   U434 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_21_port, B1 => 
                           n36245, B2 => REGISTERS_22_21_port, ZN => n35821);
   U435 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_21_port, B1 => 
                           n36258, B2 => REGISTERS_9_21_port, ZN => n35822);
   U436 : NAND4_X1 port map( A1 => n35819, A2 => n35820, A3 => n35821, A4 => 
                           n35822, ZN => n35823);
   U437 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_21_port, B1 => 
                           n36263, B2 => REGISTERS_25_21_port, ZN => n35824);
   U438 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_21_port, B1 => 
                           n36264, B2 => REGISTERS_2_21_port, ZN => n35825);
   U439 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_21_port, B1 => 
                           n36261, B2 => REGISTERS_13_21_port, ZN => n35826);
   U440 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_21_port, B1 => 
                           n36259, B2 => REGISTERS_8_21_port, ZN => n35827);
   U441 : NAND4_X1 port map( A1 => n35824, A2 => n35825, A3 => n35826, A4 => 
                           n35827, ZN => n35828);
   U442 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_21_port, B1 => 
                           n36256, B2 => REGISTERS_21_21_port, ZN => n35829);
   U443 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_21_port, B1 => 
                           n36252, B2 => REGISTERS_7_21_port, ZN => n35830);
   U444 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_21_port, B1 => 
                           n36249, B2 => REGISTERS_5_21_port, C1 => n36247, C2 
                           => REGISTERS_18_21_port, ZN => n35831);
   U445 : NAND3_X1 port map( A1 => n35829, A2 => n35830, A3 => n35831, ZN => 
                           n35832);
   U446 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_21_port, B1 => 
                           n36246, B2 => REGISTERS_19_21_port, ZN => n35833);
   U447 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_21_port, B1 => 
                           n36257, B2 => REGISTERS_23_21_port, ZN => n35834);
   U448 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_21_port, B1 => 
                           n36241, B2 => REGISTERS_10_21_port, ZN => n35835);
   U449 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_21_port, B1 => 
                           n36266, B2 => REGISTERS_27_21_port, ZN => n35836);
   U450 : NAND4_X1 port map( A1 => n35833, A2 => n35834, A3 => n35835, A4 => 
                           n35836, ZN => n35837);
   U451 : OR4_X1 port map( A1 => n35823, A2 => n35828, A3 => n35832, A4 => 
                           n35837, ZN => OUTB(21));
   U452 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_20_port, B1 => 
                           n36237, B2 => REGISTERS_14_20_port, ZN => n35838);
   U453 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_20_port, B1 => 
                           n36242, B2 => REGISTERS_4_20_port, ZN => n35839);
   U454 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_20_port, B1 => 
                           n36245, B2 => REGISTERS_22_20_port, ZN => n35840);
   U455 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_20_port, B1 => 
                           n36258, B2 => REGISTERS_9_20_port, ZN => n35841);
   U456 : NAND4_X1 port map( A1 => n35838, A2 => n35839, A3 => n35840, A4 => 
                           n35841, ZN => n35842);
   U457 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_20_port, B1 => 
                           n36263, B2 => REGISTERS_25_20_port, ZN => n35843);
   U458 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_20_port, B1 => 
                           n36264, B2 => REGISTERS_2_20_port, ZN => n35844);
   U459 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_20_port, B1 => 
                           n36261, B2 => REGISTERS_13_20_port, ZN => n35845);
   U460 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_20_port, B1 => 
                           n36259, B2 => REGISTERS_8_20_port, ZN => n35846);
   U461 : NAND4_X1 port map( A1 => n35843, A2 => n35844, A3 => n35845, A4 => 
                           n35846, ZN => n35847);
   U462 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_20_port, B1 => 
                           n36256, B2 => REGISTERS_21_20_port, ZN => n35848);
   U463 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_20_port, B1 => 
                           n36252, B2 => REGISTERS_7_20_port, ZN => n35849);
   U464 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_20_port, B1 => 
                           n36249, B2 => REGISTERS_5_20_port, C1 => n36247, C2 
                           => REGISTERS_18_20_port, ZN => n35850);
   U465 : NAND3_X1 port map( A1 => n35848, A2 => n35849, A3 => n35850, ZN => 
                           n35851);
   U466 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_20_port, B1 => 
                           n36246, B2 => REGISTERS_19_20_port, ZN => n35852);
   U467 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_20_port, B1 => 
                           n36257, B2 => REGISTERS_23_20_port, ZN => n35853);
   U468 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_20_port, B1 => 
                           n36241, B2 => REGISTERS_10_20_port, ZN => n35854);
   U469 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_20_port, B1 => 
                           n36266, B2 => REGISTERS_27_20_port, ZN => n35855);
   U470 : NAND4_X1 port map( A1 => n35852, A2 => n35853, A3 => n35854, A4 => 
                           n35855, ZN => n35856);
   U471 : OR4_X1 port map( A1 => n35842, A2 => n35847, A3 => n35851, A4 => 
                           n35856, ZN => OUTB(20));
   U472 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_19_port, B1 => 
                           n36237, B2 => REGISTERS_14_19_port, ZN => n35857);
   U473 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_19_port, B1 => 
                           n36242, B2 => REGISTERS_4_19_port, ZN => n35858);
   U474 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_19_port, B1 => 
                           n36245, B2 => REGISTERS_22_19_port, ZN => n35859);
   U475 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_19_port, B1 => 
                           n36258, B2 => REGISTERS_9_19_port, ZN => n35860);
   U476 : NAND4_X1 port map( A1 => n35857, A2 => n35858, A3 => n35859, A4 => 
                           n35860, ZN => n35861);
   U477 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_19_port, B1 => 
                           n36263, B2 => REGISTERS_25_19_port, ZN => n35862);
   U478 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_19_port, B1 => 
                           n36264, B2 => REGISTERS_2_19_port, ZN => n35863);
   U479 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_19_port, B1 => 
                           n36261, B2 => REGISTERS_13_19_port, ZN => n35864);
   U480 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_19_port, B1 => 
                           n36259, B2 => REGISTERS_8_19_port, ZN => n35865);
   U481 : NAND4_X1 port map( A1 => n35862, A2 => n35863, A3 => n35864, A4 => 
                           n35865, ZN => n35866);
   U482 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_19_port, B1 => 
                           n36256, B2 => REGISTERS_21_19_port, ZN => n35867);
   U483 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_19_port, B1 => 
                           n36252, B2 => REGISTERS_7_19_port, ZN => n35868);
   U484 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_19_port, B1 => 
                           n36249, B2 => REGISTERS_5_19_port, C1 => n36247, C2 
                           => REGISTERS_18_19_port, ZN => n35869);
   U485 : NAND3_X1 port map( A1 => n35867, A2 => n35868, A3 => n35869, ZN => 
                           n35870);
   U486 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_19_port, B1 => 
                           n36246, B2 => REGISTERS_19_19_port, ZN => n35871);
   U487 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_19_port, B1 => 
                           n36257, B2 => REGISTERS_23_19_port, ZN => n35872);
   U488 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_19_port, B1 => 
                           n36241, B2 => REGISTERS_10_19_port, ZN => n35873);
   U489 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_19_port, B1 => 
                           n36266, B2 => REGISTERS_27_19_port, ZN => n35874);
   U490 : NAND4_X1 port map( A1 => n35871, A2 => n35872, A3 => n35873, A4 => 
                           n35874, ZN => n35875);
   U491 : OR4_X1 port map( A1 => n35861, A2 => n35866, A3 => n35870, A4 => 
                           n35875, ZN => OUTB(19));
   U492 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_18_port, B1 => 
                           n36237, B2 => REGISTERS_14_18_port, ZN => n35876);
   U493 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_18_port, B1 => 
                           n36242, B2 => REGISTERS_4_18_port, ZN => n35877);
   U494 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_18_port, B1 => 
                           n36245, B2 => REGISTERS_22_18_port, ZN => n35878);
   U495 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_18_port, B1 => 
                           n36258, B2 => REGISTERS_9_18_port, ZN => n35879);
   U496 : NAND4_X1 port map( A1 => n35876, A2 => n35877, A3 => n35878, A4 => 
                           n35879, ZN => n35880);
   U497 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_18_port, B1 => 
                           n36263, B2 => REGISTERS_25_18_port, ZN => n35881);
   U498 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_18_port, B1 => 
                           n36264, B2 => REGISTERS_2_18_port, ZN => n35882);
   U499 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_18_port, B1 => 
                           n36261, B2 => REGISTERS_13_18_port, ZN => n35883);
   U500 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_18_port, B1 => 
                           n36259, B2 => REGISTERS_8_18_port, ZN => n35884);
   U501 : NAND4_X1 port map( A1 => n35881, A2 => n35882, A3 => n35883, A4 => 
                           n35884, ZN => n35885);
   U502 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_18_port, B1 => 
                           n36256, B2 => REGISTERS_21_18_port, ZN => n35886);
   U503 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_18_port, B1 => 
                           n36252, B2 => REGISTERS_7_18_port, ZN => n35887);
   U504 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_18_port, B1 => 
                           n36249, B2 => REGISTERS_5_18_port, C1 => n36247, C2 
                           => REGISTERS_18_18_port, ZN => n35888);
   U505 : NAND3_X1 port map( A1 => n35886, A2 => n35887, A3 => n35888, ZN => 
                           n35889);
   U506 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_18_port, B1 => 
                           n36246, B2 => REGISTERS_19_18_port, ZN => n35890);
   U507 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_18_port, B1 => 
                           n36257, B2 => REGISTERS_23_18_port, ZN => n35891);
   U508 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_18_port, B1 => 
                           n36241, B2 => REGISTERS_10_18_port, ZN => n35892);
   U509 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_18_port, B1 => 
                           n36266, B2 => REGISTERS_27_18_port, ZN => n35893);
   U510 : NAND4_X1 port map( A1 => n35890, A2 => n35891, A3 => n35892, A4 => 
                           n35893, ZN => n35894);
   U511 : OR4_X1 port map( A1 => n35880, A2 => n35885, A3 => n35889, A4 => 
                           n35894, ZN => OUTB(18));
   U512 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_17_port, B1 => 
                           n36237, B2 => REGISTERS_14_17_port, ZN => n35895);
   U513 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_17_port, B1 => 
                           n36242, B2 => REGISTERS_4_17_port, ZN => n35896);
   U514 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_17_port, B1 => 
                           n36245, B2 => REGISTERS_22_17_port, ZN => n35897);
   U515 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_17_port, B1 => 
                           n36258, B2 => REGISTERS_9_17_port, ZN => n35898);
   U516 : NAND4_X1 port map( A1 => n35895, A2 => n35896, A3 => n35897, A4 => 
                           n35898, ZN => n35899);
   U517 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_17_port, B1 => 
                           n36263, B2 => REGISTERS_25_17_port, ZN => n35900);
   U518 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_17_port, B1 => 
                           n36264, B2 => REGISTERS_2_17_port, ZN => n35901);
   U519 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_17_port, B1 => 
                           n36261, B2 => REGISTERS_13_17_port, ZN => n35902);
   U520 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_17_port, B1 => 
                           n36259, B2 => REGISTERS_8_17_port, ZN => n35903);
   U521 : NAND4_X1 port map( A1 => n35900, A2 => n35901, A3 => n35902, A4 => 
                           n35903, ZN => n35904);
   U522 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_17_port, B1 => 
                           n36256, B2 => REGISTERS_21_17_port, ZN => n35905);
   U523 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_17_port, B1 => 
                           n36252, B2 => REGISTERS_7_17_port, ZN => n35906);
   U524 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_17_port, B1 => 
                           n36249, B2 => REGISTERS_5_17_port, C1 => n36247, C2 
                           => REGISTERS_18_17_port, ZN => n35907);
   U525 : NAND3_X1 port map( A1 => n35905, A2 => n35906, A3 => n35907, ZN => 
                           n35908);
   U526 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_17_port, B1 => 
                           n36246, B2 => REGISTERS_19_17_port, ZN => n35909);
   U527 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_17_port, B1 => 
                           n36257, B2 => REGISTERS_23_17_port, ZN => n35910);
   U528 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_17_port, B1 => 
                           n36241, B2 => REGISTERS_10_17_port, ZN => n35911);
   U529 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_17_port, B1 => 
                           n36266, B2 => REGISTERS_27_17_port, ZN => n35912);
   U530 : NAND4_X1 port map( A1 => n35909, A2 => n35910, A3 => n35911, A4 => 
                           n35912, ZN => n35913);
   U531 : OR4_X1 port map( A1 => n35899, A2 => n35904, A3 => n35908, A4 => 
                           n35913, ZN => OUTB(17));
   U532 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_16_port, B1 => 
                           n36237, B2 => REGISTERS_14_16_port, ZN => n35914);
   U533 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_16_port, B1 => 
                           n36242, B2 => REGISTERS_4_16_port, ZN => n35915);
   U534 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_16_port, B1 => 
                           n36245, B2 => REGISTERS_22_16_port, ZN => n35916);
   U535 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_16_port, B1 => 
                           n36258, B2 => REGISTERS_9_16_port, ZN => n35917);
   U536 : NAND4_X1 port map( A1 => n35914, A2 => n35915, A3 => n35916, A4 => 
                           n35917, ZN => n35918);
   U537 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_16_port, B1 => 
                           n36263, B2 => REGISTERS_25_16_port, ZN => n35919);
   U538 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_16_port, B1 => 
                           n36264, B2 => REGISTERS_2_16_port, ZN => n35920);
   U539 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_16_port, B1 => 
                           n36261, B2 => REGISTERS_13_16_port, ZN => n35921);
   U540 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_16_port, B1 => 
                           n36259, B2 => REGISTERS_8_16_port, ZN => n35922);
   U541 : NAND4_X1 port map( A1 => n35919, A2 => n35920, A3 => n35921, A4 => 
                           n35922, ZN => n35923);
   U542 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_16_port, B1 => 
                           n36256, B2 => REGISTERS_21_16_port, ZN => n35924);
   U543 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_16_port, B1 => 
                           n36252, B2 => REGISTERS_7_16_port, ZN => n35925);
   U544 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_16_port, B1 => 
                           n36249, B2 => REGISTERS_5_16_port, C1 => n36247, C2 
                           => REGISTERS_18_16_port, ZN => n35926);
   U545 : NAND3_X1 port map( A1 => n35924, A2 => n35925, A3 => n35926, ZN => 
                           n35927);
   U546 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_16_port, B1 => 
                           n36246, B2 => REGISTERS_19_16_port, ZN => n35928);
   U547 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_16_port, B1 => 
                           n36257, B2 => REGISTERS_23_16_port, ZN => n35929);
   U548 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_16_port, B1 => 
                           n36241, B2 => REGISTERS_10_16_port, ZN => n35930);
   U549 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_16_port, B1 => 
                           n36266, B2 => REGISTERS_27_16_port, ZN => n35931);
   U550 : NAND4_X1 port map( A1 => n35928, A2 => n35929, A3 => n35930, A4 => 
                           n35931, ZN => n35932);
   U551 : OR4_X1 port map( A1 => n35918, A2 => n35923, A3 => n35927, A4 => 
                           n35932, ZN => OUTB(16));
   U552 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_15_port, B1 => 
                           n36237, B2 => REGISTERS_14_15_port, ZN => n35933);
   U553 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_15_port, B1 => 
                           n36242, B2 => REGISTERS_4_15_port, ZN => n35934);
   U554 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_15_port, B1 => 
                           n36245, B2 => REGISTERS_22_15_port, ZN => n35935);
   U555 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_15_port, B1 => 
                           n36258, B2 => REGISTERS_9_15_port, ZN => n35936);
   U556 : NAND4_X1 port map( A1 => n35933, A2 => n35934, A3 => n35935, A4 => 
                           n35936, ZN => n35937);
   U557 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_15_port, B1 => 
                           n36263, B2 => REGISTERS_25_15_port, ZN => n35938);
   U558 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_15_port, B1 => 
                           n36264, B2 => REGISTERS_2_15_port, ZN => n35939);
   U559 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_15_port, B1 => 
                           n36261, B2 => REGISTERS_13_15_port, ZN => n35940);
   U560 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_15_port, B1 => 
                           n36259, B2 => REGISTERS_8_15_port, ZN => n35941);
   U561 : NAND4_X1 port map( A1 => n35938, A2 => n35939, A3 => n35940, A4 => 
                           n35941, ZN => n35942);
   U562 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_15_port, B1 => 
                           n36256, B2 => REGISTERS_21_15_port, ZN => n35943);
   U563 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_15_port, B1 => 
                           n36252, B2 => REGISTERS_7_15_port, ZN => n35944);
   U564 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_15_port, B1 => 
                           n36249, B2 => REGISTERS_5_15_port, C1 => n36247, C2 
                           => REGISTERS_18_15_port, ZN => n35945);
   U565 : NAND3_X1 port map( A1 => n35943, A2 => n35944, A3 => n35945, ZN => 
                           n35946);
   U566 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_15_port, B1 => 
                           n36246, B2 => REGISTERS_19_15_port, ZN => n35947);
   U567 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_15_port, B1 => 
                           n36257, B2 => REGISTERS_23_15_port, ZN => n35948);
   U568 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_15_port, B1 => 
                           n36241, B2 => REGISTERS_10_15_port, ZN => n35949);
   U569 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_15_port, B1 => 
                           n36266, B2 => REGISTERS_27_15_port, ZN => n35950);
   U570 : NAND4_X1 port map( A1 => n35947, A2 => n35948, A3 => n35949, A4 => 
                           n35950, ZN => n35951);
   U571 : OR4_X1 port map( A1 => n35937, A2 => n35942, A3 => n35946, A4 => 
                           n35951, ZN => OUTB(15));
   U572 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_14_port, B1 => 
                           n36237, B2 => REGISTERS_14_14_port, ZN => n35952);
   U573 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_14_port, B1 => 
                           n36242, B2 => REGISTERS_4_14_port, ZN => n35953);
   U574 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_14_port, B1 => 
                           n36245, B2 => REGISTERS_22_14_port, ZN => n35954);
   U575 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_14_port, B1 => 
                           n36258, B2 => REGISTERS_9_14_port, ZN => n35955);
   U576 : NAND4_X1 port map( A1 => n35952, A2 => n35953, A3 => n35954, A4 => 
                           n35955, ZN => n35956);
   U577 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_14_port, B1 => 
                           n36263, B2 => REGISTERS_25_14_port, ZN => n35957);
   U578 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_14_port, B1 => 
                           n36264, B2 => REGISTERS_2_14_port, ZN => n35958);
   U579 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_14_port, B1 => 
                           n36261, B2 => REGISTERS_13_14_port, ZN => n35959);
   U580 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_14_port, B1 => 
                           n36259, B2 => REGISTERS_8_14_port, ZN => n35960);
   U581 : NAND4_X1 port map( A1 => n35957, A2 => n35958, A3 => n35959, A4 => 
                           n35960, ZN => n35961);
   U582 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_14_port, B1 => 
                           n36256, B2 => REGISTERS_21_14_port, ZN => n35962);
   U583 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_14_port, B1 => 
                           n36252, B2 => REGISTERS_7_14_port, ZN => n35963);
   U584 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_14_port, B1 => 
                           n36249, B2 => REGISTERS_5_14_port, C1 => n36247, C2 
                           => REGISTERS_18_14_port, ZN => n35964);
   U585 : NAND3_X1 port map( A1 => n35962, A2 => n35963, A3 => n35964, ZN => 
                           n35965);
   U586 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_14_port, B1 => 
                           n36246, B2 => REGISTERS_19_14_port, ZN => n35966);
   U587 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_14_port, B1 => 
                           n36257, B2 => REGISTERS_23_14_port, ZN => n35967);
   U588 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_14_port, B1 => 
                           n36241, B2 => REGISTERS_10_14_port, ZN => n35968);
   U589 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_14_port, B1 => 
                           n36266, B2 => REGISTERS_27_14_port, ZN => n35969);
   U590 : NAND4_X1 port map( A1 => n35966, A2 => n35967, A3 => n35968, A4 => 
                           n35969, ZN => n35970);
   U591 : OR4_X1 port map( A1 => n35956, A2 => n35961, A3 => n35965, A4 => 
                           n35970, ZN => OUTB(14));
   U592 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_13_port, B1 => 
                           n36237, B2 => REGISTERS_14_13_port, ZN => n35971);
   U593 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_13_port, B1 => 
                           n36242, B2 => REGISTERS_4_13_port, ZN => n35972);
   U594 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_13_port, B1 => 
                           n36245, B2 => REGISTERS_22_13_port, ZN => n35973);
   U595 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_13_port, B1 => 
                           n36258, B2 => REGISTERS_9_13_port, ZN => n35974);
   U596 : NAND4_X1 port map( A1 => n35971, A2 => n35972, A3 => n35973, A4 => 
                           n35974, ZN => n35975);
   U597 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_13_port, B1 => 
                           n36263, B2 => REGISTERS_25_13_port, ZN => n35976);
   U598 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_13_port, B1 => 
                           n36264, B2 => REGISTERS_2_13_port, ZN => n35977);
   U599 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_13_port, B1 => 
                           n36261, B2 => REGISTERS_13_13_port, ZN => n35978);
   U600 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_13_port, B1 => 
                           n36259, B2 => REGISTERS_8_13_port, ZN => n35979);
   U601 : NAND4_X1 port map( A1 => n35976, A2 => n35977, A3 => n35978, A4 => 
                           n35979, ZN => n35980);
   U602 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_13_port, B1 => 
                           n36256, B2 => REGISTERS_21_13_port, ZN => n35981);
   U603 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_13_port, B1 => 
                           n36252, B2 => REGISTERS_7_13_port, ZN => n35982);
   U604 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_13_port, B1 => 
                           n36249, B2 => REGISTERS_5_13_port, C1 => n36247, C2 
                           => REGISTERS_18_13_port, ZN => n35983);
   U605 : NAND3_X1 port map( A1 => n35981, A2 => n35982, A3 => n35983, ZN => 
                           n35984);
   U606 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_13_port, B1 => 
                           n36246, B2 => REGISTERS_19_13_port, ZN => n35985);
   U607 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_13_port, B1 => 
                           n36257, B2 => REGISTERS_23_13_port, ZN => n35986);
   U608 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_13_port, B1 => 
                           n36241, B2 => REGISTERS_10_13_port, ZN => n35987);
   U609 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_13_port, B1 => 
                           n36266, B2 => REGISTERS_27_13_port, ZN => n35988);
   U610 : NAND4_X1 port map( A1 => n35985, A2 => n35986, A3 => n35987, A4 => 
                           n35988, ZN => n35989);
   U611 : OR4_X1 port map( A1 => n35975, A2 => n35980, A3 => n35984, A4 => 
                           n35989, ZN => OUTB(13));
   U612 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_12_port, B1 => 
                           n36237, B2 => REGISTERS_14_12_port, ZN => n35990);
   U613 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_12_port, B1 => 
                           n36242, B2 => REGISTERS_4_12_port, ZN => n35991);
   U614 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_12_port, B1 => 
                           n36245, B2 => REGISTERS_22_12_port, ZN => n35992);
   U615 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_12_port, B1 => 
                           n36258, B2 => REGISTERS_9_12_port, ZN => n35993);
   U616 : NAND4_X1 port map( A1 => n35990, A2 => n35991, A3 => n35992, A4 => 
                           n35993, ZN => n35994);
   U617 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_12_port, B1 => 
                           n36263, B2 => REGISTERS_25_12_port, ZN => n35995);
   U618 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_12_port, B1 => 
                           n36264, B2 => REGISTERS_2_12_port, ZN => n35996);
   U619 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_12_port, B1 => 
                           n36261, B2 => REGISTERS_13_12_port, ZN => n35997);
   U620 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_12_port, B1 => 
                           n36259, B2 => REGISTERS_8_12_port, ZN => n35998);
   U621 : NAND4_X1 port map( A1 => n35995, A2 => n35996, A3 => n35997, A4 => 
                           n35998, ZN => n35999);
   U622 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_12_port, B1 => 
                           n36256, B2 => REGISTERS_21_12_port, ZN => n36000);
   U623 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_12_port, B1 => 
                           n36252, B2 => REGISTERS_7_12_port, ZN => n36001);
   U624 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_12_port, B1 => 
                           n36249, B2 => REGISTERS_5_12_port, C1 => n36247, C2 
                           => REGISTERS_18_12_port, ZN => n36002);
   U625 : NAND3_X1 port map( A1 => n36000, A2 => n36001, A3 => n36002, ZN => 
                           n36003);
   U626 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_12_port, B1 => 
                           n36246, B2 => REGISTERS_19_12_port, ZN => n36004);
   U627 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_12_port, B1 => 
                           n36257, B2 => REGISTERS_23_12_port, ZN => n36005);
   U628 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_12_port, B1 => 
                           n36241, B2 => REGISTERS_10_12_port, ZN => n36006);
   U629 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_12_port, B1 => 
                           n36266, B2 => REGISTERS_27_12_port, ZN => n36007);
   U630 : NAND4_X1 port map( A1 => n36004, A2 => n36005, A3 => n36006, A4 => 
                           n36007, ZN => n36008);
   U631 : OR4_X1 port map( A1 => n35994, A2 => n35999, A3 => n36003, A4 => 
                           n36008, ZN => OUTB(12));
   U632 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_11_port, B1 => 
                           n36237, B2 => REGISTERS_14_11_port, ZN => n36009);
   U633 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_11_port, B1 => 
                           n36242, B2 => REGISTERS_4_11_port, ZN => n36010);
   U634 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_11_port, B1 => 
                           n36245, B2 => REGISTERS_22_11_port, ZN => n36011);
   U635 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_11_port, B1 => 
                           n36258, B2 => REGISTERS_9_11_port, ZN => n36012);
   U636 : NAND4_X1 port map( A1 => n36009, A2 => n36010, A3 => n36011, A4 => 
                           n36012, ZN => n36013);
   U637 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_11_port, B1 => 
                           n36263, B2 => REGISTERS_25_11_port, ZN => n36014);
   U638 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_11_port, B1 => 
                           n36264, B2 => REGISTERS_2_11_port, ZN => n36015);
   U639 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_11_port, B1 => 
                           n36261, B2 => REGISTERS_13_11_port, ZN => n36016);
   U640 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_11_port, B1 => 
                           n36259, B2 => REGISTERS_8_11_port, ZN => n36017);
   U641 : NAND4_X1 port map( A1 => n36014, A2 => n36015, A3 => n36016, A4 => 
                           n36017, ZN => n36018);
   U642 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_11_port, B1 => 
                           n36256, B2 => REGISTERS_21_11_port, ZN => n36019);
   U643 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_11_port, B1 => 
                           n36252, B2 => REGISTERS_7_11_port, ZN => n36020);
   U644 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_11_port, B1 => 
                           n36249, B2 => REGISTERS_5_11_port, C1 => n36247, C2 
                           => REGISTERS_18_11_port, ZN => n36021);
   U645 : NAND3_X1 port map( A1 => n36019, A2 => n36020, A3 => n36021, ZN => 
                           n36022);
   U646 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_11_port, B1 => 
                           n36246, B2 => REGISTERS_19_11_port, ZN => n36023);
   U647 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_11_port, B1 => 
                           n36257, B2 => REGISTERS_23_11_port, ZN => n36024);
   U648 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_11_port, B1 => 
                           n36241, B2 => REGISTERS_10_11_port, ZN => n36025);
   U649 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_11_port, B1 => 
                           n36266, B2 => REGISTERS_27_11_port, ZN => n36026);
   U650 : NAND4_X1 port map( A1 => n36023, A2 => n36024, A3 => n36025, A4 => 
                           n36026, ZN => n36027);
   U651 : OR4_X1 port map( A1 => n36013, A2 => n36018, A3 => n36022, A4 => 
                           n36027, ZN => OUTB(11));
   U652 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_10_port, B1 => 
                           n36237, B2 => REGISTERS_14_10_port, ZN => n36028);
   U653 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_10_port, B1 => 
                           n36242, B2 => REGISTERS_4_10_port, ZN => n36029);
   U654 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_10_port, B1 => 
                           n36245, B2 => REGISTERS_22_10_port, ZN => n36030);
   U655 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_10_port, B1 => 
                           n36258, B2 => REGISTERS_9_10_port, ZN => n36031);
   U656 : NAND4_X1 port map( A1 => n36028, A2 => n36029, A3 => n36030, A4 => 
                           n36031, ZN => n36032);
   U657 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_10_port, B1 => 
                           n36263, B2 => REGISTERS_25_10_port, ZN => n36033);
   U658 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_10_port, B1 => 
                           n36264, B2 => REGISTERS_2_10_port, ZN => n36034);
   U659 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_10_port, B1 => 
                           n36261, B2 => REGISTERS_13_10_port, ZN => n36035);
   U660 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_10_port, B1 => 
                           n36259, B2 => REGISTERS_8_10_port, ZN => n36036);
   U661 : NAND4_X1 port map( A1 => n36033, A2 => n36034, A3 => n36035, A4 => 
                           n36036, ZN => n36037);
   U662 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_10_port, B1 => 
                           n36256, B2 => REGISTERS_21_10_port, ZN => n36038);
   U663 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_10_port, B1 => 
                           n36252, B2 => REGISTERS_7_10_port, ZN => n36039);
   U664 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_10_port, B1 => 
                           n36249, B2 => REGISTERS_5_10_port, C1 => n36247, C2 
                           => REGISTERS_18_10_port, ZN => n36040);
   U665 : NAND3_X1 port map( A1 => n36038, A2 => n36039, A3 => n36040, ZN => 
                           n36041);
   U666 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_10_port, B1 => 
                           n36246, B2 => REGISTERS_19_10_port, ZN => n36042);
   U667 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_10_port, B1 => 
                           n36257, B2 => REGISTERS_23_10_port, ZN => n36043);
   U668 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_10_port, B1 => 
                           n36241, B2 => REGISTERS_10_10_port, ZN => n36044);
   U669 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_10_port, B1 => 
                           n36266, B2 => REGISTERS_27_10_port, ZN => n36045);
   U670 : NAND4_X1 port map( A1 => n36042, A2 => n36043, A3 => n36044, A4 => 
                           n36045, ZN => n36046);
   U671 : OR4_X1 port map( A1 => n36032, A2 => n36037, A3 => n36041, A4 => 
                           n36046, ZN => OUTB(10));
   U672 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_9_port, B1 => 
                           n36237, B2 => REGISTERS_14_9_port, ZN => n36047);
   U673 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_9_port, B1 => 
                           n36242, B2 => REGISTERS_4_9_port, ZN => n36048);
   U674 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_9_port, B1 => 
                           n36245, B2 => REGISTERS_22_9_port, ZN => n36049);
   U675 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_9_port, B1 => 
                           n36258, B2 => REGISTERS_9_9_port, ZN => n36050);
   U676 : NAND4_X1 port map( A1 => n36047, A2 => n36048, A3 => n36049, A4 => 
                           n36050, ZN => n36051);
   U677 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_9_port, B1 => 
                           n36263, B2 => REGISTERS_25_9_port, ZN => n36052);
   U678 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_9_port, B1 => 
                           n36264, B2 => REGISTERS_2_9_port, ZN => n36053);
   U679 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_9_port, B1 => 
                           n36261, B2 => REGISTERS_13_9_port, ZN => n36054);
   U680 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_9_port, B1 => 
                           n36259, B2 => REGISTERS_8_9_port, ZN => n36055);
   U681 : NAND4_X1 port map( A1 => n36052, A2 => n36053, A3 => n36054, A4 => 
                           n36055, ZN => n36056);
   U682 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_9_port, B1 => 
                           n36256, B2 => REGISTERS_21_9_port, ZN => n36057);
   U683 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_9_port, B1 => 
                           n36252, B2 => REGISTERS_7_9_port, ZN => n36058);
   U684 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_9_port, B1 => 
                           n36249, B2 => REGISTERS_5_9_port, C1 => n36247, C2 
                           => REGISTERS_18_9_port, ZN => n36059);
   U685 : NAND3_X1 port map( A1 => n36057, A2 => n36058, A3 => n36059, ZN => 
                           n36060);
   U686 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_9_port, B1 => 
                           n36246, B2 => REGISTERS_19_9_port, ZN => n36061);
   U687 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_9_port, B1 => 
                           n36257, B2 => REGISTERS_23_9_port, ZN => n36062);
   U688 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_9_port, B1 => 
                           n36241, B2 => REGISTERS_10_9_port, ZN => n36063);
   U689 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_9_port, B1 => 
                           n36266, B2 => REGISTERS_27_9_port, ZN => n36064);
   U690 : NAND4_X1 port map( A1 => n36061, A2 => n36062, A3 => n36063, A4 => 
                           n36064, ZN => n36065);
   U691 : OR4_X1 port map( A1 => n36051, A2 => n36056, A3 => n36060, A4 => 
                           n36065, ZN => OUTB(9));
   U692 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_8_port, B1 => 
                           n36237, B2 => REGISTERS_14_8_port, ZN => n36066);
   U693 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_8_port, B1 => 
                           n36242, B2 => REGISTERS_4_8_port, ZN => n36067);
   U694 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_8_port, B1 => 
                           n36245, B2 => REGISTERS_22_8_port, ZN => n36068);
   U695 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_8_port, B1 => 
                           n36258, B2 => REGISTERS_9_8_port, ZN => n36069);
   U696 : NAND4_X1 port map( A1 => n36066, A2 => n36067, A3 => n36068, A4 => 
                           n36069, ZN => n36070);
   U697 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_8_port, B1 => 
                           n36263, B2 => REGISTERS_25_8_port, ZN => n36071);
   U698 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_8_port, B1 => 
                           n36264, B2 => REGISTERS_2_8_port, ZN => n36072);
   U699 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_8_port, B1 => 
                           n36261, B2 => REGISTERS_13_8_port, ZN => n36073);
   U700 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_8_port, B1 => 
                           n36259, B2 => REGISTERS_8_8_port, ZN => n36074);
   U701 : NAND4_X1 port map( A1 => n36071, A2 => n36072, A3 => n36073, A4 => 
                           n36074, ZN => n36075);
   U702 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_8_port, B1 => 
                           n36256, B2 => REGISTERS_21_8_port, ZN => n36076);
   U703 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_8_port, B1 => 
                           n36252, B2 => REGISTERS_7_8_port, ZN => n36077);
   U704 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_8_port, B1 => 
                           n36249, B2 => REGISTERS_5_8_port, C1 => n36247, C2 
                           => REGISTERS_18_8_port, ZN => n36078);
   U705 : NAND3_X1 port map( A1 => n36076, A2 => n36077, A3 => n36078, ZN => 
                           n36079);
   U706 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_8_port, B1 => 
                           n36246, B2 => REGISTERS_19_8_port, ZN => n36080);
   U707 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_8_port, B1 => 
                           n36257, B2 => REGISTERS_23_8_port, ZN => n36081);
   U708 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_8_port, B1 => 
                           n36241, B2 => REGISTERS_10_8_port, ZN => n36082);
   U709 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_8_port, B1 => 
                           n36266, B2 => REGISTERS_27_8_port, ZN => n36083);
   U710 : NAND4_X1 port map( A1 => n36080, A2 => n36081, A3 => n36082, A4 => 
                           n36083, ZN => n36084);
   U711 : OR4_X1 port map( A1 => n36070, A2 => n36075, A3 => n36079, A4 => 
                           n36084, ZN => OUTB(8));
   U712 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_7_port, B1 => 
                           n36237, B2 => REGISTERS_14_7_port, ZN => n36085);
   U713 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_7_port, B1 => 
                           n36242, B2 => REGISTERS_4_7_port, ZN => n36086);
   U714 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_7_port, B1 => 
                           n36245, B2 => REGISTERS_22_7_port, ZN => n36087);
   U715 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_7_port, B1 => 
                           n36258, B2 => REGISTERS_9_7_port, ZN => n36088);
   U716 : NAND4_X1 port map( A1 => n36085, A2 => n36086, A3 => n36087, A4 => 
                           n36088, ZN => n36089);
   U717 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_7_port, B1 => 
                           n36263, B2 => REGISTERS_25_7_port, ZN => n36090);
   U718 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_7_port, B1 => 
                           n36264, B2 => REGISTERS_2_7_port, ZN => n36091);
   U719 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_7_port, B1 => 
                           n36261, B2 => REGISTERS_13_7_port, ZN => n36092);
   U720 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_7_port, B1 => 
                           n36259, B2 => REGISTERS_8_7_port, ZN => n36093);
   U721 : NAND4_X1 port map( A1 => n36090, A2 => n36091, A3 => n36092, A4 => 
                           n36093, ZN => n36094);
   U722 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_7_port, B1 => 
                           n36256, B2 => REGISTERS_21_7_port, ZN => n36095);
   U723 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_7_port, B1 => 
                           n36252, B2 => REGISTERS_7_7_port, ZN => n36096);
   U724 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_7_port, B1 => 
                           n36249, B2 => REGISTERS_5_7_port, C1 => n36247, C2 
                           => REGISTERS_18_7_port, ZN => n36097);
   U725 : NAND3_X1 port map( A1 => n36095, A2 => n36096, A3 => n36097, ZN => 
                           n36098);
   U726 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_7_port, B1 => 
                           n36246, B2 => REGISTERS_19_7_port, ZN => n36099);
   U727 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_7_port, B1 => 
                           n36257, B2 => REGISTERS_23_7_port, ZN => n36100);
   U728 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_7_port, B1 => 
                           n36241, B2 => REGISTERS_10_7_port, ZN => n36101);
   U729 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_7_port, B1 => 
                           n36266, B2 => REGISTERS_27_7_port, ZN => n36102);
   U730 : NAND4_X1 port map( A1 => n36099, A2 => n36100, A3 => n36101, A4 => 
                           n36102, ZN => n36103);
   U731 : OR4_X1 port map( A1 => n36089, A2 => n36094, A3 => n36098, A4 => 
                           n36103, ZN => OUTB(7));
   U732 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_6_port, B1 => 
                           n36237, B2 => REGISTERS_14_6_port, ZN => n36104);
   U733 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_6_port, B1 => 
                           n36242, B2 => REGISTERS_4_6_port, ZN => n36105);
   U734 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_6_port, B1 => 
                           n36245, B2 => REGISTERS_22_6_port, ZN => n36106);
   U735 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_6_port, B1 => 
                           n36258, B2 => REGISTERS_9_6_port, ZN => n36107);
   U736 : NAND4_X1 port map( A1 => n36104, A2 => n36105, A3 => n36106, A4 => 
                           n36107, ZN => n36108);
   U737 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_6_port, B1 => 
                           n36263, B2 => REGISTERS_25_6_port, ZN => n36109);
   U738 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_6_port, B1 => 
                           n36264, B2 => REGISTERS_2_6_port, ZN => n36110);
   U739 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_6_port, B1 => 
                           n36261, B2 => REGISTERS_13_6_port, ZN => n36111);
   U740 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_6_port, B1 => 
                           n36259, B2 => REGISTERS_8_6_port, ZN => n36112);
   U741 : NAND4_X1 port map( A1 => n36109, A2 => n36110, A3 => n36111, A4 => 
                           n36112, ZN => n36113);
   U742 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_6_port, B1 => 
                           n36256, B2 => REGISTERS_21_6_port, ZN => n36114);
   U743 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_6_port, B1 => 
                           n36252, B2 => REGISTERS_7_6_port, ZN => n36115);
   U744 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_6_port, B1 => 
                           n36249, B2 => REGISTERS_5_6_port, C1 => n36247, C2 
                           => REGISTERS_18_6_port, ZN => n36116);
   U745 : NAND3_X1 port map( A1 => n36114, A2 => n36115, A3 => n36116, ZN => 
                           n36117);
   U746 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_6_port, B1 => 
                           n36246, B2 => REGISTERS_19_6_port, ZN => n36118);
   U747 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_6_port, B1 => 
                           n36257, B2 => REGISTERS_23_6_port, ZN => n36119);
   U748 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_6_port, B1 => 
                           n36241, B2 => REGISTERS_10_6_port, ZN => n36120);
   U749 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_6_port, B1 => 
                           n36266, B2 => REGISTERS_27_6_port, ZN => n36121);
   U750 : NAND4_X1 port map( A1 => n36118, A2 => n36119, A3 => n36120, A4 => 
                           n36121, ZN => n36122);
   U751 : OR4_X1 port map( A1 => n36108, A2 => n36113, A3 => n36117, A4 => 
                           n36122, ZN => OUTB(6));
   U752 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_5_port, B1 => 
                           n36237, B2 => REGISTERS_14_5_port, ZN => n36123);
   U753 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_5_port, B1 => 
                           n36242, B2 => REGISTERS_4_5_port, ZN => n36124);
   U754 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_5_port, B1 => 
                           n36245, B2 => REGISTERS_22_5_port, ZN => n36125);
   U755 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_5_port, B1 => 
                           n36258, B2 => REGISTERS_9_5_port, ZN => n36126);
   U756 : NAND4_X1 port map( A1 => n36123, A2 => n36124, A3 => n36125, A4 => 
                           n36126, ZN => n36127);
   U757 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_5_port, B1 => 
                           n36263, B2 => REGISTERS_25_5_port, ZN => n36128);
   U758 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_5_port, B1 => 
                           n36264, B2 => REGISTERS_2_5_port, ZN => n36129);
   U759 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_5_port, B1 => 
                           n36261, B2 => REGISTERS_13_5_port, ZN => n36130);
   U760 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_5_port, B1 => 
                           n36259, B2 => REGISTERS_8_5_port, ZN => n36131);
   U761 : NAND4_X1 port map( A1 => n36128, A2 => n36129, A3 => n36130, A4 => 
                           n36131, ZN => n36132);
   U762 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_5_port, B1 => 
                           n36256, B2 => REGISTERS_21_5_port, ZN => n36133);
   U763 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_5_port, B1 => 
                           n36252, B2 => REGISTERS_7_5_port, ZN => n36134);
   U764 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_5_port, B1 => 
                           n36249, B2 => REGISTERS_5_5_port, C1 => n36247, C2 
                           => REGISTERS_18_5_port, ZN => n36135);
   U765 : NAND3_X1 port map( A1 => n36133, A2 => n36134, A3 => n36135, ZN => 
                           n36136);
   U766 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_5_port, B1 => 
                           n36246, B2 => REGISTERS_19_5_port, ZN => n36137);
   U767 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_5_port, B1 => 
                           n36257, B2 => REGISTERS_23_5_port, ZN => n36138);
   U768 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_5_port, B1 => 
                           n36241, B2 => REGISTERS_10_5_port, ZN => n36139);
   U769 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_5_port, B1 => 
                           n36266, B2 => REGISTERS_27_5_port, ZN => n36140);
   U770 : NAND4_X1 port map( A1 => n36137, A2 => n36138, A3 => n36139, A4 => 
                           n36140, ZN => n36141);
   U771 : OR4_X1 port map( A1 => n36127, A2 => n36132, A3 => n36136, A4 => 
                           n36141, ZN => OUTB(5));
   U772 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_4_port, B1 => 
                           n36237, B2 => REGISTERS_14_4_port, ZN => n36142);
   U773 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_4_port, B1 => 
                           n36242, B2 => REGISTERS_4_4_port, ZN => n36143);
   U774 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_4_port, B1 => 
                           n36245, B2 => REGISTERS_22_4_port, ZN => n36144);
   U775 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_4_port, B1 => 
                           n36258, B2 => REGISTERS_9_4_port, ZN => n36145);
   U776 : NAND4_X1 port map( A1 => n36142, A2 => n36143, A3 => n36144, A4 => 
                           n36145, ZN => n36146);
   U777 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_4_port, B1 => 
                           n36263, B2 => REGISTERS_25_4_port, ZN => n36147);
   U778 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_4_port, B1 => 
                           n36264, B2 => REGISTERS_2_4_port, ZN => n36148);
   U779 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_4_port, B1 => 
                           n36261, B2 => REGISTERS_13_4_port, ZN => n36149);
   U780 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_4_port, B1 => 
                           n36259, B2 => REGISTERS_8_4_port, ZN => n36150);
   U781 : NAND4_X1 port map( A1 => n36147, A2 => n36148, A3 => n36149, A4 => 
                           n36150, ZN => n36151);
   U782 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_4_port, B1 => 
                           n36256, B2 => REGISTERS_21_4_port, ZN => n36152);
   U783 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_4_port, B1 => 
                           n36252, B2 => REGISTERS_7_4_port, ZN => n36153);
   U784 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_4_port, B1 => 
                           n36249, B2 => REGISTERS_5_4_port, C1 => n36247, C2 
                           => REGISTERS_18_4_port, ZN => n36154);
   U785 : NAND3_X1 port map( A1 => n36152, A2 => n36153, A3 => n36154, ZN => 
                           n36155);
   U786 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_4_port, B1 => 
                           n36246, B2 => REGISTERS_19_4_port, ZN => n36156);
   U787 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_4_port, B1 => 
                           n36257, B2 => REGISTERS_23_4_port, ZN => n36157);
   U788 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_4_port, B1 => 
                           n36241, B2 => REGISTERS_10_4_port, ZN => n36158);
   U789 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_4_port, B1 => 
                           n36266, B2 => REGISTERS_27_4_port, ZN => n36159);
   U790 : NAND4_X1 port map( A1 => n36156, A2 => n36157, A3 => n36158, A4 => 
                           n36159, ZN => n36160);
   U791 : OR4_X1 port map( A1 => n36146, A2 => n36151, A3 => n36155, A4 => 
                           n36160, ZN => OUTB(4));
   U792 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_3_port, B1 => 
                           n36237, B2 => REGISTERS_14_3_port, ZN => n36161);
   U793 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_3_port, B1 => 
                           n36242, B2 => REGISTERS_4_3_port, ZN => n36162);
   U794 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_3_port, B1 => 
                           n36245, B2 => REGISTERS_22_3_port, ZN => n36163);
   U795 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_3_port, B1 => 
                           n36258, B2 => REGISTERS_9_3_port, ZN => n36164);
   U796 : NAND4_X1 port map( A1 => n36161, A2 => n36162, A3 => n36163, A4 => 
                           n36164, ZN => n36165);
   U797 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_3_port, B1 => 
                           n36263, B2 => REGISTERS_25_3_port, ZN => n36166);
   U798 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_3_port, B1 => 
                           n36264, B2 => REGISTERS_2_3_port, ZN => n36167);
   U799 : AOI22_X1 port map( A1 => n36855, A2 => REGISTERS_31_3_port, B1 => 
                           n36261, B2 => REGISTERS_13_3_port, ZN => n36168);
   U800 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_3_port, B1 => 
                           n36259, B2 => REGISTERS_8_3_port, ZN => n36169);
   U801 : NAND4_X1 port map( A1 => n36166, A2 => n36167, A3 => n36168, A4 => 
                           n36169, ZN => n36170);
   U802 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_3_port, B1 => 
                           n36256, B2 => REGISTERS_21_3_port, ZN => n36171);
   U803 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_3_port, B1 => 
                           n36252, B2 => REGISTERS_7_3_port, ZN => n36172);
   U804 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_3_port, B1 => 
                           n36249, B2 => REGISTERS_5_3_port, C1 => n36247, C2 
                           => REGISTERS_18_3_port, ZN => n36173);
   U805 : NAND3_X1 port map( A1 => n36171, A2 => n36172, A3 => n36173, ZN => 
                           n36174);
   U806 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_3_port, B1 => 
                           n36246, B2 => REGISTERS_19_3_port, ZN => n36175);
   U807 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_3_port, B1 => 
                           n36257, B2 => REGISTERS_23_3_port, ZN => n36176);
   U808 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_3_port, B1 => 
                           n36241, B2 => REGISTERS_10_3_port, ZN => n36177);
   U809 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_3_port, B1 => 
                           n36266, B2 => REGISTERS_27_3_port, ZN => n36178);
   U810 : NAND4_X1 port map( A1 => n36175, A2 => n36176, A3 => n36177, A4 => 
                           n36178, ZN => n36179);
   U811 : OR4_X1 port map( A1 => n36165, A2 => n36170, A3 => n36174, A4 => 
                           n36179, ZN => OUTB(3));
   U812 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_2_port, B1 => 
                           n36237, B2 => REGISTERS_14_2_port, ZN => n36180);
   U813 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_2_port, B1 => 
                           n36242, B2 => REGISTERS_4_2_port, ZN => n36181);
   U814 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_2_port, B1 => 
                           n36245, B2 => REGISTERS_22_2_port, ZN => n36182);
   U815 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_2_port, B1 => 
                           n36258, B2 => REGISTERS_9_2_port, ZN => n36183);
   U816 : NAND4_X1 port map( A1 => n36180, A2 => n36181, A3 => n36182, A4 => 
                           n36183, ZN => n36184);
   U817 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_2_port, B1 => 
                           n36263, B2 => REGISTERS_25_2_port, ZN => n36185);
   U818 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_2_port, B1 => 
                           n36264, B2 => REGISTERS_2_2_port, ZN => n36186);
   U819 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_2_port, B1 => 
                           n36261, B2 => REGISTERS_13_2_port, ZN => n36187);
   U820 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_2_port, B1 => 
                           n36259, B2 => REGISTERS_8_2_port, ZN => n36188);
   U821 : NAND4_X1 port map( A1 => n36185, A2 => n36186, A3 => n36187, A4 => 
                           n36188, ZN => n36189);
   U822 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_2_port, B1 => 
                           n36256, B2 => REGISTERS_21_2_port, ZN => n36190);
   U823 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_2_port, B1 => 
                           n36252, B2 => REGISTERS_7_2_port, ZN => n36191);
   U824 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_2_port, B1 => 
                           n36249, B2 => REGISTERS_5_2_port, C1 => n36247, C2 
                           => REGISTERS_18_2_port, ZN => n36192);
   U825 : NAND3_X1 port map( A1 => n36190, A2 => n36191, A3 => n36192, ZN => 
                           n36193);
   U826 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_2_port, B1 => 
                           n36246, B2 => REGISTERS_19_2_port, ZN => n36194);
   U827 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_2_port, B1 => 
                           n36257, B2 => REGISTERS_23_2_port, ZN => n36195);
   U828 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_2_port, B1 => 
                           n36241, B2 => REGISTERS_10_2_port, ZN => n36196);
   U829 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_2_port, B1 => 
                           n36266, B2 => REGISTERS_27_2_port, ZN => n36197);
   U830 : NAND4_X1 port map( A1 => n36194, A2 => n36195, A3 => n36196, A4 => 
                           n36197, ZN => n36198);
   U831 : OR4_X1 port map( A1 => n36184, A2 => n36189, A3 => n36193, A4 => 
                           n36198, ZN => OUTB(2));
   U832 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_1_port, B1 => 
                           n36237, B2 => REGISTERS_14_1_port, ZN => n36199);
   U833 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_1_port, B1 => 
                           n36242, B2 => REGISTERS_4_1_port, ZN => n36200);
   U834 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_1_port, B1 => 
                           n36245, B2 => REGISTERS_22_1_port, ZN => n36201);
   U835 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_1_port, B1 => 
                           n36258, B2 => REGISTERS_9_1_port, ZN => n36202);
   U836 : NAND4_X1 port map( A1 => n36199, A2 => n36200, A3 => n36201, A4 => 
                           n36202, ZN => n36203);
   U837 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_1_port, B1 => 
                           n36263, B2 => REGISTERS_25_1_port, ZN => n36204);
   U838 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_1_port, B1 => 
                           n36264, B2 => REGISTERS_2_1_port, ZN => n36205);
   U839 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_1_port, B1 => 
                           n36261, B2 => REGISTERS_13_1_port, ZN => n36206);
   U840 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_1_port, B1 => 
                           n36259, B2 => REGISTERS_8_1_port, ZN => n36207);
   U841 : NAND4_X1 port map( A1 => n36204, A2 => n36205, A3 => n36206, A4 => 
                           n36207, ZN => n36208);
   U842 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_1_port, B1 => 
                           n36256, B2 => REGISTERS_21_1_port, ZN => n36209);
   U843 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_1_port, B1 => 
                           n36252, B2 => REGISTERS_7_1_port, ZN => n36210);
   U844 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_1_port, B1 => 
                           n36249, B2 => REGISTERS_5_1_port, C1 => n36247, C2 
                           => REGISTERS_18_1_port, ZN => n36211);
   U845 : NAND3_X1 port map( A1 => n36209, A2 => n36210, A3 => n36211, ZN => 
                           n36212);
   U846 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_1_port, B1 => 
                           n36246, B2 => REGISTERS_19_1_port, ZN => n36213);
   U847 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_1_port, B1 => 
                           n36257, B2 => REGISTERS_23_1_port, ZN => n36214);
   U848 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_1_port, B1 => 
                           n36241, B2 => REGISTERS_10_1_port, ZN => n36215);
   U849 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_1_port, B1 => 
                           n36266, B2 => REGISTERS_27_1_port, ZN => n36216);
   U850 : NAND4_X1 port map( A1 => n36213, A2 => n36214, A3 => n36215, A4 => 
                           n36216, ZN => n36217);
   U851 : OR4_X1 port map( A1 => n36203, A2 => n36208, A3 => n36212, A4 => 
                           n36217, ZN => OUTB(1));
   U852 : AOI22_X1 port map( A1 => n36240, A2 => REGISTERS_30_0_port, B1 => 
                           n36237, B2 => REGISTERS_14_0_port, ZN => n36218);
   U853 : AOI22_X1 port map( A1 => n36238, A2 => REGISTERS_3_0_port, B1 => 
                           n36242, B2 => REGISTERS_4_0_port, ZN => n36219);
   U854 : AOI22_X1 port map( A1 => n36250, A2 => REGISTERS_17_0_port, B1 => 
                           n36245, B2 => REGISTERS_22_0_port, ZN => n36220);
   U855 : AOI22_X1 port map( A1 => n36260, A2 => REGISTERS_15_0_port, B1 => 
                           n36258, B2 => REGISTERS_9_0_port, ZN => n36221);
   U856 : NAND4_X1 port map( A1 => n36218, A2 => n36219, A3 => n36220, A4 => 
                           n36221, ZN => n36222);
   U857 : AOI22_X1 port map( A1 => n36262, A2 => REGISTERS_16_0_port, B1 => 
                           n36263, B2 => REGISTERS_25_0_port, ZN => n36223);
   U858 : AOI22_X1 port map( A1 => n36265, A2 => REGISTERS_11_0_port, B1 => 
                           n36264, B2 => REGISTERS_2_0_port, ZN => n36224);
   U859 : AOI22_X1 port map( A1 => n36267, A2 => REGISTERS_31_0_port, B1 => 
                           n36261, B2 => REGISTERS_13_0_port, ZN => n36225);
   U860 : AOI22_X1 port map( A1 => n36255, A2 => REGISTERS_29_0_port, B1 => 
                           n36259, B2 => REGISTERS_8_0_port, ZN => n36226);
   U861 : NAND4_X1 port map( A1 => n36223, A2 => n36224, A3 => n36225, A4 => 
                           n36226, ZN => n36227);
   U862 : AOI22_X1 port map( A1 => n36254, A2 => REGISTERS_26_0_port, B1 => 
                           n36256, B2 => REGISTERS_21_0_port, ZN => n36228);
   U863 : AOI22_X1 port map( A1 => n36251, A2 => REGISTERS_1_0_port, B1 => 
                           n36252, B2 => REGISTERS_7_0_port, ZN => n36229);
   U864 : AOI222_X1 port map( A1 => n36248, A2 => REGISTERS_20_0_port, B1 => 
                           n36249, B2 => REGISTERS_5_0_port, C1 => n36247, C2 
                           => REGISTERS_18_0_port, ZN => n36230);
   U865 : NAND3_X1 port map( A1 => n36228, A2 => n36229, A3 => n36230, ZN => 
                           n36231);
   U866 : AOI22_X1 port map( A1 => n36244, A2 => REGISTERS_28_0_port, B1 => 
                           n36246, B2 => REGISTERS_19_0_port, ZN => n36232);
   U867 : AOI22_X1 port map( A1 => n36243, A2 => REGISTERS_6_0_port, B1 => 
                           n36257, B2 => REGISTERS_23_0_port, ZN => n36233);
   U868 : AOI22_X1 port map( A1 => n36253, A2 => REGISTERS_24_0_port, B1 => 
                           n36241, B2 => REGISTERS_10_0_port, ZN => n36234);
   U869 : AOI22_X1 port map( A1 => n36239, A2 => REGISTERS_12_0_port, B1 => 
                           n36266, B2 => REGISTERS_27_0_port, ZN => n36235);
   U870 : NAND4_X1 port map( A1 => n36232, A2 => n36233, A3 => n36234, A4 => 
                           n36235, ZN => n36236);
   U871 : OR4_X1 port map( A1 => n36222, A2 => n36227, A3 => n36231, A4 => 
                           n36236, ZN => OUTB(0));
   U872 : BUF_X2 port map( A => n36844, Z => n36237);
   U873 : BUF_X2 port map( A => n36845, Z => n36238);
   U874 : BUF_X2 port map( A => n36841, Z => n36239);
   U875 : BUF_X2 port map( A => n36843, Z => n36240);
   U876 : BUF_X2 port map( A => n36840, Z => n36241);
   U877 : BUF_X2 port map( A => n36846, Z => n36242);
   U878 : BUF_X2 port map( A => n36837, Z => n36243);
   U879 : BUF_X2 port map( A => n36835, Z => n36244);
   U880 : BUF_X2 port map( A => n36848, Z => n36245);
   U881 : BUF_X2 port map( A => n36836, Z => n36246);
   U882 : BUF_X2 port map( A => n36834, Z => n36247);
   U883 : BUF_X2 port map( A => n36832, Z => n36248);
   U884 : BUF_X2 port map( A => n36833, Z => n36249);
   U885 : BUF_X2 port map( A => n36847, Z => n36250);
   U886 : BUF_X2 port map( A => n36830, Z => n36251);
   U887 : BUF_X2 port map( A => n36831, Z => n36252);
   U888 : BUF_X2 port map( A => n36839, Z => n36253);
   U889 : BUF_X2 port map( A => n36828, Z => n36254);
   U890 : BUF_X2 port map( A => n36857, Z => n36255);
   U891 : BUF_X2 port map( A => n36829, Z => n36256);
   U892 : BUF_X2 port map( A => n36838, Z => n36257);
   U893 : BUF_X2 port map( A => n36850, Z => n36258);
   U894 : BUF_X2 port map( A => n36858, Z => n36259);
   U895 : BUF_X2 port map( A => n36849, Z => n36260);
   U896 : BUF_X2 port map( A => n36856, Z => n36261);
   U897 : BUF_X2 port map( A => n36851, Z => n36262);
   U898 : BUF_X2 port map( A => n36852, Z => n36263);
   U899 : BUF_X2 port map( A => n36854, Z => n36264);
   U900 : BUF_X2 port map( A => n36853, Z => n36265);
   U901 : BUF_X2 port map( A => n36842, Z => n36266);
   U902 : BUF_X2 port map( A => n36855, Z => n36267);
   U903 : NOR3_X2 port map( A1 => ADD_RDA(2), A2 => n36357, A3 => n36356, ZN =>
                           n36784);
   U904 : BUF_X1 port map( A => n36784, Z => n36286);
   U905 : BUF_X1 port map( A => n36771, Z => n36277);
   U906 : BUF_X1 port map( A => n36760, Z => n36270);
   U907 : BUF_X1 port map( A => n36800, Z => n36298);
   U908 : BUF_X1 port map( A => n36787, Z => n36289);
   U909 : BUF_X1 port map( A => n36788, Z => n36290);
   U910 : BUF_X1 port map( A => n36786, Z => n36288);
   U911 : BUF_X1 port map( A => n36782, Z => n36284);
   U912 : BUF_X1 port map( A => n36776, Z => n36282);
   U913 : BUF_X1 port map( A => n36763, Z => n36273);
   U914 : BUF_X1 port map( A => n36761, Z => n36271);
   U915 : BUF_X1 port map( A => n36759, Z => n36269);
   U916 : BUF_X1 port map( A => n36798, Z => n36296);
   U917 : BUF_X1 port map( A => n36796, Z => n36294);
   U918 : BUF_X1 port map( A => n36794, Z => n36292);
   U919 : BUF_X1 port map( A => n36772, Z => n36278);
   U920 : BUF_X1 port map( A => n36783, Z => n36285);
   U921 : BUF_X1 port map( A => n36764, Z => n36274);
   U922 : BUF_X1 port map( A => n36762, Z => n36272);
   U923 : BUF_X1 port map( A => n36775, Z => n36281);
   U924 : BUF_X1 port map( A => n36799, Z => n36297);
   U925 : BUF_X1 port map( A => n36797, Z => n36295);
   U926 : BUF_X1 port map( A => n36795, Z => n36293);
   U927 : BUF_X1 port map( A => n36793, Z => n36291);
   U928 : BUF_X1 port map( A => n36781, Z => n36283);
   U929 : BUF_X1 port map( A => n36773, Z => n36279);
   U930 : BUF_X1 port map( A => n36774, Z => n36280);
   U931 : BUF_X1 port map( A => n36769, Z => n36275);
   U932 : BUF_X1 port map( A => n36770, Z => n36276);
   U933 : BUF_X1 port map( A => n36758, Z => n36268);
   U934 : BUF_X1 port map( A => n36785, Z => n36287);
   U935 : INV_X1 port map( A => ADD_RDA(2), ZN => n36352);
   U936 : INV_X1 port map( A => ADD_RDA(4), ZN => n36350);
   U937 : INV_X1 port map( A => ADD_RDA(1), ZN => n36357);
   U938 : INV_X1 port map( A => ADD_RDB(3), ZN => n36810);
   U939 : OR4_X1 port map( A1 => n36717, A2 => n36716, A3 => n36715, A4 => 
                           n36714, ZN => OUTA(6));
   U940 : OR4_X1 port map( A1 => n36697, A2 => n36696, A3 => n36695, A4 => 
                           n36694, ZN => OUTA(5));
   U941 : OR4_X1 port map( A1 => n36657, A2 => n36656, A3 => n36655, A4 => 
                           n36654, ZN => OUTA(3));
   U942 : OR4_X1 port map( A1 => n36677, A2 => n36676, A3 => n36675, A4 => 
                           n36674, ZN => OUTA(4));
   U943 : OR4_X1 port map( A1 => n36637, A2 => n36636, A3 => n36635, A4 => 
                           n36634, ZN => OUTA(30));
   U944 : OR4_X1 port map( A1 => n36511, A2 => n36510, A3 => n36509, A4 => 
                           n36508, ZN => OUTA(1));
   U945 : OR4_X1 port map( A1 => n36427, A2 => n36426, A3 => n36425, A4 => 
                           n36424, ZN => OUTA(12));
   U946 : OR4_X1 port map( A1 => n36447, A2 => n36446, A3 => n36445, A4 => 
                           n36444, ZN => OUTA(13));
   U947 : OR4_X1 port map( A1 => n36387, A2 => n36386, A3 => n36385, A4 => 
                           n36384, ZN => OUTA(10));
   U948 : OR4_X1 port map( A1 => n36407, A2 => n36406, A3 => n36405, A4 => 
                           n36404, ZN => OUTA(11));
   U949 : OR4_X1 port map( A1 => n36467, A2 => n36466, A3 => n36465, A4 => 
                           n36464, ZN => OUTA(14));
   U950 : OR4_X1 port map( A1 => n36487, A2 => n36486, A3 => n36485, A4 => 
                           n36484, ZN => OUTA(15));
   U951 : OR4_X1 port map( A1 => n36737, A2 => n36736, A3 => n36735, A4 => 
                           n36734, ZN => OUTA(7));
   U952 : OR4_X1 port map( A1 => n36577, A2 => n36576, A3 => n36575, A4 => 
                           n36574, ZN => OUTA(28));
   U953 : OR4_X1 port map( A1 => n36537, A2 => n36536, A3 => n36535, A4 => 
                           n36534, ZN => OUTA(26));
   U954 : OR4_X1 port map( A1 => n36557, A2 => n36556, A3 => n36555, A4 => 
                           n36554, ZN => OUTA(27));
   U955 : OR4_X1 port map( A1 => n36617, A2 => n36616, A3 => n36615, A4 => 
                           n36614, ZN => OUTA(2));
   U956 : OR4_X1 port map( A1 => n36597, A2 => n36596, A3 => n36595, A4 => 
                           n36594, ZN => OUTA(29));
   U957 : OR4_X1 port map( A1 => n36757, A2 => n36756, A3 => n36755, A4 => 
                           n36754, ZN => OUTA(8));
   U958 : OR4_X1 port map( A1 => n36808, A2 => n36807, A3 => n36806, A4 => 
                           n36805, ZN => OUTA(9));
   U959 : NOR2_X1 port map( A1 => n36349, A2 => n36358, ZN => n36764);
   U960 : BUF_X1 port map( A => N288, Z => n36316);
   U961 : BUF_X1 port map( A => N300, Z => n36304);
   U962 : BUF_X1 port map( A => N287, Z => n36317);
   U963 : BUF_X1 port map( A => N283, Z => n36321);
   U964 : BUF_X1 port map( A => N284, Z => n36320);
   U965 : BUF_X1 port map( A => N285, Z => n36319);
   U966 : BUF_X1 port map( A => N301, Z => n36303);
   U967 : BUF_X1 port map( A => N286, Z => n36318);
   U968 : BUF_X1 port map( A => N293, Z => n36311);
   U969 : BUF_X1 port map( A => N294, Z => n36310);
   U970 : BUF_X1 port map( A => N295, Z => n36309);
   U971 : BUF_X1 port map( A => N296, Z => n36308);
   U972 : BUF_X1 port map( A => N289, Z => n36315);
   U973 : BUF_X1 port map( A => N299, Z => n36305);
   U974 : BUF_X1 port map( A => N290, Z => n36314);
   U975 : BUF_X1 port map( A => N291, Z => n36313);
   U976 : BUF_X1 port map( A => N298, Z => n36306);
   U977 : BUF_X1 port map( A => N297, Z => n36307);
   U978 : BUF_X1 port map( A => N292, Z => n36312);
   U979 : BUF_X1 port map( A => N276, Z => n36328);
   U980 : BUF_X1 port map( A => N277, Z => n36327);
   U981 : BUF_X1 port map( A => N305, Z => n36299);
   U982 : BUF_X1 port map( A => N243, Z => n36329);
   U983 : BUF_X1 port map( A => N278, Z => n36326);
   U984 : BUF_X1 port map( A => N302, Z => n36302);
   U985 : BUF_X1 port map( A => N303, Z => n36301);
   U986 : BUF_X1 port map( A => N304, Z => n36300);
   U987 : BUF_X1 port map( A => N282, Z => n36322);
   U988 : BUF_X1 port map( A => N281, Z => n36323);
   U989 : BUF_X1 port map( A => N280, Z => n36324);
   U990 : INV_X1 port map( A => ADD_WR(0), ZN => n36332);
   U991 : BUF_X1 port map( A => N279, Z => n36325);
   U992 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(6), ZN => N250);
   U993 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(5), ZN => N249);
   U994 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(3), ZN => N247);
   U995 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(17), ZN => N261);
   U996 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(18), ZN => N262);
   U997 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(19), ZN => N263);
   U998 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(16), ZN => N260);
   U999 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(15), ZN => N259);
   U1000 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(14), ZN => N258);
   U1001 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(13), ZN => N257);
   U1002 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(24), ZN => N268);
   U1003 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(20), ZN => N264);
   U1004 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(12), ZN => N256);
   U1005 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(11), ZN => N255);
   U1006 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(10), ZN => N254);
   U1007 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(9), ZN => N253);
   U1008 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(8), ZN => N252);
   U1009 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(7), ZN => N251);
   U1010 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(27), ZN => N271);
   U1011 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(26), ZN => N270);
   U1012 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(4), ZN => N248);
   U1013 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(30), ZN => N274);
   U1014 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(2), ZN => N246);
   U1015 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(1), ZN => N245);
   U1016 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(0), ZN => N244);
   U1017 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(31), ZN => N275);
   U1018 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(25), ZN => N269);
   U1019 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(29), ZN => N273);
   U1020 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(28), ZN => N272);
   U1021 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(22), ZN => N266);
   U1022 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(21), ZN => N265);
   U1023 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(23), ZN => N267);
   U1024 : NOR2_X1 port map( A1 => n36823, A2 => n36826, ZN => n36855);
   U1025 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => ADD_WR(2)
                           , ZN => n36340);
   U1026 : NAND3_X1 port map( A1 => WE, A2 => ADD_WR(3), A3 => ADD_WR(4), ZN =>
                           n36334);
   U1027 : OAI21_X1 port map( B1 => n36340, B2 => n36334, A => RESET, ZN => 
                           N243);
   U1028 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n36332, 
                           ZN => n36341);
   U1029 : OAI21_X1 port map( B1 => n36334, B2 => n36341, A => RESET, ZN => 
                           N276);
   U1030 : INV_X1 port map( A => ADD_WR(1), ZN => n36330);
   U1031 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n36330, 
                           ZN => n36342);
   U1032 : OAI21_X1 port map( B1 => n36334, B2 => n36342, A => RESET, ZN => 
                           N277);
   U1033 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n36332, A3 => n36330, ZN 
                           => n36343);
   U1034 : OAI21_X1 port map( B1 => n36334, B2 => n36343, A => RESET, ZN => 
                           N278);
   U1035 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n36330, ZN => n36331);
   U1036 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n36331, ZN => n36344);
   U1037 : OAI21_X1 port map( B1 => n36334, B2 => n36344, A => RESET, ZN => 
                           N279);
   U1038 : NAND2_X1 port map( A1 => n36331, A2 => n36332, ZN => n36345);
   U1039 : OAI21_X1 port map( B1 => n36334, B2 => n36345, A => RESET, ZN => 
                           N280);
   U1040 : NOR2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), ZN => n36333);
   U1041 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n36333, ZN => n36347);
   U1042 : OAI21_X1 port map( B1 => n36334, B2 => n36347, A => RESET, ZN => 
                           N281);
   U1043 : NAND2_X1 port map( A1 => n36333, A2 => n36332, ZN => n36337);
   U1044 : OAI21_X1 port map( B1 => n36334, B2 => n36337, A => RESET, ZN => 
                           N282);
   U1045 : INV_X1 port map( A => ADD_WR(3), ZN => n36339);
   U1046 : NAND3_X1 port map( A1 => WE, A2 => ADD_WR(4), A3 => n36339, ZN => 
                           n36335);
   U1047 : OAI21_X1 port map( B1 => n36340, B2 => n36335, A => RESET, ZN => 
                           N283);
   U1048 : OAI21_X1 port map( B1 => n36341, B2 => n36335, A => RESET, ZN => 
                           N284);
   U1049 : OAI21_X1 port map( B1 => n36342, B2 => n36335, A => RESET, ZN => 
                           N285);
   U1050 : OAI21_X1 port map( B1 => n36343, B2 => n36335, A => RESET, ZN => 
                           N286);
   U1051 : OAI21_X1 port map( B1 => n36344, B2 => n36335, A => RESET, ZN => 
                           N287);
   U1052 : OAI21_X1 port map( B1 => n36345, B2 => n36335, A => RESET, ZN => 
                           N288);
   U1053 : OAI21_X1 port map( B1 => n36347, B2 => n36335, A => RESET, ZN => 
                           N289);
   U1054 : OAI21_X1 port map( B1 => n36337, B2 => n36335, A => RESET, ZN => 
                           N290);
   U1055 : INV_X1 port map( A => ADD_WR(4), ZN => n36338);
   U1056 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => WE, A3 => n36338, ZN => 
                           n36336);
   U1057 : OAI21_X1 port map( B1 => n36340, B2 => n36336, A => RESET, ZN => 
                           N291);
   U1058 : OAI21_X1 port map( B1 => n36341, B2 => n36336, A => RESET, ZN => 
                           N292);
   U1059 : OAI21_X1 port map( B1 => n36342, B2 => n36336, A => RESET, ZN => 
                           N293);
   U1060 : OAI21_X1 port map( B1 => n36343, B2 => n36336, A => RESET, ZN => 
                           N294);
   U1061 : OAI21_X1 port map( B1 => n36344, B2 => n36336, A => RESET, ZN => 
                           N295);
   U1062 : OAI21_X1 port map( B1 => n36345, B2 => n36336, A => RESET, ZN => 
                           N296);
   U1063 : OAI21_X1 port map( B1 => n36347, B2 => n36336, A => RESET, ZN => 
                           N297);
   U1064 : OAI21_X1 port map( B1 => n36337, B2 => n36336, A => RESET, ZN => 
                           N298);
   U1065 : NAND3_X1 port map( A1 => WE, A2 => n36339, A3 => n36338, ZN => 
                           n36346);
   U1066 : OAI21_X1 port map( B1 => n36340, B2 => n36346, A => RESET, ZN => 
                           N299);
   U1067 : OAI21_X1 port map( B1 => n36341, B2 => n36346, A => RESET, ZN => 
                           N300);
   U1068 : OAI21_X1 port map( B1 => n36342, B2 => n36346, A => RESET, ZN => 
                           N301);
   U1069 : OAI21_X1 port map( B1 => n36343, B2 => n36346, A => RESET, ZN => 
                           N302);
   U1070 : OAI21_X1 port map( B1 => n36344, B2 => n36346, A => RESET, ZN => 
                           N303);
   U1071 : OAI21_X1 port map( B1 => n36345, B2 => n36346, A => RESET, ZN => 
                           N304);
   U1072 : OAI21_X1 port map( B1 => n36347, B2 => n36346, A => RESET, ZN => 
                           N305);
   U1073 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDA(2), A3 => n36357, ZN 
                           => n36365);
   U1074 : INV_X1 port map( A => ADD_RDA(3), ZN => n36348);
   U1075 : NAND3_X1 port map( A1 => ADD_RDA(0), A2 => n36350, A3 => n36348, ZN 
                           => n36360);
   U1076 : NOR2_X1 port map( A1 => n36365, A2 => n36360, ZN => n36759);
   U1077 : NOR2_X1 port map( A1 => ADD_RDA(3), A2 => ADD_RDA(0), ZN => n36351);
   U1078 : NAND2_X1 port map( A1 => ADD_RDA(4), A2 => n36351, ZN => n36364);
   U1079 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDA(1), A3 => ADD_RDA(2), 
                           ZN => n36367);
   U1080 : NOR2_X1 port map( A1 => n36364, A2 => n36367, ZN => n36758);
   U1081 : NAND3_X1 port map( A1 => ADD_RDA(4), A2 => ADD_RDA(3), A3 => 
                           ADD_RDA(0), ZN => n36359);
   U1082 : NAND3_X1 port map( A1 => RESET, A2 => n36357, A3 => n36352, ZN => 
                           n36363);
   U1083 : NOR2_X1 port map( A1 => n36359, A2 => n36363, ZN => n36761);
   U1084 : NAND3_X1 port map( A1 => ADD_RDA(4), A2 => ADD_RDA(0), A3 => n36348,
                           ZN => n36349);
   U1085 : NOR2_X1 port map( A1 => n36349, A2 => n36365, ZN => n36760);
   U1086 : NOR2_X1 port map( A1 => n36349, A2 => n36363, ZN => n36763);
   U1087 : NOR2_X1 port map( A1 => n36349, A2 => n36367, ZN => n36762);
   U1088 : NAND3_X1 port map( A1 => ADD_RDA(1), A2 => RESET, A3 => n36352, ZN 
                           => n36358);
   U1089 : INV_X1 port map( A => ADD_RDA(0), ZN => n36354);
   U1090 : NAND3_X1 port map( A1 => ADD_RDA(3), A2 => n36350, A3 => n36354, ZN 
                           => n36361);
   U1091 : NOR2_X1 port map( A1 => n36367, A2 => n36361, ZN => n36770);
   U1092 : NAND3_X1 port map( A1 => ADD_RDA(3), A2 => ADD_RDA(0), A3 => n36350,
                           ZN => n36366);
   U1093 : NOR2_X1 port map( A1 => n36365, A2 => n36366, ZN => n36769);
   U1094 : NOR2_X1 port map( A1 => n36358, A2 => n36359, ZN => n36772);
   U1095 : NAND3_X1 port map( A1 => RESET, A2 => n36351, A3 => n36350, ZN => 
                           n36356);
   U1096 : NOR3_X1 port map( A1 => ADD_RDA(1), A2 => n36352, A3 => n36356, ZN 
                           => n36771);
   U1097 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n36278, B1 => 
                           REGISTERS_4_0_port, B2 => n36277, ZN => n36355);
   U1098 : NAND2_X1 port map( A1 => ADD_RDA(1), A2 => ADD_RDA(2), ZN => n36353)
                           ;
   U1099 : NOR2_X1 port map( A1 => n36353, A2 => n36356, ZN => n36774);
   U1100 : NAND3_X1 port map( A1 => ADD_RDA(3), A2 => ADD_RDA(4), A3 => n36354,
                           ZN => n36362);
   U1101 : NOR2_X1 port map( A1 => n36365, A2 => n36362, ZN => n36773);
   U1102 : NOR2_X1 port map( A1 => n36358, A2 => n36362, ZN => n36776);
   U1103 : NOR2_X1 port map( A1 => n36360, A2 => n36367, ZN => n36775);
   U1104 : NOR2_X1 port map( A1 => n36358, A2 => n36361, ZN => n36782);
   U1105 : NOR2_X1 port map( A1 => n36363, A2 => n36366, ZN => n36781);
   U1106 : NOR2_X1 port map( A1 => n36358, A2 => n36364, ZN => n36783);
   U1107 : NOR2_X1 port map( A1 => n36358, A2 => n36360, ZN => n36786);
   U1108 : NOR2_X1 port map( A1 => n36367, A2 => n36359, ZN => n36785);
   U1109 : NOR2_X1 port map( A1 => n36367, A2 => n36362, ZN => n36788);
   U1110 : NOR2_X1 port map( A1 => n36363, A2 => n36361, ZN => n36787);
   U1111 : NOR2_X1 port map( A1 => n36358, A2 => n36366, ZN => n36794);
   U1112 : NOR2_X1 port map( A1 => n36365, A2 => n36359, ZN => n36793);
   U1113 : NOR2_X1 port map( A1 => n36360, A2 => n36363, ZN => n36796);
   U1114 : NOR2_X1 port map( A1 => n36364, A2 => n36363, ZN => n36795);
   U1115 : NOR2_X1 port map( A1 => n36365, A2 => n36361, ZN => n36798);
   U1116 : NOR2_X1 port map( A1 => n36363, A2 => n36362, ZN => n36797);
   U1117 : NOR2_X1 port map( A1 => n36365, A2 => n36364, ZN => n36800);
   U1118 : NOR2_X1 port map( A1 => n36367, A2 => n36366, ZN => n36799);
   U1119 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_10_port, B1 => 
                           n36268, B2 => REGISTERS_22_10_port, ZN => n36371);
   U1120 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_10_port, B1 => 
                           n36270, B2 => REGISTERS_21_10_port, ZN => n36370);
   U1121 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_10_port, B1 => 
                           n36272, B2 => REGISTERS_23_10_port, ZN => n36369);
   U1122 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_10_port, ZN => 
                           n36368);
   U1123 : NAND4_X1 port map( A1 => n36371, A2 => n36370, A3 => n36369, A4 => 
                           n36368, ZN => n36387);
   U1124 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_10_port, B1 => 
                           n36275, B2 => REGISTERS_13_10_port, ZN => n36375);
   U1125 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_10_port, B1 => 
                           n36277, B2 => REGISTERS_4_10_port, ZN => n36374);
   U1126 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_10_port, B1 => 
                           n36279, B2 => REGISTERS_28_10_port, ZN => n36373);
   U1127 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_10_port, B1 => 
                           n36281, B2 => REGISTERS_7_10_port, ZN => n36372);
   U1128 : NAND4_X1 port map( A1 => n36375, A2 => n36374, A3 => n36373, A4 => 
                           n36372, ZN => n36386);
   U1129 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_10_port, B1 => 
                           n36283, B2 => REGISTERS_9_10_port, ZN => n36379);
   U1130 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_10_port, B1 => 
                           n36285, B2 => REGISTERS_18_10_port, ZN => n36378);
   U1131 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_10_port, B1 => 
                           n36287, B2 => REGISTERS_31_10_port, ZN => n36377);
   U1132 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_10_port, B1 => 
                           n36289, B2 => REGISTERS_8_10_port, ZN => n36376);
   U1133 : NAND4_X1 port map( A1 => n36379, A2 => n36378, A3 => n36377, A4 => 
                           n36376, ZN => n36385);
   U1134 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_10_port, B1 => 
                           n36291, B2 => REGISTERS_29_10_port, ZN => n36383);
   U1135 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_10_port, B1 => 
                           n36293, B2 => REGISTERS_16_10_port, ZN => n36382);
   U1136 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_10_port, B1 => 
                           n36295, B2 => REGISTERS_24_10_port, ZN => n36381);
   U1137 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_10_port, B1 => 
                           n36297, B2 => REGISTERS_15_10_port, ZN => n36380);
   U1138 : NAND4_X1 port map( A1 => n36383, A2 => n36382, A3 => n36381, A4 => 
                           n36380, ZN => n36384);
   U1139 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_11_port, B1 => 
                           n36268, B2 => REGISTERS_22_11_port, ZN => n36391);
   U1140 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_11_port, B1 => 
                           n36270, B2 => REGISTERS_21_11_port, ZN => n36390);
   U1141 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_11_port, B1 => 
                           n36272, B2 => REGISTERS_23_11_port, ZN => n36389);
   U1142 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_11_port, ZN => 
                           n36388);
   U1143 : NAND4_X1 port map( A1 => n36391, A2 => n36390, A3 => n36389, A4 => 
                           n36388, ZN => n36407);
   U1144 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_11_port, B1 => 
                           n36275, B2 => REGISTERS_13_11_port, ZN => n36395);
   U1145 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_11_port, B1 => 
                           n36277, B2 => REGISTERS_4_11_port, ZN => n36394);
   U1146 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_11_port, B1 => 
                           n36279, B2 => REGISTERS_28_11_port, ZN => n36393);
   U1147 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_11_port, B1 => 
                           n36281, B2 => REGISTERS_7_11_port, ZN => n36392);
   U1148 : NAND4_X1 port map( A1 => n36395, A2 => n36394, A3 => n36393, A4 => 
                           n36392, ZN => n36406);
   U1149 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_11_port, B1 => 
                           n36283, B2 => REGISTERS_9_11_port, ZN => n36399);
   U1150 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_11_port, B1 => 
                           n36285, B2 => REGISTERS_18_11_port, ZN => n36398);
   U1151 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_11_port, B1 => 
                           n36287, B2 => REGISTERS_31_11_port, ZN => n36397);
   U1152 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_11_port, B1 => 
                           n36289, B2 => REGISTERS_8_11_port, ZN => n36396);
   U1153 : NAND4_X1 port map( A1 => n36399, A2 => n36398, A3 => n36397, A4 => 
                           n36396, ZN => n36405);
   U1154 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_11_port, B1 => 
                           n36291, B2 => REGISTERS_29_11_port, ZN => n36403);
   U1155 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_11_port, B1 => 
                           n36293, B2 => REGISTERS_16_11_port, ZN => n36402);
   U1156 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_11_port, B1 => 
                           n36295, B2 => REGISTERS_24_11_port, ZN => n36401);
   U1157 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_11_port, B1 => 
                           n36297, B2 => REGISTERS_15_11_port, ZN => n36400);
   U1158 : NAND4_X1 port map( A1 => n36403, A2 => n36402, A3 => n36401, A4 => 
                           n36400, ZN => n36404);
   U1159 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_12_port, B1 => 
                           n36268, B2 => REGISTERS_22_12_port, ZN => n36411);
   U1160 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_12_port, B1 => 
                           n36270, B2 => REGISTERS_21_12_port, ZN => n36410);
   U1161 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_12_port, B1 => 
                           n36272, B2 => REGISTERS_23_12_port, ZN => n36409);
   U1162 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_12_port, ZN => 
                           n36408);
   U1163 : NAND4_X1 port map( A1 => n36411, A2 => n36410, A3 => n36409, A4 => 
                           n36408, ZN => n36427);
   U1164 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_12_port, B1 => 
                           n36275, B2 => REGISTERS_13_12_port, ZN => n36415);
   U1165 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_12_port, B1 => 
                           n36277, B2 => REGISTERS_4_12_port, ZN => n36414);
   U1166 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_12_port, B1 => 
                           n36279, B2 => REGISTERS_28_12_port, ZN => n36413);
   U1167 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_12_port, B1 => 
                           n36281, B2 => REGISTERS_7_12_port, ZN => n36412);
   U1168 : NAND4_X1 port map( A1 => n36415, A2 => n36414, A3 => n36413, A4 => 
                           n36412, ZN => n36426);
   U1169 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_12_port, B1 => 
                           n36283, B2 => REGISTERS_9_12_port, ZN => n36419);
   U1170 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_12_port, B1 => 
                           n36285, B2 => REGISTERS_18_12_port, ZN => n36418);
   U1171 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_12_port, B1 => 
                           n36287, B2 => REGISTERS_31_12_port, ZN => n36417);
   U1172 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_12_port, B1 => 
                           n36289, B2 => REGISTERS_8_12_port, ZN => n36416);
   U1173 : NAND4_X1 port map( A1 => n36419, A2 => n36418, A3 => n36417, A4 => 
                           n36416, ZN => n36425);
   U1174 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_12_port, B1 => 
                           n36291, B2 => REGISTERS_29_12_port, ZN => n36423);
   U1175 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_12_port, B1 => 
                           n36293, B2 => REGISTERS_16_12_port, ZN => n36422);
   U1176 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_12_port, B1 => 
                           n36295, B2 => REGISTERS_24_12_port, ZN => n36421);
   U1177 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_12_port, B1 => 
                           n36297, B2 => REGISTERS_15_12_port, ZN => n36420);
   U1178 : NAND4_X1 port map( A1 => n36423, A2 => n36422, A3 => n36421, A4 => 
                           n36420, ZN => n36424);
   U1179 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_13_port, B1 => 
                           n36268, B2 => REGISTERS_22_13_port, ZN => n36431);
   U1180 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_13_port, B1 => 
                           n36270, B2 => REGISTERS_21_13_port, ZN => n36430);
   U1181 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_13_port, B1 => 
                           n36272, B2 => REGISTERS_23_13_port, ZN => n36429);
   U1182 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_13_port, ZN => 
                           n36428);
   U1183 : NAND4_X1 port map( A1 => n36431, A2 => n36430, A3 => n36429, A4 => 
                           n36428, ZN => n36447);
   U1184 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_13_port, B1 => 
                           n36275, B2 => REGISTERS_13_13_port, ZN => n36435);
   U1185 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_13_port, B1 => 
                           n36277, B2 => REGISTERS_4_13_port, ZN => n36434);
   U1186 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_13_port, B1 => 
                           n36279, B2 => REGISTERS_28_13_port, ZN => n36433);
   U1187 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_13_port, B1 => 
                           n36281, B2 => REGISTERS_7_13_port, ZN => n36432);
   U1188 : NAND4_X1 port map( A1 => n36435, A2 => n36434, A3 => n36433, A4 => 
                           n36432, ZN => n36446);
   U1189 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_13_port, B1 => 
                           n36283, B2 => REGISTERS_9_13_port, ZN => n36439);
   U1190 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_13_port, B1 => 
                           n36285, B2 => REGISTERS_18_13_port, ZN => n36438);
   U1191 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_13_port, B1 => 
                           n36287, B2 => REGISTERS_31_13_port, ZN => n36437);
   U1192 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_13_port, B1 => 
                           n36289, B2 => REGISTERS_8_13_port, ZN => n36436);
   U1193 : NAND4_X1 port map( A1 => n36439, A2 => n36438, A3 => n36437, A4 => 
                           n36436, ZN => n36445);
   U1194 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_13_port, B1 => 
                           n36291, B2 => REGISTERS_29_13_port, ZN => n36443);
   U1195 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_13_port, B1 => 
                           n36293, B2 => REGISTERS_16_13_port, ZN => n36442);
   U1196 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_13_port, B1 => 
                           n36295, B2 => REGISTERS_24_13_port, ZN => n36441);
   U1197 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_13_port, B1 => 
                           n36297, B2 => REGISTERS_15_13_port, ZN => n36440);
   U1198 : NAND4_X1 port map( A1 => n36443, A2 => n36442, A3 => n36441, A4 => 
                           n36440, ZN => n36444);
   U1199 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_14_port, B1 => 
                           n36268, B2 => REGISTERS_22_14_port, ZN => n36451);
   U1200 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_14_port, B1 => 
                           n36270, B2 => REGISTERS_21_14_port, ZN => n36450);
   U1201 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_14_port, B1 => 
                           n36272, B2 => REGISTERS_23_14_port, ZN => n36449);
   U1202 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_14_port, ZN => 
                           n36448);
   U1203 : NAND4_X1 port map( A1 => n36451, A2 => n36450, A3 => n36449, A4 => 
                           n36448, ZN => n36467);
   U1204 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_14_port, B1 => 
                           n36275, B2 => REGISTERS_13_14_port, ZN => n36455);
   U1205 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_14_port, B1 => 
                           n36277, B2 => REGISTERS_4_14_port, ZN => n36454);
   U1206 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_14_port, B1 => 
                           n36279, B2 => REGISTERS_28_14_port, ZN => n36453);
   U1207 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_14_port, B1 => 
                           n36281, B2 => REGISTERS_7_14_port, ZN => n36452);
   U1208 : NAND4_X1 port map( A1 => n36455, A2 => n36454, A3 => n36453, A4 => 
                           n36452, ZN => n36466);
   U1209 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_14_port, B1 => 
                           n36283, B2 => REGISTERS_9_14_port, ZN => n36459);
   U1210 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_14_port, B1 => 
                           n36285, B2 => REGISTERS_18_14_port, ZN => n36458);
   U1211 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_14_port, B1 => 
                           n36287, B2 => REGISTERS_31_14_port, ZN => n36457);
   U1212 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_14_port, B1 => 
                           n36289, B2 => REGISTERS_8_14_port, ZN => n36456);
   U1213 : NAND4_X1 port map( A1 => n36459, A2 => n36458, A3 => n36457, A4 => 
                           n36456, ZN => n36465);
   U1214 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_14_port, B1 => 
                           n36291, B2 => REGISTERS_29_14_port, ZN => n36463);
   U1215 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_14_port, B1 => 
                           n36293, B2 => REGISTERS_16_14_port, ZN => n36462);
   U1216 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_14_port, B1 => 
                           n36295, B2 => REGISTERS_24_14_port, ZN => n36461);
   U1217 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_14_port, B1 => 
                           n36297, B2 => REGISTERS_15_14_port, ZN => n36460);
   U1218 : NAND4_X1 port map( A1 => n36463, A2 => n36462, A3 => n36461, A4 => 
                           n36460, ZN => n36464);
   U1219 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_15_port, B1 => 
                           n36268, B2 => REGISTERS_22_15_port, ZN => n36471);
   U1220 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_15_port, B1 => 
                           n36270, B2 => REGISTERS_21_15_port, ZN => n36470);
   U1221 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_15_port, B1 => 
                           n36272, B2 => REGISTERS_23_15_port, ZN => n36469);
   U1222 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_15_port, ZN => 
                           n36468);
   U1223 : NAND4_X1 port map( A1 => n36471, A2 => n36470, A3 => n36469, A4 => 
                           n36468, ZN => n36487);
   U1224 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_15_port, B1 => 
                           n36275, B2 => REGISTERS_13_15_port, ZN => n36475);
   U1225 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_15_port, B1 => 
                           n36277, B2 => REGISTERS_4_15_port, ZN => n36474);
   U1226 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_15_port, B1 => 
                           n36279, B2 => REGISTERS_28_15_port, ZN => n36473);
   U1227 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_15_port, B1 => 
                           n36281, B2 => REGISTERS_7_15_port, ZN => n36472);
   U1228 : NAND4_X1 port map( A1 => n36475, A2 => n36474, A3 => n36473, A4 => 
                           n36472, ZN => n36486);
   U1229 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_15_port, B1 => 
                           n36283, B2 => REGISTERS_9_15_port, ZN => n36479);
   U1230 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_15_port, B1 => 
                           n36285, B2 => REGISTERS_18_15_port, ZN => n36478);
   U1231 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_15_port, B1 => 
                           n36287, B2 => REGISTERS_31_15_port, ZN => n36477);
   U1232 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_15_port, B1 => 
                           n36289, B2 => REGISTERS_8_15_port, ZN => n36476);
   U1233 : NAND4_X1 port map( A1 => n36479, A2 => n36478, A3 => n36477, A4 => 
                           n36476, ZN => n36485);
   U1234 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_15_port, B1 => 
                           n36291, B2 => REGISTERS_29_15_port, ZN => n36483);
   U1235 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_15_port, B1 => 
                           n36293, B2 => REGISTERS_16_15_port, ZN => n36482);
   U1236 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_15_port, B1 => 
                           n36295, B2 => REGISTERS_24_15_port, ZN => n36481);
   U1237 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_15_port, B1 => 
                           n36297, B2 => REGISTERS_15_15_port, ZN => n36480);
   U1238 : NAND4_X1 port map( A1 => n36483, A2 => n36482, A3 => n36481, A4 => 
                           n36480, ZN => n36484);
   U1239 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_16_port, B1 => 
                           n36277, B2 => REGISTERS_4_16_port, ZN => n36488);
   U1240 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_17_port, B1 => 
                           n36277, B2 => REGISTERS_4_17_port, ZN => n36489);
   U1241 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_18_port, B1 => 
                           n36277, B2 => REGISTERS_4_18_port, ZN => n36490);
   U1242 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_19_port, B1 => 
                           n36277, B2 => REGISTERS_4_19_port, ZN => n36491);
   U1243 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_1_port, B1 => 
                           n36268, B2 => REGISTERS_22_1_port, ZN => n36495);
   U1244 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_1_port, B1 => 
                           n36270, B2 => REGISTERS_21_1_port, ZN => n36494);
   U1245 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_1_port, B1 => 
                           n36272, B2 => REGISTERS_23_1_port, ZN => n36493);
   U1246 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_1_port, ZN => 
                           n36492);
   U1247 : NAND4_X1 port map( A1 => n36495, A2 => n36494, A3 => n36493, A4 => 
                           n36492, ZN => n36511);
   U1248 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_1_port, B1 => 
                           n36275, B2 => REGISTERS_13_1_port, ZN => n36499);
   U1249 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_1_port, B1 => 
                           n36277, B2 => REGISTERS_4_1_port, ZN => n36498);
   U1250 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_1_port, B1 => 
                           n36279, B2 => REGISTERS_28_1_port, ZN => n36497);
   U1251 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_1_port, B1 => 
                           n36281, B2 => REGISTERS_7_1_port, ZN => n36496);
   U1252 : NAND4_X1 port map( A1 => n36499, A2 => n36498, A3 => n36497, A4 => 
                           n36496, ZN => n36510);
   U1253 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_1_port, B1 => 
                           n36283, B2 => REGISTERS_9_1_port, ZN => n36503);
   U1254 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_1_port, B1 => 
                           n36285, B2 => REGISTERS_18_1_port, ZN => n36502);
   U1255 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_1_port, B1 => 
                           n36287, B2 => REGISTERS_31_1_port, ZN => n36501);
   U1256 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_1_port, B1 => 
                           n36289, B2 => REGISTERS_8_1_port, ZN => n36500);
   U1257 : NAND4_X1 port map( A1 => n36503, A2 => n36502, A3 => n36501, A4 => 
                           n36500, ZN => n36509);
   U1258 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_1_port, B1 => 
                           n36291, B2 => REGISTERS_29_1_port, ZN => n36507);
   U1259 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_1_port, B1 => 
                           n36293, B2 => REGISTERS_16_1_port, ZN => n36506);
   U1260 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_1_port, B1 => 
                           n36295, B2 => REGISTERS_24_1_port, ZN => n36505);
   U1261 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_1_port, B1 => 
                           n36297, B2 => REGISTERS_15_1_port, ZN => n36504);
   U1262 : NAND4_X1 port map( A1 => n36507, A2 => n36506, A3 => n36505, A4 => 
                           n36504, ZN => n36508);
   U1263 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_20_port, B1 => 
                           n36277, B2 => REGISTERS_4_20_port, ZN => n36512);
   U1264 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_21_port, B1 => 
                           n36277, B2 => REGISTERS_4_21_port, ZN => n36513);
   U1265 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_22_port, B1 => 
                           n36277, B2 => REGISTERS_4_22_port, ZN => n36514);
   U1266 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_23_port, B1 => 
                           n36277, B2 => REGISTERS_4_23_port, ZN => n36515);
   U1267 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_24_port, B1 => 
                           n36277, B2 => REGISTERS_4_24_port, ZN => n36516);
   U1268 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_25_port, B1 => 
                           n36277, B2 => REGISTERS_4_25_port, ZN => n36517);
   U1269 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_26_port, B1 => 
                           n36758, B2 => REGISTERS_22_26_port, ZN => n36521);
   U1270 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_26_port, B1 => 
                           n36760, B2 => REGISTERS_21_26_port, ZN => n36520);
   U1271 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_26_port, B1 => 
                           n36762, B2 => REGISTERS_23_26_port, ZN => n36519);
   U1272 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_26_port, ZN => 
                           n36518);
   U1273 : NAND4_X1 port map( A1 => n36521, A2 => n36520, A3 => n36519, A4 => 
                           n36518, ZN => n36537);
   U1274 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_26_port, B1 => 
                           n36275, B2 => REGISTERS_13_26_port, ZN => n36525);
   U1275 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_26_port, B1 => 
                           n36277, B2 => REGISTERS_4_26_port, ZN => n36524);
   U1276 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_26_port, B1 => 
                           n36279, B2 => REGISTERS_28_26_port, ZN => n36523);
   U1277 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_26_port, B1 => 
                           n36775, B2 => REGISTERS_7_26_port, ZN => n36522);
   U1278 : NAND4_X1 port map( A1 => n36525, A2 => n36524, A3 => n36523, A4 => 
                           n36522, ZN => n36536);
   U1279 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_26_port, B1 => 
                           n36283, B2 => REGISTERS_9_26_port, ZN => n36529);
   U1280 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_26_port, B1 => 
                           n36783, B2 => REGISTERS_18_26_port, ZN => n36528);
   U1281 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_26_port, B1 => 
                           n36785, B2 => REGISTERS_31_26_port, ZN => n36527);
   U1282 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_26_port, B1 => 
                           n36289, B2 => REGISTERS_8_26_port, ZN => n36526);
   U1283 : NAND4_X1 port map( A1 => n36529, A2 => n36528, A3 => n36527, A4 => 
                           n36526, ZN => n36535);
   U1284 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_26_port, B1 => 
                           n36291, B2 => REGISTERS_29_26_port, ZN => n36533);
   U1285 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_26_port, B1 => 
                           n36293, B2 => REGISTERS_16_26_port, ZN => n36532);
   U1286 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_26_port, B1 => 
                           n36295, B2 => REGISTERS_24_26_port, ZN => n36531);
   U1287 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_26_port, B1 => 
                           n36297, B2 => REGISTERS_15_26_port, ZN => n36530);
   U1288 : NAND4_X1 port map( A1 => n36533, A2 => n36532, A3 => n36531, A4 => 
                           n36530, ZN => n36534);
   U1289 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_27_port, B1 => 
                           n36758, B2 => REGISTERS_22_27_port, ZN => n36541);
   U1290 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_27_port, B1 => 
                           n36760, B2 => REGISTERS_21_27_port, ZN => n36540);
   U1291 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_27_port, B1 => 
                           n36762, B2 => REGISTERS_23_27_port, ZN => n36539);
   U1292 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_27_port, ZN => 
                           n36538);
   U1293 : NAND4_X1 port map( A1 => n36541, A2 => n36540, A3 => n36539, A4 => 
                           n36538, ZN => n36557);
   U1294 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_27_port, B1 => 
                           n36769, B2 => REGISTERS_13_27_port, ZN => n36545);
   U1295 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_27_port, B1 => 
                           n36277, B2 => REGISTERS_4_27_port, ZN => n36544);
   U1296 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_27_port, B1 => 
                           n36773, B2 => REGISTERS_28_27_port, ZN => n36543);
   U1297 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_27_port, B1 => 
                           n36775, B2 => REGISTERS_7_27_port, ZN => n36542);
   U1298 : NAND4_X1 port map( A1 => n36545, A2 => n36544, A3 => n36543, A4 => 
                           n36542, ZN => n36556);
   U1299 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_27_port, B1 => 
                           n36781, B2 => REGISTERS_9_27_port, ZN => n36549);
   U1300 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_27_port, B1 => 
                           n36783, B2 => REGISTERS_18_27_port, ZN => n36548);
   U1301 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_27_port, B1 => 
                           n36785, B2 => REGISTERS_31_27_port, ZN => n36547);
   U1302 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_27_port, B1 => 
                           n36787, B2 => REGISTERS_8_27_port, ZN => n36546);
   U1303 : NAND4_X1 port map( A1 => n36549, A2 => n36548, A3 => n36547, A4 => 
                           n36546, ZN => n36555);
   U1304 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_27_port, B1 => 
                           n36793, B2 => REGISTERS_29_27_port, ZN => n36553);
   U1305 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_27_port, B1 => 
                           n36795, B2 => REGISTERS_16_27_port, ZN => n36552);
   U1306 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_27_port, B1 => 
                           n36797, B2 => REGISTERS_24_27_port, ZN => n36551);
   U1307 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_27_port, B1 => 
                           n36799, B2 => REGISTERS_15_27_port, ZN => n36550);
   U1308 : NAND4_X1 port map( A1 => n36553, A2 => n36552, A3 => n36551, A4 => 
                           n36550, ZN => n36554);
   U1309 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_28_port, B1 => 
                           n36758, B2 => REGISTERS_22_28_port, ZN => n36561);
   U1310 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_28_port, B1 => 
                           n36270, B2 => REGISTERS_21_28_port, ZN => n36560);
   U1311 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_28_port, B1 => 
                           n36762, B2 => REGISTERS_23_28_port, ZN => n36559);
   U1312 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_28_port, ZN => 
                           n36558);
   U1313 : NAND4_X1 port map( A1 => n36561, A2 => n36560, A3 => n36559, A4 => 
                           n36558, ZN => n36577);
   U1314 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_28_port, B1 => 
                           n36769, B2 => REGISTERS_13_28_port, ZN => n36565);
   U1315 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_28_port, B1 => 
                           n36277, B2 => REGISTERS_4_28_port, ZN => n36564);
   U1316 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_28_port, B1 => 
                           n36773, B2 => REGISTERS_28_28_port, ZN => n36563);
   U1317 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_28_port, B1 => 
                           n36281, B2 => REGISTERS_7_28_port, ZN => n36562);
   U1318 : NAND4_X1 port map( A1 => n36565, A2 => n36564, A3 => n36563, A4 => 
                           n36562, ZN => n36576);
   U1319 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_28_port, B1 => 
                           n36781, B2 => REGISTERS_9_28_port, ZN => n36569);
   U1320 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_28_port, B1 => 
                           n36783, B2 => REGISTERS_18_28_port, ZN => n36568);
   U1321 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_28_port, B1 => 
                           n36785, B2 => REGISTERS_31_28_port, ZN => n36567);
   U1322 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_28_port, B1 => 
                           n36787, B2 => REGISTERS_8_28_port, ZN => n36566);
   U1323 : NAND4_X1 port map( A1 => n36569, A2 => n36568, A3 => n36567, A4 => 
                           n36566, ZN => n36575);
   U1324 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_28_port, B1 => 
                           n36793, B2 => REGISTERS_29_28_port, ZN => n36573);
   U1325 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_28_port, B1 => 
                           n36795, B2 => REGISTERS_16_28_port, ZN => n36572);
   U1326 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_28_port, B1 => 
                           n36797, B2 => REGISTERS_24_28_port, ZN => n36571);
   U1327 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_28_port, B1 => 
                           n36799, B2 => REGISTERS_15_28_port, ZN => n36570);
   U1328 : NAND4_X1 port map( A1 => n36573, A2 => n36572, A3 => n36571, A4 => 
                           n36570, ZN => n36574);
   U1329 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_29_port, B1 => 
                           n36758, B2 => REGISTERS_22_29_port, ZN => n36581);
   U1330 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_29_port, B1 => 
                           n36760, B2 => REGISTERS_21_29_port, ZN => n36580);
   U1331 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_29_port, B1 => 
                           n36762, B2 => REGISTERS_23_29_port, ZN => n36579);
   U1332 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_29_port, ZN => 
                           n36578);
   U1333 : NAND4_X1 port map( A1 => n36581, A2 => n36580, A3 => n36579, A4 => 
                           n36578, ZN => n36597);
   U1334 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_29_port, B1 => 
                           n36769, B2 => REGISTERS_13_29_port, ZN => n36585);
   U1335 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_29_port, B1 => 
                           n36277, B2 => REGISTERS_4_29_port, ZN => n36584);
   U1336 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_29_port, B1 => 
                           n36773, B2 => REGISTERS_28_29_port, ZN => n36583);
   U1337 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_29_port, B1 => 
                           n36775, B2 => REGISTERS_7_29_port, ZN => n36582);
   U1338 : NAND4_X1 port map( A1 => n36585, A2 => n36584, A3 => n36583, A4 => 
                           n36582, ZN => n36596);
   U1339 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_29_port, B1 => 
                           n36781, B2 => REGISTERS_9_29_port, ZN => n36589);
   U1340 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_29_port, B1 => 
                           n36783, B2 => REGISTERS_18_29_port, ZN => n36588);
   U1341 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_29_port, B1 => 
                           n36785, B2 => REGISTERS_31_29_port, ZN => n36587);
   U1342 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_29_port, B1 => 
                           n36787, B2 => REGISTERS_8_29_port, ZN => n36586);
   U1343 : NAND4_X1 port map( A1 => n36589, A2 => n36588, A3 => n36587, A4 => 
                           n36586, ZN => n36595);
   U1344 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_29_port, B1 => 
                           n36793, B2 => REGISTERS_29_29_port, ZN => n36593);
   U1345 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_29_port, B1 => 
                           n36795, B2 => REGISTERS_16_29_port, ZN => n36592);
   U1346 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_29_port, B1 => 
                           n36797, B2 => REGISTERS_24_29_port, ZN => n36591);
   U1347 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_29_port, B1 => 
                           n36799, B2 => REGISTERS_15_29_port, ZN => n36590);
   U1348 : NAND4_X1 port map( A1 => n36593, A2 => n36592, A3 => n36591, A4 => 
                           n36590, ZN => n36594);
   U1349 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_2_port, B1 => 
                           n36758, B2 => REGISTERS_22_2_port, ZN => n36601);
   U1350 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_2_port, B1 => 
                           n36760, B2 => REGISTERS_21_2_port, ZN => n36600);
   U1351 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_2_port, B1 => 
                           n36762, B2 => REGISTERS_23_2_port, ZN => n36599);
   U1352 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_2_port, ZN => 
                           n36598);
   U1353 : NAND4_X1 port map( A1 => n36601, A2 => n36600, A3 => n36599, A4 => 
                           n36598, ZN => n36617);
   U1354 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_2_port, B1 => 
                           n36769, B2 => REGISTERS_13_2_port, ZN => n36605);
   U1355 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_2_port, B1 => 
                           n36277, B2 => REGISTERS_4_2_port, ZN => n36604);
   U1356 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_2_port, B1 => 
                           n36773, B2 => REGISTERS_28_2_port, ZN => n36603);
   U1357 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_2_port, B1 => 
                           n36775, B2 => REGISTERS_7_2_port, ZN => n36602);
   U1358 : NAND4_X1 port map( A1 => n36605, A2 => n36604, A3 => n36603, A4 => 
                           n36602, ZN => n36616);
   U1359 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_2_port, B1 => 
                           n36781, B2 => REGISTERS_9_2_port, ZN => n36609);
   U1360 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_2_port, B1 => 
                           n36783, B2 => REGISTERS_18_2_port, ZN => n36608);
   U1361 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_2_port, B1 => 
                           n36785, B2 => REGISTERS_31_2_port, ZN => n36607);
   U1362 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_2_port, B1 => 
                           n36787, B2 => REGISTERS_8_2_port, ZN => n36606);
   U1363 : NAND4_X1 port map( A1 => n36609, A2 => n36608, A3 => n36607, A4 => 
                           n36606, ZN => n36615);
   U1364 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_2_port, B1 => 
                           n36793, B2 => REGISTERS_29_2_port, ZN => n36613);
   U1365 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_2_port, B1 => 
                           n36795, B2 => REGISTERS_16_2_port, ZN => n36612);
   U1366 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_2_port, B1 => 
                           n36797, B2 => REGISTERS_24_2_port, ZN => n36611);
   U1367 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_2_port, B1 => 
                           n36799, B2 => REGISTERS_15_2_port, ZN => n36610);
   U1368 : NAND4_X1 port map( A1 => n36613, A2 => n36612, A3 => n36611, A4 => 
                           n36610, ZN => n36614);
   U1369 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_30_port, B1 => 
                           n36758, B2 => REGISTERS_22_30_port, ZN => n36621);
   U1370 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_30_port, B1 => 
                           n36760, B2 => REGISTERS_21_30_port, ZN => n36620);
   U1371 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_30_port, B1 => 
                           n36272, B2 => REGISTERS_23_30_port, ZN => n36619);
   U1372 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_30_port, ZN => 
                           n36618);
   U1373 : NAND4_X1 port map( A1 => n36621, A2 => n36620, A3 => n36619, A4 => 
                           n36618, ZN => n36637);
   U1374 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_30_port, B1 => 
                           n36769, B2 => REGISTERS_13_30_port, ZN => n36625);
   U1375 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_30_port, B1 => 
                           n36771, B2 => REGISTERS_4_30_port, ZN => n36624);
   U1376 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_30_port, B1 => 
                           n36773, B2 => REGISTERS_28_30_port, ZN => n36623);
   U1377 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_30_port, B1 => 
                           n36775, B2 => REGISTERS_7_30_port, ZN => n36622);
   U1378 : NAND4_X1 port map( A1 => n36625, A2 => n36624, A3 => n36623, A4 => 
                           n36622, ZN => n36636);
   U1379 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_30_port, B1 => 
                           n36781, B2 => REGISTERS_9_30_port, ZN => n36629);
   U1380 : AOI22_X1 port map( A1 => n36784, A2 => REGISTERS_2_30_port, B1 => 
                           n36783, B2 => REGISTERS_18_30_port, ZN => n36628);
   U1381 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_30_port, B1 => 
                           n36785, B2 => REGISTERS_31_30_port, ZN => n36627);
   U1382 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_30_port, B1 => 
                           n36787, B2 => REGISTERS_8_30_port, ZN => n36626);
   U1383 : NAND4_X1 port map( A1 => n36629, A2 => n36628, A3 => n36627, A4 => 
                           n36626, ZN => n36635);
   U1384 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_30_port, B1 => 
                           n36793, B2 => REGISTERS_29_30_port, ZN => n36633);
   U1385 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_30_port, B1 => 
                           n36795, B2 => REGISTERS_16_30_port, ZN => n36632);
   U1386 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_30_port, B1 => 
                           n36797, B2 => REGISTERS_24_30_port, ZN => n36631);
   U1387 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_30_port, B1 => 
                           n36799, B2 => REGISTERS_15_30_port, ZN => n36630);
   U1388 : NAND4_X1 port map( A1 => n36633, A2 => n36632, A3 => n36631, A4 => 
                           n36630, ZN => n36634);
   U1389 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_3_port, B1 => 
                           n36758, B2 => REGISTERS_22_3_port, ZN => n36641);
   U1390 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_3_port, B1 => 
                           n36760, B2 => REGISTERS_21_3_port, ZN => n36640);
   U1391 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_3_port, B1 => 
                           n36762, B2 => REGISTERS_23_3_port, ZN => n36639);
   U1392 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_3_port, ZN => 
                           n36638);
   U1393 : NAND4_X1 port map( A1 => n36641, A2 => n36640, A3 => n36639, A4 => 
                           n36638, ZN => n36657);
   U1394 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_3_port, B1 => 
                           n36769, B2 => REGISTERS_13_3_port, ZN => n36645);
   U1395 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_3_port, B1 => 
                           n36771, B2 => REGISTERS_4_3_port, ZN => n36644);
   U1396 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_3_port, B1 => 
                           n36773, B2 => REGISTERS_28_3_port, ZN => n36643);
   U1397 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_3_port, B1 => 
                           n36775, B2 => REGISTERS_7_3_port, ZN => n36642);
   U1398 : NAND4_X1 port map( A1 => n36645, A2 => n36644, A3 => n36643, A4 => 
                           n36642, ZN => n36656);
   U1399 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_3_port, B1 => 
                           n36781, B2 => REGISTERS_9_3_port, ZN => n36649);
   U1400 : AOI22_X1 port map( A1 => n36784, A2 => REGISTERS_2_3_port, B1 => 
                           n36783, B2 => REGISTERS_18_3_port, ZN => n36648);
   U1401 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_3_port, B1 => 
                           n36785, B2 => REGISTERS_31_3_port, ZN => n36647);
   U1402 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_3_port, B1 => 
                           n36787, B2 => REGISTERS_8_3_port, ZN => n36646);
   U1403 : NAND4_X1 port map( A1 => n36649, A2 => n36648, A3 => n36647, A4 => 
                           n36646, ZN => n36655);
   U1404 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_3_port, B1 => 
                           n36793, B2 => REGISTERS_29_3_port, ZN => n36653);
   U1405 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_3_port, B1 => 
                           n36795, B2 => REGISTERS_16_3_port, ZN => n36652);
   U1406 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_3_port, B1 => 
                           n36797, B2 => REGISTERS_24_3_port, ZN => n36651);
   U1407 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_3_port, B1 => 
                           n36799, B2 => REGISTERS_15_3_port, ZN => n36650);
   U1408 : NAND4_X1 port map( A1 => n36653, A2 => n36652, A3 => n36651, A4 => 
                           n36650, ZN => n36654);
   U1409 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_4_port, B1 => 
                           n36758, B2 => REGISTERS_22_4_port, ZN => n36661);
   U1410 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_4_port, B1 => 
                           n36760, B2 => REGISTERS_21_4_port, ZN => n36660);
   U1411 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_4_port, B1 => 
                           n36762, B2 => REGISTERS_23_4_port, ZN => n36659);
   U1412 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_4_port, ZN => 
                           n36658);
   U1413 : NAND4_X1 port map( A1 => n36661, A2 => n36660, A3 => n36659, A4 => 
                           n36658, ZN => n36677);
   U1414 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_4_port, B1 => 
                           n36769, B2 => REGISTERS_13_4_port, ZN => n36665);
   U1415 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_4_port, B1 => 
                           n36771, B2 => REGISTERS_4_4_port, ZN => n36664);
   U1416 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_4_port, B1 => 
                           n36773, B2 => REGISTERS_28_4_port, ZN => n36663);
   U1417 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_4_port, B1 => 
                           n36775, B2 => REGISTERS_7_4_port, ZN => n36662);
   U1418 : NAND4_X1 port map( A1 => n36665, A2 => n36664, A3 => n36663, A4 => 
                           n36662, ZN => n36676);
   U1419 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_4_port, B1 => 
                           n36781, B2 => REGISTERS_9_4_port, ZN => n36669);
   U1420 : AOI22_X1 port map( A1 => n36784, A2 => REGISTERS_2_4_port, B1 => 
                           n36783, B2 => REGISTERS_18_4_port, ZN => n36668);
   U1421 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_4_port, B1 => 
                           n36785, B2 => REGISTERS_31_4_port, ZN => n36667);
   U1422 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_4_port, B1 => 
                           n36787, B2 => REGISTERS_8_4_port, ZN => n36666);
   U1423 : NAND4_X1 port map( A1 => n36669, A2 => n36668, A3 => n36667, A4 => 
                           n36666, ZN => n36675);
   U1424 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_4_port, B1 => 
                           n36793, B2 => REGISTERS_29_4_port, ZN => n36673);
   U1425 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_4_port, B1 => 
                           n36795, B2 => REGISTERS_16_4_port, ZN => n36672);
   U1426 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_4_port, B1 => 
                           n36797, B2 => REGISTERS_24_4_port, ZN => n36671);
   U1427 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_4_port, B1 => 
                           n36799, B2 => REGISTERS_15_4_port, ZN => n36670);
   U1428 : NAND4_X1 port map( A1 => n36673, A2 => n36672, A3 => n36671, A4 => 
                           n36670, ZN => n36674);
   U1429 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_5_port, B1 => 
                           n36758, B2 => REGISTERS_22_5_port, ZN => n36681);
   U1430 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_5_port, B1 => 
                           n36760, B2 => REGISTERS_21_5_port, ZN => n36680);
   U1431 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_5_port, B1 => 
                           n36762, B2 => REGISTERS_23_5_port, ZN => n36679);
   U1432 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_5_port, ZN => 
                           n36678);
   U1433 : NAND4_X1 port map( A1 => n36681, A2 => n36680, A3 => n36679, A4 => 
                           n36678, ZN => n36697);
   U1434 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_5_port, B1 => 
                           n36769, B2 => REGISTERS_13_5_port, ZN => n36685);
   U1435 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_5_port, B1 => 
                           n36771, B2 => REGISTERS_4_5_port, ZN => n36684);
   U1436 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_5_port, B1 => 
                           n36773, B2 => REGISTERS_28_5_port, ZN => n36683);
   U1437 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_5_port, B1 => 
                           n36775, B2 => REGISTERS_7_5_port, ZN => n36682);
   U1438 : NAND4_X1 port map( A1 => n36685, A2 => n36684, A3 => n36683, A4 => 
                           n36682, ZN => n36696);
   U1439 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_5_port, B1 => 
                           n36781, B2 => REGISTERS_9_5_port, ZN => n36689);
   U1440 : AOI22_X1 port map( A1 => n36784, A2 => REGISTERS_2_5_port, B1 => 
                           n36783, B2 => REGISTERS_18_5_port, ZN => n36688);
   U1441 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_5_port, B1 => 
                           n36785, B2 => REGISTERS_31_5_port, ZN => n36687);
   U1442 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_5_port, B1 => 
                           n36787, B2 => REGISTERS_8_5_port, ZN => n36686);
   U1443 : NAND4_X1 port map( A1 => n36689, A2 => n36688, A3 => n36687, A4 => 
                           n36686, ZN => n36695);
   U1444 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_5_port, B1 => 
                           n36793, B2 => REGISTERS_29_5_port, ZN => n36693);
   U1445 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_5_port, B1 => 
                           n36795, B2 => REGISTERS_16_5_port, ZN => n36692);
   U1446 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_5_port, B1 => 
                           n36797, B2 => REGISTERS_24_5_port, ZN => n36691);
   U1447 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_5_port, B1 => 
                           n36799, B2 => REGISTERS_15_5_port, ZN => n36690);
   U1448 : NAND4_X1 port map( A1 => n36693, A2 => n36692, A3 => n36691, A4 => 
                           n36690, ZN => n36694);
   U1449 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_6_port, B1 => 
                           n36758, B2 => REGISTERS_22_6_port, ZN => n36701);
   U1450 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_6_port, B1 => 
                           n36760, B2 => REGISTERS_21_6_port, ZN => n36700);
   U1451 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_6_port, B1 => 
                           n36762, B2 => REGISTERS_23_6_port, ZN => n36699);
   U1452 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_6_port, ZN => 
                           n36698);
   U1453 : NAND4_X1 port map( A1 => n36701, A2 => n36700, A3 => n36699, A4 => 
                           n36698, ZN => n36717);
   U1454 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_6_port, B1 => 
                           n36769, B2 => REGISTERS_13_6_port, ZN => n36705);
   U1455 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_6_port, B1 => 
                           n36771, B2 => REGISTERS_4_6_port, ZN => n36704);
   U1456 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_6_port, B1 => 
                           n36773, B2 => REGISTERS_28_6_port, ZN => n36703);
   U1457 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_6_port, B1 => 
                           n36775, B2 => REGISTERS_7_6_port, ZN => n36702);
   U1458 : NAND4_X1 port map( A1 => n36705, A2 => n36704, A3 => n36703, A4 => 
                           n36702, ZN => n36716);
   U1459 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_6_port, B1 => 
                           n36781, B2 => REGISTERS_9_6_port, ZN => n36709);
   U1460 : AOI22_X1 port map( A1 => n36784, A2 => REGISTERS_2_6_port, B1 => 
                           n36783, B2 => REGISTERS_18_6_port, ZN => n36708);
   U1461 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_6_port, B1 => 
                           n36785, B2 => REGISTERS_31_6_port, ZN => n36707);
   U1462 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_6_port, B1 => 
                           n36787, B2 => REGISTERS_8_6_port, ZN => n36706);
   U1463 : NAND4_X1 port map( A1 => n36709, A2 => n36708, A3 => n36707, A4 => 
                           n36706, ZN => n36715);
   U1464 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_6_port, B1 => 
                           n36793, B2 => REGISTERS_29_6_port, ZN => n36713);
   U1465 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_6_port, B1 => 
                           n36795, B2 => REGISTERS_16_6_port, ZN => n36712);
   U1466 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_6_port, B1 => 
                           n36797, B2 => REGISTERS_24_6_port, ZN => n36711);
   U1467 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_6_port, B1 => 
                           n36799, B2 => REGISTERS_15_6_port, ZN => n36710);
   U1468 : NAND4_X1 port map( A1 => n36713, A2 => n36712, A3 => n36711, A4 => 
                           n36710, ZN => n36714);
   U1469 : AOI22_X1 port map( A1 => n36269, A2 => REGISTERS_5_7_port, B1 => 
                           n36268, B2 => REGISTERS_22_7_port, ZN => n36721);
   U1470 : AOI22_X1 port map( A1 => n36271, A2 => REGISTERS_25_7_port, B1 => 
                           n36270, B2 => REGISTERS_21_7_port, ZN => n36720);
   U1471 : AOI22_X1 port map( A1 => n36273, A2 => REGISTERS_17_7_port, B1 => 
                           n36272, B2 => REGISTERS_23_7_port, ZN => n36719);
   U1472 : NAND2_X1 port map( A1 => n36764, A2 => REGISTERS_19_7_port, ZN => 
                           n36718);
   U1473 : NAND4_X1 port map( A1 => n36721, A2 => n36720, A3 => n36719, A4 => 
                           n36718, ZN => n36737);
   U1474 : AOI22_X1 port map( A1 => n36276, A2 => REGISTERS_14_7_port, B1 => 
                           n36275, B2 => REGISTERS_13_7_port, ZN => n36725);
   U1475 : AOI22_X1 port map( A1 => n36278, A2 => REGISTERS_27_7_port, B1 => 
                           n36277, B2 => REGISTERS_4_7_port, ZN => n36724);
   U1476 : AOI22_X1 port map( A1 => n36280, A2 => REGISTERS_6_7_port, B1 => 
                           n36279, B2 => REGISTERS_28_7_port, ZN => n36723);
   U1477 : AOI22_X1 port map( A1 => n36282, A2 => REGISTERS_26_7_port, B1 => 
                           n36281, B2 => REGISTERS_7_7_port, ZN => n36722);
   U1478 : NAND4_X1 port map( A1 => n36725, A2 => n36724, A3 => n36723, A4 => 
                           n36722, ZN => n36736);
   U1479 : AOI22_X1 port map( A1 => n36284, A2 => REGISTERS_10_7_port, B1 => 
                           n36283, B2 => REGISTERS_9_7_port, ZN => n36729);
   U1480 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_7_port, B1 => 
                           n36285, B2 => REGISTERS_18_7_port, ZN => n36728);
   U1481 : AOI22_X1 port map( A1 => n36288, A2 => REGISTERS_3_7_port, B1 => 
                           n36287, B2 => REGISTERS_31_7_port, ZN => n36727);
   U1482 : AOI22_X1 port map( A1 => n36290, A2 => REGISTERS_30_7_port, B1 => 
                           n36289, B2 => REGISTERS_8_7_port, ZN => n36726);
   U1483 : NAND4_X1 port map( A1 => n36729, A2 => n36728, A3 => n36727, A4 => 
                           n36726, ZN => n36735);
   U1484 : AOI22_X1 port map( A1 => n36292, A2 => REGISTERS_11_7_port, B1 => 
                           n36291, B2 => REGISTERS_29_7_port, ZN => n36733);
   U1485 : AOI22_X1 port map( A1 => n36294, A2 => REGISTERS_1_7_port, B1 => 
                           n36293, B2 => REGISTERS_16_7_port, ZN => n36732);
   U1486 : AOI22_X1 port map( A1 => n36296, A2 => REGISTERS_12_7_port, B1 => 
                           n36295, B2 => REGISTERS_24_7_port, ZN => n36731);
   U1487 : AOI22_X1 port map( A1 => n36298, A2 => REGISTERS_20_7_port, B1 => 
                           n36297, B2 => REGISTERS_15_7_port, ZN => n36730);
   U1488 : NAND4_X1 port map( A1 => n36733, A2 => n36732, A3 => n36731, A4 => 
                           n36730, ZN => n36734);
   U1489 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_8_port, B1 => 
                           n36268, B2 => REGISTERS_22_8_port, ZN => n36741);
   U1490 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_8_port, B1 => 
                           n36760, B2 => REGISTERS_21_8_port, ZN => n36740);
   U1491 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_8_port, B1 => 
                           n36762, B2 => REGISTERS_23_8_port, ZN => n36739);
   U1492 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_8_port, ZN => 
                           n36738);
   U1493 : NAND4_X1 port map( A1 => n36741, A2 => n36740, A3 => n36739, A4 => 
                           n36738, ZN => n36757);
   U1494 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_8_port, B1 => 
                           n36769, B2 => REGISTERS_13_8_port, ZN => n36745);
   U1495 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_8_port, B1 => 
                           n36277, B2 => REGISTERS_4_8_port, ZN => n36744);
   U1496 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_8_port, B1 => 
                           n36773, B2 => REGISTERS_28_8_port, ZN => n36743);
   U1497 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_8_port, B1 => 
                           n36775, B2 => REGISTERS_7_8_port, ZN => n36742);
   U1498 : NAND4_X1 port map( A1 => n36745, A2 => n36744, A3 => n36743, A4 => 
                           n36742, ZN => n36756);
   U1499 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_8_port, B1 => 
                           n36781, B2 => REGISTERS_9_8_port, ZN => n36749);
   U1500 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_8_port, B1 => 
                           n36783, B2 => REGISTERS_18_8_port, ZN => n36748);
   U1501 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_8_port, B1 => 
                           n36785, B2 => REGISTERS_31_8_port, ZN => n36747);
   U1502 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_8_port, B1 => 
                           n36787, B2 => REGISTERS_8_8_port, ZN => n36746);
   U1503 : NAND4_X1 port map( A1 => n36749, A2 => n36748, A3 => n36747, A4 => 
                           n36746, ZN => n36755);
   U1504 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_8_port, B1 => 
                           n36793, B2 => REGISTERS_29_8_port, ZN => n36753);
   U1505 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_8_port, B1 => 
                           n36795, B2 => REGISTERS_16_8_port, ZN => n36752);
   U1506 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_8_port, B1 => 
                           n36797, B2 => REGISTERS_24_8_port, ZN => n36751);
   U1507 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_8_port, B1 => 
                           n36799, B2 => REGISTERS_15_8_port, ZN => n36750);
   U1508 : NAND4_X1 port map( A1 => n36753, A2 => n36752, A3 => n36751, A4 => 
                           n36750, ZN => n36754);
   U1509 : AOI22_X1 port map( A1 => n36759, A2 => REGISTERS_5_9_port, B1 => 
                           n36758, B2 => REGISTERS_22_9_port, ZN => n36768);
   U1510 : AOI22_X1 port map( A1 => n36761, A2 => REGISTERS_25_9_port, B1 => 
                           n36760, B2 => REGISTERS_21_9_port, ZN => n36767);
   U1511 : AOI22_X1 port map( A1 => n36763, A2 => REGISTERS_17_9_port, B1 => 
                           n36762, B2 => REGISTERS_23_9_port, ZN => n36766);
   U1512 : NAND2_X1 port map( A1 => n36274, A2 => REGISTERS_19_9_port, ZN => 
                           n36765);
   U1513 : NAND4_X1 port map( A1 => n36768, A2 => n36767, A3 => n36766, A4 => 
                           n36765, ZN => n36808);
   U1514 : AOI22_X1 port map( A1 => n36770, A2 => REGISTERS_14_9_port, B1 => 
                           n36769, B2 => REGISTERS_13_9_port, ZN => n36780);
   U1515 : AOI22_X1 port map( A1 => n36772, A2 => REGISTERS_27_9_port, B1 => 
                           n36277, B2 => REGISTERS_4_9_port, ZN => n36779);
   U1516 : AOI22_X1 port map( A1 => n36774, A2 => REGISTERS_6_9_port, B1 => 
                           n36773, B2 => REGISTERS_28_9_port, ZN => n36778);
   U1517 : AOI22_X1 port map( A1 => n36776, A2 => REGISTERS_26_9_port, B1 => 
                           n36775, B2 => REGISTERS_7_9_port, ZN => n36777);
   U1518 : NAND4_X1 port map( A1 => n36780, A2 => n36779, A3 => n36778, A4 => 
                           n36777, ZN => n36807);
   U1519 : AOI22_X1 port map( A1 => n36782, A2 => REGISTERS_10_9_port, B1 => 
                           n36781, B2 => REGISTERS_9_9_port, ZN => n36792);
   U1520 : AOI22_X1 port map( A1 => n36286, A2 => REGISTERS_2_9_port, B1 => 
                           n36285, B2 => REGISTERS_18_9_port, ZN => n36791);
   U1521 : AOI22_X1 port map( A1 => n36786, A2 => REGISTERS_3_9_port, B1 => 
                           n36287, B2 => REGISTERS_31_9_port, ZN => n36790);
   U1522 : AOI22_X1 port map( A1 => n36788, A2 => REGISTERS_30_9_port, B1 => 
                           n36787, B2 => REGISTERS_8_9_port, ZN => n36789);
   U1523 : NAND4_X1 port map( A1 => n36792, A2 => n36791, A3 => n36790, A4 => 
                           n36789, ZN => n36806);
   U1524 : AOI22_X1 port map( A1 => n36794, A2 => REGISTERS_11_9_port, B1 => 
                           n36793, B2 => REGISTERS_29_9_port, ZN => n36804);
   U1525 : AOI22_X1 port map( A1 => n36796, A2 => REGISTERS_1_9_port, B1 => 
                           n36795, B2 => REGISTERS_16_9_port, ZN => n36803);
   U1526 : AOI22_X1 port map( A1 => n36798, A2 => REGISTERS_12_9_port, B1 => 
                           n36797, B2 => REGISTERS_24_9_port, ZN => n36802);
   U1527 : AOI22_X1 port map( A1 => n36800, A2 => REGISTERS_20_9_port, B1 => 
                           n36799, B2 => REGISTERS_15_9_port, ZN => n36801);
   U1528 : NAND4_X1 port map( A1 => n36804, A2 => n36803, A3 => n36802, A4 => 
                           n36801, ZN => n36805);
   U1529 : NAND3_X1 port map( A1 => ADD_RDB(0), A2 => ADD_RDB(4), A3 => n36810,
                           ZN => n36816);
   U1530 : INV_X1 port map( A => ADD_RDB(1), ZN => n36820);
   U1531 : NAND3_X1 port map( A1 => ADD_RDB(2), A2 => RESET, A3 => n36820, ZN 
                           => n36827);
   U1532 : NOR2_X1 port map( A1 => n36816, A2 => n36827, ZN => n36829);
   U1533 : INV_X1 port map( A => ADD_RDB(2), ZN => n36814);
   U1534 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDB(1), A3 => n36814, ZN 
                           => n36821);
   U1535 : INV_X1 port map( A => ADD_RDB(0), ZN => n36809);
   U1536 : NAND3_X1 port map( A1 => ADD_RDB(3), A2 => ADD_RDB(4), A3 => n36809,
                           ZN => n36813);
   U1537 : NOR2_X1 port map( A1 => n36821, A2 => n36813, ZN => n36828);
   U1538 : INV_X1 port map( A => ADD_RDB(4), ZN => n36817);
   U1539 : NAND3_X1 port map( A1 => ADD_RDB(0), A2 => n36810, A3 => n36817, ZN 
                           => n36815);
   U1540 : NAND3_X1 port map( A1 => RESET, A2 => ADD_RDB(2), A3 => ADD_RDB(1), 
                           ZN => n36823);
   U1541 : NOR2_X1 port map( A1 => n36815, A2 => n36823, ZN => n36831);
   U1542 : NAND3_X1 port map( A1 => RESET, A2 => n36814, A3 => n36820, ZN => 
                           n36825);
   U1543 : NOR2_X1 port map( A1 => n36815, A2 => n36825, ZN => n36830);
   U1544 : NOR2_X1 port map( A1 => n36827, A2 => n36815, ZN => n36833);
   U1545 : NAND3_X1 port map( A1 => ADD_RDB(4), A2 => n36810, A3 => n36809, ZN 
                           => n36818);
   U1546 : NOR2_X1 port map( A1 => n36818, A2 => n36827, ZN => n36832);
   U1547 : NOR2_X1 port map( A1 => n36821, A2 => n36818, ZN => n36834);
   U1548 : NOR2_X1 port map( A1 => n36821, A2 => n36816, ZN => n36836);
   U1549 : NOR2_X1 port map( A1 => n36813, A2 => n36827, ZN => n36835);
   U1550 : NOR2_X1 port map( A1 => n36816, A2 => n36823, ZN => n36838);
   U1551 : NAND2_X1 port map( A1 => ADD_RDB(2), A2 => ADD_RDB(1), ZN => n36811)
                           ;
   U1552 : NOR2_X1 port map( A1 => ADD_RDB(0), A2 => ADD_RDB(4), ZN => n36812);
   U1553 : NAND3_X1 port map( A1 => RESET, A2 => n36812, A3 => n36810, ZN => 
                           n36819);
   U1554 : NOR2_X1 port map( A1 => n36811, A2 => n36819, ZN => n36837);
   U1555 : NAND2_X1 port map( A1 => ADD_RDB(3), A2 => n36812, ZN => n36824);
   U1556 : NOR2_X1 port map( A1 => n36821, A2 => n36824, ZN => n36840);
   U1557 : NOR2_X1 port map( A1 => n36813, A2 => n36825, ZN => n36839);
   U1558 : NAND3_X1 port map( A1 => ADD_RDB(3), A2 => ADD_RDB(0), A3 => 
                           ADD_RDB(4), ZN => n36826);
   U1559 : NOR2_X1 port map( A1 => n36821, A2 => n36826, ZN => n36842);
   U1560 : NOR2_X1 port map( A1 => n36827, A2 => n36824, ZN => n36841);
   U1561 : NOR2_X1 port map( A1 => n36823, A2 => n36824, ZN => n36844);
   U1562 : NOR2_X1 port map( A1 => n36813, A2 => n36823, ZN => n36843);
   U1563 : NOR3_X1 port map( A1 => ADD_RDB(1), A2 => n36814, A3 => n36819, ZN 
                           => n36846);
   U1564 : NOR2_X1 port map( A1 => n36821, A2 => n36815, ZN => n36845);
   U1565 : NOR2_X1 port map( A1 => n36818, A2 => n36823, ZN => n36848);
   U1566 : NOR2_X1 port map( A1 => n36816, A2 => n36825, ZN => n36847);
   U1567 : NAND3_X1 port map( A1 => ADD_RDB(0), A2 => ADD_RDB(3), A3 => n36817,
                           ZN => n36822);
   U1568 : NOR2_X1 port map( A1 => n36825, A2 => n36822, ZN => n36850);
   U1569 : NOR2_X1 port map( A1 => n36823, A2 => n36822, ZN => n36849);
   U1570 : NOR2_X1 port map( A1 => n36825, A2 => n36826, ZN => n36852);
   U1571 : NOR2_X1 port map( A1 => n36818, A2 => n36825, ZN => n36851);
   U1572 : NOR3_X1 port map( A1 => ADD_RDB(2), A2 => n36820, A3 => n36819, ZN 
                           => n36854);
   U1573 : NOR2_X1 port map( A1 => n36821, A2 => n36822, ZN => n36853);
   U1574 : NOR2_X1 port map( A1 => n36827, A2 => n36822, ZN => n36856);
   U1575 : NOR2_X1 port map( A1 => n36825, A2 => n36824, ZN => n36858);
   U1576 : NOR2_X1 port map( A1 => n36827, A2 => n36826, ZN => n36857);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_syn.all;

entity DLX_syn is

   port( Clk, Rst : in std_logic;  IRAM_DATA_OUT, DRAM_DATA_OUT : in 
         std_logic_vector (31 downto 0);  DRAM_DATA_IN : out std_logic_vector 
         (31 downto 0);  DRAM_ADDRESS : out std_logic_vector (11 downto 0);  
         DRAM_ENABLE, DRAM_RW : out std_logic;  DRAM_SEL : out std_logic_vector
         (2 downto 0);  IRAM_ADDRESS : out std_logic_vector (7 downto 0));

end DLX_syn;

architecture SYN_structural of DLX_syn is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X4
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component branch_predictor
      port( RST : in std_logic;  PC_IN, PC_FAIL, IR_IN : in std_logic_vector 
            (31 downto 0);  IR_FAIL : in std_logic_vector (15 downto 0);  
            WRONG_PRE, RIGHT_PRE : in std_logic;  NPC_OUT, LINK_ADD : out 
            std_logic_vector (31 downto 0);  SEL, TAKEN : out std_logic);
   end component;
   
   component register_file_N32_addBit5
      port( RESET, RE, WE : in std_logic;  ADD_WR, ADD_RDA, ADD_RDB : in 
            std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
            downto 0);  OUTA, OUTB : out std_logic_vector (31 downto 0));
   end component;
   
   signal DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, IR_CU_31, IR_CU_28, IR_CU_27, 
      IR_CU_26, IR_CU_9_port, IR_CU_8_port, IR_CU_7_port, IR_CU_6_port, 
      IR_CU_5_port, IR_CU_4_port, IR_CU_1_port, IR_CU_0_port, BR_EN_i, 
      ALU_OPCODE_i_3_port, ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, 
      ALU_OPCODE_i_0_port, WB_MUX_SEL_i_1_port, RF_WE_i, 
      CU_I_aluOpcode_i_0_port, CU_I_aluOpcode_i_1_port, CU_I_aluOpcode_i_2_port
      , CU_I_aluOpcode_i_3_port, CU_I_aluOpcode_i_4_port, CU_I_cw2_1_port, 
      CU_I_cw_0_port, CU_I_cw_1_port, CU_I_cw_3_port, CU_I_cw_4_port, 
      CU_I_cw_6_port, CU_I_cw_7_port, CU_I_cw_10_port, DataP_LMD_out_0_port, 
      DataP_LMD_out_1_port, DataP_LMD_out_2_port, DataP_LMD_out_3_port, 
      DataP_LMD_out_4_port, DataP_LMD_out_5_port, DataP_LMD_out_6_port, 
      DataP_LMD_out_7_port, DataP_LMD_out_8_port, DataP_LMD_out_9_port, 
      DataP_LMD_out_10_port, DataP_LMD_out_11_port, DataP_LMD_out_12_port, 
      DataP_LMD_out_13_port, DataP_LMD_out_14_port, DataP_LMD_out_15_port, 
      DataP_LMD_out_16_port, DataP_LMD_out_17_port, DataP_LMD_out_18_port, 
      DataP_LMD_out_19_port, DataP_LMD_out_20_port, DataP_LMD_out_21_port, 
      DataP_LMD_out_22_port, DataP_LMD_out_23_port, DataP_LMD_out_24_port, 
      DataP_LMD_out_25_port, DataP_LMD_out_26_port, DataP_LMD_out_27_port, 
      DataP_LMD_out_28_port, DataP_LMD_out_29_port, DataP_LMD_out_30_port, 
      DataP_LMD_out_31_port, DataP_link_addr_W_0_port, DataP_link_addr_W_1_port
      , DataP_link_addr_W_2_port, DataP_link_addr_W_3_port, 
      DataP_link_addr_W_4_port, DataP_link_addr_W_5_port, 
      DataP_link_addr_W_6_port, DataP_link_addr_W_7_port, 
      DataP_link_addr_W_8_port, DataP_link_addr_W_9_port, 
      DataP_link_addr_W_10_port, DataP_link_addr_W_11_port, 
      DataP_link_addr_W_12_port, DataP_link_addr_W_13_port, 
      DataP_link_addr_W_14_port, DataP_link_addr_W_15_port, 
      DataP_link_addr_W_16_port, DataP_link_addr_W_17_port, 
      DataP_link_addr_W_18_port, DataP_link_addr_W_19_port, 
      DataP_link_addr_W_20_port, DataP_link_addr_W_21_port, 
      DataP_link_addr_W_22_port, DataP_link_addr_W_23_port, 
      DataP_link_addr_W_24_port, DataP_link_addr_W_25_port, 
      DataP_link_addr_W_26_port, DataP_link_addr_W_27_port, 
      DataP_link_addr_W_28_port, DataP_link_addr_W_29_port, 
      DataP_link_addr_W_30_port, DataP_link_addr_W_31_port, 
      DataP_FWD_MUX_BR_S_0_port, DataP_FWD_MUX_BR_S_1_port, 
      DataP_alu_b_in_0_port, DataP_alu_b_in_1_port, DataP_alu_b_in_2_port, 
      DataP_alu_b_in_3_port, DataP_alu_b_in_6_port, DataP_alu_b_in_7_port, 
      DataP_alu_b_in_8_port, DataP_alu_b_in_9_port, DataP_alu_b_in_10_port, 
      DataP_alu_b_in_11_port, DataP_alu_b_in_12_port, DataP_alu_b_in_13_port, 
      DataP_alu_b_in_15_port, DataP_alu_b_in_16_port, DataP_alu_b_in_17_port, 
      DataP_alu_b_in_18_port, DataP_alu_b_in_19_port, DataP_alu_b_in_20_port, 
      DataP_alu_b_in_21_port, DataP_alu_b_in_22_port, DataP_alu_b_in_23_port, 
      DataP_alu_b_in_24_port, DataP_alu_b_in_26_port, DataP_alu_b_in_27_port, 
      DataP_alu_b_in_28_port, DataP_alu_b_in_29_port, DataP_alu_b_in_30_port, 
      DataP_alu_b_in_31_port, DataP_alu_a_in_0_port, DataP_alu_a_in_2_port, 
      DataP_alu_a_in_3_port, DataP_alu_a_in_4_port, DataP_alu_a_in_5_port, 
      DataP_alu_a_in_6_port, DataP_alu_a_in_7_port, DataP_alu_a_in_8_port, 
      DataP_alu_a_in_9_port, DataP_alu_a_in_10_port, DataP_alu_a_in_11_port, 
      DataP_alu_a_in_12_port, DataP_alu_a_in_13_port, DataP_alu_a_in_14_port, 
      DataP_alu_a_in_15_port, DataP_alu_a_in_16_port, DataP_alu_a_in_17_port, 
      DataP_alu_a_in_18_port, DataP_alu_a_in_19_port, DataP_alu_a_in_20_port, 
      DataP_alu_a_in_21_port, DataP_alu_a_in_22_port, DataP_alu_a_in_23_port, 
      DataP_alu_a_in_24_port, DataP_alu_a_in_25_port, DataP_alu_a_in_26_port, 
      DataP_alu_a_in_27_port, DataP_alu_a_in_28_port, DataP_alu_a_in_29_port, 
      DataP_alu_a_in_30_port, DataP_alu_a_in_31_port, DataP_alu_out_W_0_port, 
      DataP_alu_out_W_1_port, DataP_alu_out_W_2_port, DataP_alu_out_W_3_port, 
      DataP_alu_out_W_4_port, DataP_alu_out_W_5_port, DataP_alu_out_W_6_port, 
      DataP_alu_out_W_7_port, DataP_alu_out_W_8_port, DataP_alu_out_W_9_port, 
      DataP_alu_out_W_10_port, DataP_alu_out_W_11_port, DataP_alu_out_W_12_port
      , DataP_alu_out_W_13_port, DataP_alu_out_W_14_port, 
      DataP_alu_out_W_15_port, DataP_alu_out_W_16_port, DataP_alu_out_W_17_port
      , DataP_alu_out_W_18_port, DataP_alu_out_W_19_port, 
      DataP_alu_out_W_20_port, DataP_alu_out_W_21_port, DataP_alu_out_W_22_port
      , DataP_alu_out_W_23_port, DataP_alu_out_W_24_port, 
      DataP_alu_out_W_25_port, DataP_alu_out_W_26_port, DataP_alu_out_W_27_port
      , DataP_alu_out_W_28_port, DataP_alu_out_W_29_port, 
      DataP_alu_out_W_30_port, DataP_alu_out_W_31_port, DataP_alu_out_M_12_port
      , DataP_alu_out_M_13_port, DataP_alu_out_M_14_port, 
      DataP_alu_out_M_15_port, DataP_alu_out_M_16_port, DataP_alu_out_M_17_port
      , DataP_alu_out_M_18_port, DataP_alu_out_M_19_port, 
      DataP_alu_out_M_20_port, DataP_alu_out_M_21_port, DataP_alu_out_M_22_port
      , DataP_alu_out_M_23_port, DataP_alu_out_M_24_port, 
      DataP_alu_out_M_25_port, DataP_alu_out_M_26_port, DataP_alu_out_M_27_port
      , DataP_alu_out_M_28_port, DataP_alu_out_M_29_port, 
      DataP_alu_out_M_30_port, DataP_alu_out_M_31_port, DataP_opcode_W_0_port, 
      DataP_opcode_W_1_port, DataP_opcode_W_2_port, DataP_opcode_W_3_port, 
      DataP_opcode_W_4_port, DataP_opcode_W_5_port, DataP_opcode_M_0_port, 
      DataP_opcode_M_1_port, DataP_opcode_M_2_port, DataP_opcode_M_3_port, 
      DataP_opcode_M_4_port, DataP_dest_M_0_port, DataP_dest_M_1_port, 
      DataP_dest_M_2_port, DataP_dest_M_3_port, DataP_dest_M_4_port, DataP_pr_E
      , DataP_opcode_E_0_port, DataP_opcode_E_1_port, DataP_opcode_E_3_port, 
      DataP_opcode_E_4_port, DataP_Rs2_0_port, DataP_Rs2_1_port, 
      DataP_Rs2_2_port, DataP_Rs2_3_port, DataP_Rs2_4_port, DataP_Rs1_1_port, 
      DataP_Rs1_2_port, DataP_IMM_s_0_port, DataP_IMM_s_1_port, 
      DataP_IMM_s_2_port, DataP_IMM_s_3_port, DataP_IMM_s_4_port, 
      DataP_IMM_s_5_port, DataP_IMM_s_6_port, DataP_IMM_s_7_port, 
      DataP_IMM_s_8_port, DataP_IMM_s_9_port, DataP_IMM_s_10_port, 
      DataP_IMM_s_11_port, DataP_IMM_s_12_port, DataP_IMM_s_13_port, 
      DataP_IMM_s_14_port, DataP_IMM_s_15_port, DataP_IMM_s_16_port, 
      DataP_IMM_s_17_port, DataP_IMM_s_18_port, DataP_IMM_s_19_port, 
      DataP_IMM_s_20_port, DataP_IMM_s_21_port, DataP_IMM_s_22_port, 
      DataP_IMM_s_23_port, DataP_IMM_s_24_port, DataP_IMM_s_30_port, 
      DataP_B_s_0_port, DataP_B_s_1_port, DataP_B_s_2_port, DataP_B_s_3_port, 
      DataP_B_s_4_port, DataP_B_s_5_port, DataP_B_s_6_port, DataP_B_s_7_port, 
      DataP_B_s_8_port, DataP_B_s_9_port, DataP_B_s_10_port, DataP_B_s_11_port,
      DataP_B_s_12_port, DataP_B_s_13_port, DataP_B_s_14_port, 
      DataP_B_s_15_port, DataP_B_s_16_port, DataP_B_s_17_port, 
      DataP_B_s_18_port, DataP_B_s_19_port, DataP_B_s_20_port, 
      DataP_B_s_21_port, DataP_B_s_22_port, DataP_B_s_23_port, 
      DataP_B_s_24_port, DataP_B_s_25_port, DataP_B_s_26_port, 
      DataP_B_s_27_port, DataP_B_s_28_port, DataP_B_s_29_port, 
      DataP_B_s_30_port, DataP_B_s_31_port, DataP_A_s_0_port, DataP_A_s_1_port,
      DataP_A_s_2_port, DataP_A_s_3_port, DataP_A_s_4_port, DataP_A_s_5_port, 
      DataP_A_s_6_port, DataP_A_s_7_port, DataP_A_s_8_port, DataP_A_s_9_port, 
      DataP_A_s_10_port, DataP_A_s_11_port, DataP_A_s_12_port, 
      DataP_A_s_13_port, DataP_A_s_14_port, DataP_A_s_15_port, 
      DataP_A_s_16_port, DataP_A_s_17_port, DataP_A_s_18_port, 
      DataP_A_s_19_port, DataP_A_s_20_port, DataP_A_s_21_port, 
      DataP_A_s_22_port, DataP_A_s_23_port, DataP_A_s_24_port, 
      DataP_A_s_25_port, DataP_A_s_26_port, DataP_A_s_27_port, 
      DataP_A_s_28_port, DataP_A_s_29_port, DataP_A_s_30_port, 
      DataP_A_s_31_port, DataP_npc_E_9_port, DataP_imm_out_16_port, 
      DataP_imm_out_17_port, DataP_imm_out_18_port, DataP_imm_out_19_port, 
      DataP_imm_out_20_port, DataP_imm_out_21_port, DataP_imm_out_22_port, 
      DataP_imm_out_23_port, DataP_imm_out_24_port, DataP_imm_out_31_port, 
      DataP_b_out_0_port, DataP_b_out_1_port, DataP_b_out_2_port, 
      DataP_b_out_3_port, DataP_b_out_4_port, DataP_b_out_5_port, 
      DataP_b_out_6_port, DataP_b_out_7_port, DataP_b_out_8_port, 
      DataP_b_out_9_port, DataP_b_out_10_port, DataP_b_out_11_port, 
      DataP_b_out_12_port, DataP_b_out_13_port, DataP_b_out_14_port, 
      DataP_b_out_15_port, DataP_b_out_16_port, DataP_b_out_17_port, 
      DataP_b_out_18_port, DataP_b_out_19_port, DataP_b_out_20_port, 
      DataP_b_out_21_port, DataP_b_out_22_port, DataP_b_out_23_port, 
      DataP_b_out_24_port, DataP_b_out_25_port, DataP_b_out_26_port, 
      DataP_b_out_27_port, DataP_b_out_28_port, DataP_b_out_29_port, 
      DataP_b_out_30_port, DataP_b_out_31_port, DataP_a_out_0_port, 
      DataP_a_out_1_port, DataP_a_out_2_port, DataP_a_out_3_port, 
      DataP_a_out_4_port, DataP_a_out_5_port, DataP_a_out_6_port, 
      DataP_a_out_7_port, DataP_a_out_8_port, DataP_a_out_9_port, 
      DataP_a_out_10_port, DataP_a_out_11_port, DataP_a_out_12_port, 
      DataP_a_out_13_port, DataP_a_out_14_port, DataP_a_out_15_port, 
      DataP_a_out_16_port, DataP_a_out_17_port, DataP_a_out_18_port, 
      DataP_a_out_19_port, DataP_a_out_20_port, DataP_a_out_21_port, 
      DataP_a_out_22_port, DataP_a_out_23_port, DataP_a_out_24_port, 
      DataP_a_out_25_port, DataP_a_out_26_port, DataP_a_out_27_port, 
      DataP_a_out_28_port, DataP_a_out_29_port, DataP_a_out_30_port, 
      DataP_a_out_31_port, DataP_WB_0_port, DataP_WB_1_port, DataP_WB_2_port, 
      DataP_WB_3_port, DataP_WB_4_port, DataP_WB_5_port, DataP_WB_6_port, 
      DataP_WB_7_port, DataP_WB_8_port, DataP_WB_9_port, DataP_WB_10_port, 
      DataP_WB_11_port, DataP_WB_12_port, DataP_WB_13_port, DataP_WB_14_port, 
      DataP_WB_15_port, DataP_WB_16_port, DataP_WB_17_port, DataP_WB_18_port, 
      DataP_WB_19_port, DataP_WB_20_port, DataP_WB_21_port, DataP_WB_22_port, 
      DataP_WB_23_port, DataP_WB_24_port, DataP_WB_25_port, DataP_WB_26_port, 
      DataP_WB_27_port, DataP_WB_28_port, DataP_WB_29_port, DataP_WB_30_port, 
      DataP_WB_31_port, DataP_add_D_0_port, DataP_add_D_1_port, 
      DataP_add_D_2_port, DataP_add_D_3_port, DataP_add_D_4_port, 
      DataP_dest_D_0_port, DataP_dest_D_1_port, DataP_dest_D_2_port, 
      DataP_dest_D_3_port, DataP_dest_D_4_port, DataP_add_S2_0_port, 
      DataP_add_S2_1_port, DataP_add_S2_2_port, DataP_add_S2_3_port, 
      DataP_add_S2_4_port, DataP_pr_D, DataP_link_addr_D_0_port, 
      DataP_link_addr_D_1_port, DataP_link_addr_D_2_port, 
      DataP_link_addr_D_3_port, DataP_link_addr_D_4_port, 
      DataP_link_addr_D_5_port, DataP_link_addr_D_6_port, 
      DataP_link_addr_D_7_port, DataP_link_addr_D_8_port, 
      DataP_link_addr_D_9_port, DataP_link_addr_D_10_port, 
      DataP_link_addr_D_11_port, DataP_link_addr_D_12_port, 
      DataP_link_addr_D_13_port, DataP_link_addr_D_14_port, 
      DataP_link_addr_D_15_port, DataP_link_addr_D_16_port, 
      DataP_link_addr_D_17_port, DataP_link_addr_D_18_port, 
      DataP_link_addr_D_19_port, DataP_link_addr_D_20_port, 
      DataP_link_addr_D_21_port, DataP_link_addr_D_22_port, 
      DataP_link_addr_D_23_port, DataP_link_addr_D_24_port, 
      DataP_link_addr_D_25_port, DataP_link_addr_D_26_port, 
      DataP_link_addr_D_27_port, DataP_link_addr_D_28_port, 
      DataP_link_addr_D_29_port, DataP_link_addr_D_30_port, 
      DataP_link_addr_D_31_port, DataP_prediction, DataP_npc_mux_sel, 
      DataP_link_addr_F_0_port, DataP_link_addr_F_1_port, 
      DataP_link_addr_F_2_port, DataP_link_addr_F_3_port, 
      DataP_link_addr_F_4_port, DataP_link_addr_F_5_port, 
      DataP_link_addr_F_6_port, DataP_link_addr_F_7_port, 
      DataP_link_addr_F_8_port, DataP_link_addr_F_9_port, 
      DataP_link_addr_F_10_port, DataP_link_addr_F_11_port, 
      DataP_link_addr_F_12_port, DataP_link_addr_F_13_port, 
      DataP_link_addr_F_14_port, DataP_link_addr_F_15_port, 
      DataP_link_addr_F_16_port, DataP_link_addr_F_17_port, 
      DataP_link_addr_F_18_port, DataP_link_addr_F_19_port, 
      DataP_link_addr_F_20_port, DataP_link_addr_F_21_port, 
      DataP_link_addr_F_22_port, DataP_link_addr_F_23_port, 
      DataP_link_addr_F_24_port, DataP_link_addr_F_25_port, 
      DataP_link_addr_F_26_port, DataP_link_addr_F_27_port, 
      DataP_link_addr_F_28_port, DataP_link_addr_F_29_port, 
      DataP_link_addr_F_30_port, DataP_link_addr_F_31_port, 
      DataP_npc_pre_0_port, DataP_npc_pre_1_port, DataP_npc_pre_2_port, 
      DataP_npc_pre_3_port, DataP_npc_pre_4_port, DataP_npc_pre_5_port, 
      DataP_npc_pre_6_port, DataP_npc_pre_7_port, DataP_npc_pre_8_port, 
      DataP_npc_pre_9_port, DataP_npc_pre_10_port, DataP_npc_pre_11_port, 
      DataP_npc_pre_12_port, DataP_npc_pre_13_port, DataP_npc_pre_14_port, 
      DataP_npc_pre_15_port, DataP_npc_pre_16_port, DataP_npc_pre_17_port, 
      DataP_npc_pre_18_port, DataP_npc_pre_19_port, DataP_npc_pre_20_port, 
      DataP_npc_pre_21_port, DataP_npc_pre_22_port, DataP_npc_pre_23_port, 
      DataP_npc_pre_24_port, DataP_npc_pre_25_port, DataP_npc_pre_26_port, 
      DataP_npc_pre_27_port, DataP_npc_pre_28_port, DataP_npc_pre_29_port, 
      DataP_npc_pre_30_port, DataP_npc_pre_31_port, DataP_right_br, 
      DataP_wrong_br, DataP_npc_M_0_port, DataP_npc_M_1_port, 
      DataP_npc_M_2_port, DataP_npc_M_3_port, DataP_npc_M_4_port, 
      DataP_npc_M_5_port, DataP_npc_M_6_port, DataP_npc_M_7_port, 
      DataP_npc_M_8_port, DataP_npc_M_9_port, DataP_npc_M_10_port, 
      DataP_npc_M_11_port, DataP_npc_M_12_port, DataP_npc_M_13_port, 
      DataP_npc_M_14_port, DataP_npc_M_15_port, DataP_npc_M_16_port, 
      DataP_npc_M_17_port, DataP_npc_M_18_port, DataP_npc_M_19_port, 
      DataP_npc_M_20_port, DataP_npc_M_21_port, DataP_npc_M_22_port, 
      DataP_npc_M_23_port, DataP_npc_M_24_port, DataP_npc_M_25_port, 
      DataP_npc_M_26_port, DataP_npc_M_27_port, DataP_npc_M_28_port, 
      DataP_npc_M_29_port, DataP_npc_M_30_port, DataP_npc_M_31_port, 
      DataP_pc_out_0, DataP_pc_out_1, DataP_pc_out_10_port, 
      DataP_pc_out_11_port, DataP_pc_out_12_port, DataP_pc_out_13_port, 
      DataP_pc_out_14_port, DataP_pc_out_15_port, DataP_pc_out_16_port, 
      DataP_pc_out_17_port, DataP_pc_out_18_port, DataP_pc_out_19_port, 
      DataP_pc_out_20_port, DataP_pc_out_21_port, DataP_pc_out_22_port, 
      DataP_pc_out_23_port, DataP_pc_out_24_port, DataP_pc_out_25_port, 
      DataP_pc_out_26_port, DataP_pc_out_27_port, DataP_pc_out_28_port, 
      DataP_pc_out_29_port, DataP_pc_out_30_port, DataP_pc_out_31_port, 
      DataP_npc_0_port, DataP_npc_1_port, DataP_npc_2_port, DataP_npc_3_port, 
      DataP_npc_4_port, DataP_npc_5_port, DataP_npc_6_port, DataP_npc_7_port, 
      DataP_npc_8_port, DataP_npc_9_port, DataP_npc_10_port, DataP_npc_11_port,
      DataP_npc_12_port, DataP_npc_13_port, DataP_npc_14_port, 
      DataP_npc_15_port, DataP_npc_16_port, DataP_npc_17_port, 
      DataP_npc_18_port, DataP_npc_19_port, DataP_npc_20_port, 
      DataP_npc_21_port, DataP_npc_22_port, DataP_npc_23_port, 
      DataP_npc_24_port, DataP_npc_25_port, DataP_npc_26_port, 
      DataP_npc_27_port, DataP_npc_28_port, DataP_npc_29_port, 
      DataP_npc_30_port, DataP_npc_31_port, DataP_IR1_11_port, 
      DataP_IR1_12_port, DataP_IR1_13_port, DataP_IR1_14_port, 
      DataP_IR1_15_port, DataP_IR1_21_port, DataP_IR1_22_port, 
      DataP_IR1_23_port, DataP_IR1_24_port, DataP_IR1_25_port, DataP_PC_reg_N33
      , DataP_PC_reg_N32, DataP_PC_reg_N31, DataP_PC_reg_N30, DataP_PC_reg_N29,
      DataP_PC_reg_N28, DataP_PC_reg_N27, DataP_PC_reg_N26, DataP_PC_reg_N25, 
      DataP_PC_reg_N24, DataP_PC_reg_N23, DataP_PC_reg_N22, DataP_PC_reg_N21, 
      DataP_PC_reg_N20, DataP_PC_reg_N19, DataP_PC_reg_N18, DataP_PC_reg_N17, 
      DataP_PC_reg_N16, DataP_PC_reg_N15, DataP_PC_reg_N14, DataP_PC_reg_N13, 
      DataP_PC_reg_N12, DataP_PC_reg_N11, DataP_PC_reg_N10, DataP_PC_reg_N9, 
      DataP_PC_reg_N8, DataP_PC_reg_N7, DataP_PC_reg_N6, DataP_PC_reg_N5, 
      DataP_PC_reg_N4, DataP_PC_reg_N3, DataP_PC_reg_N2, DataP_NPC_add_N32, 
      DataP_NPC_add_N31, DataP_NPC_add_N30, DataP_NPC_add_N29, 
      DataP_NPC_add_N28, DataP_NPC_add_N27, DataP_NPC_add_N26, 
      DataP_NPC_add_N25, DataP_NPC_add_N24, DataP_NPC_add_N23, 
      DataP_NPC_add_N22, DataP_NPC_add_N21, DataP_NPC_add_N20, 
      DataP_NPC_add_N19, DataP_NPC_add_N18, DataP_NPC_add_N17, 
      DataP_NPC_add_N16, DataP_NPC_add_N15, DataP_NPC_add_N14, 
      DataP_NPC_add_N13, DataP_NPC_add_N12, DataP_NPC_add_N11, 
      DataP_NPC_add_N10, DataP_NPC_add_N9, DataP_NPC_add_N8, DataP_NPC_add_N7, 
      DataP_NPC_add_N6, DataP_NPC_add_N5, DataP_NPC_add_N4, DataP_NPC_add_N3, 
      DataP_NPC_add_N2, DataP_NPC_add_N1, DataP_NPC_add_N0, 
      DataP_FORWARDING_BR_N12, DataP_ALU_C_shifter_N108, 
      DataP_ALU_C_shifter_N107, DataP_ALU_C_shifter_N106, 
      DataP_ALU_C_shifter_N105, DataP_ALU_C_shifter_N104, 
      DataP_ALU_C_shifter_N103, DataP_ALU_C_shifter_N102, 
      DataP_ALU_C_shifter_N101, DataP_ALU_C_shifter_N100, 
      DataP_ALU_C_shifter_N99, DataP_ALU_C_shifter_N97, DataP_ALU_C_shifter_N96
      , DataP_ALU_C_shifter_N93, DataP_ALU_C_shifter_N84, 
      DataP_ALU_C_shifter_N83, DataP_ALU_C_shifter_N82, DataP_ALU_C_shifter_N81
      , DataP_ALU_C_shifter_N80, DataP_ALU_C_shifter_N79, 
      DataP_ALU_C_shifter_N78, DataP_ALU_C_shifter_N77, DataP_ALU_C_shifter_N76
      , DataP_ALU_C_shifter_N75, DataP_ALU_C_shifter_N74, 
      DataP_ALU_C_shifter_N73, DataP_ALU_C_shifter_N72, DataP_ALU_C_shifter_N71
      , DataP_ALU_C_shifter_N70, DataP_ALU_C_shifter_N69, 
      DataP_ALU_C_shifter_N67, DataP_ALU_C_shifter_N66, DataP_ALU_C_shifter_N65
      , DataP_ALU_C_shifter_N64, DataP_ALU_C_shifter_N61, 
      DataP_ALU_C_shifter_N59, DataP_ALU_C_shifter_N52, DataP_ALU_C_shifter_N51
      , DataP_ALU_C_shifter_N50, DataP_ALU_C_shifter_N49, 
      DataP_ALU_C_shifter_N47, DataP_ALU_C_shifter_N46, DataP_ALU_C_shifter_N45
      , DataP_ALU_C_shifter_N43, DataP_ALU_C_shifter_N42, 
      DataP_ALU_C_shifter_N41, DataP_ALU_C_shifter_N40, DataP_ALU_C_shifter_N39
      , DataP_ALU_C_shifter_N38, DataP_ALU_C_shifter_N37, 
      DataP_ALU_C_shifter_N36, DataP_ALU_C_shifter_N34, DataP_ALU_C_shifter_N33
      , DataP_ALU_C_shifter_N32, DataP_ALU_C_shifter_N29, 
      DataP_ALU_C_shifter_N20, DataP_ALU_C_shifter_N19, DataP_ALU_C_comp_N50, 
      DataP_ALU_C_comp_N24, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n294, n296, n297, n299, n300, n301, n303, n304, n308, n311, n313, n317, 
      n319, n322, n323, n326, n330, n332, n333, n337, n340, n341, n345, n350, 
      n353, n354, n355, n356, n357, n358, n399, n432, n443, n476, n477, n478, 
      n479, n480, n482, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n497, n504, n514, n515, n516, n520, n521, n523, n524, n528, 
      n529, n530, n536, n538, n540, n607, n1358, n1372, n1449, n1450, n1451, 
      n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, 
      n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, 
      n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, 
      n1546, sra_131_SH_4_port, lt_x_135_B_12_port, lt_x_135_B_5_port, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
      n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
      n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
      n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, 
      n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
      n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, 
      n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
      n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
      n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
      n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
      n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, 
      n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
      n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, 
      n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
      n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, 
      n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, 
      n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, 
      n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, 
      n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
      n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, 
      n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, 
      n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, 
      n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, 
      n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, 
      n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
      n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
      n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
      n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
      n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, 
      n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, 
      n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, 
      n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
      n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, 
      n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, 
      n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, 
      n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
      n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, 
      n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, 
      n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, 
      n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, 
      n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
      n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
      n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
      n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
      n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
      n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
      n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
      n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
      n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
      n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
      n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
      n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
      n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
      n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
      n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
      n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
      n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
      n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
      n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, 
      n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, 
      n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
      n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, 
      n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, 
      n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, 
      n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
      n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, 
      n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
      n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
      n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, 
      n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, 
      n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, 
      n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
      n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, 
      n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, 
      n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, 
      n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, 
      n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, 
      n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, 
      n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, 
      n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, 
      n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, 
      n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, 
      n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
      n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, 
      n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
      n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, 
      n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
      n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
      n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, 
      n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
      n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
      n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
      n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
      n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
      n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, 
      n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
      n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
      n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
      n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4220, n4221, n4222, n4223, n4224, n_1004, n_1005, n_1006, n_1007,
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358 : 
      std_logic;

begin
   DRAM_ADDRESS <= ( DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, 
      DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, 
      DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, 
      DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, 
      DRAM_ADDRESS_0_port );
   IRAM_ADDRESS <= ( IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   
   DataP_Reg_F : register_file_N32_addBit5 port map( RESET => Rst, RE => n1546,
                           WE => RF_WE_i, ADD_WR(4) => n1629, ADD_WR(3) => 
                           n2146, ADD_WR(2) => DataP_add_D_2_port, ADD_WR(1) =>
                           n2229, ADD_WR(0) => DataP_add_D_0_port, ADD_RDA(4) 
                           => n494, ADD_RDA(3) => n493, ADD_RDA(2) => n492, 
                           ADD_RDA(1) => n491, ADD_RDA(0) => n490, ADD_RDB(4) 
                           => DataP_add_S2_4_port, ADD_RDB(3) => 
                           DataP_add_S2_3_port, ADD_RDB(2) => 
                           DataP_add_S2_2_port, ADD_RDB(1) => 
                           DataP_add_S2_1_port, ADD_RDB(0) => 
                           DataP_add_S2_0_port, DATAIN(31) => DataP_WB_31_port,
                           DATAIN(30) => DataP_WB_30_port, DATAIN(29) => 
                           DataP_WB_29_port, DATAIN(28) => DataP_WB_28_port, 
                           DATAIN(27) => DataP_WB_27_port, DATAIN(26) => 
                           DataP_WB_26_port, DATAIN(25) => DataP_WB_25_port, 
                           DATAIN(24) => DataP_WB_24_port, DATAIN(23) => 
                           DataP_WB_23_port, DATAIN(22) => DataP_WB_22_port, 
                           DATAIN(21) => DataP_WB_21_port, DATAIN(20) => 
                           DataP_WB_20_port, DATAIN(19) => DataP_WB_19_port, 
                           DATAIN(18) => DataP_WB_18_port, DATAIN(17) => 
                           DataP_WB_17_port, DATAIN(16) => DataP_WB_16_port, 
                           DATAIN(15) => DataP_WB_15_port, DATAIN(14) => 
                           DataP_WB_14_port, DATAIN(13) => DataP_WB_13_port, 
                           DATAIN(12) => DataP_WB_12_port, DATAIN(11) => 
                           DataP_WB_11_port, DATAIN(10) => DataP_WB_10_port, 
                           DATAIN(9) => DataP_WB_9_port, DATAIN(8) => 
                           DataP_WB_8_port, DATAIN(7) => DataP_WB_7_port, 
                           DATAIN(6) => DataP_WB_6_port, DATAIN(5) => 
                           DataP_WB_5_port, DATAIN(4) => DataP_WB_4_port, 
                           DATAIN(3) => DataP_WB_3_port, DATAIN(2) => 
                           DataP_WB_2_port, DATAIN(1) => DataP_WB_1_port, 
                           DATAIN(0) => DataP_WB_0_port, OUTA(31) => 
                           DataP_a_out_31_port, OUTA(30) => DataP_a_out_30_port
                           , OUTA(29) => DataP_a_out_29_port, OUTA(28) => 
                           DataP_a_out_28_port, OUTA(27) => DataP_a_out_27_port
                           , OUTA(26) => DataP_a_out_26_port, OUTA(25) => 
                           DataP_a_out_25_port, OUTA(24) => DataP_a_out_24_port
                           , OUTA(23) => DataP_a_out_23_port, OUTA(22) => 
                           DataP_a_out_22_port, OUTA(21) => DataP_a_out_21_port
                           , OUTA(20) => DataP_a_out_20_port, OUTA(19) => 
                           DataP_a_out_19_port, OUTA(18) => DataP_a_out_18_port
                           , OUTA(17) => DataP_a_out_17_port, OUTA(16) => 
                           DataP_a_out_16_port, OUTA(15) => DataP_a_out_15_port
                           , OUTA(14) => DataP_a_out_14_port, OUTA(13) => 
                           DataP_a_out_13_port, OUTA(12) => DataP_a_out_12_port
                           , OUTA(11) => DataP_a_out_11_port, OUTA(10) => 
                           DataP_a_out_10_port, OUTA(9) => DataP_a_out_9_port, 
                           OUTA(8) => DataP_a_out_8_port, OUTA(7) => 
                           DataP_a_out_7_port, OUTA(6) => DataP_a_out_6_port, 
                           OUTA(5) => DataP_a_out_5_port, OUTA(4) => 
                           DataP_a_out_4_port, OUTA(3) => DataP_a_out_3_port, 
                           OUTA(2) => DataP_a_out_2_port, OUTA(1) => 
                           DataP_a_out_1_port, OUTA(0) => DataP_a_out_0_port, 
                           OUTB(31) => DataP_b_out_31_port, OUTB(30) => 
                           DataP_b_out_30_port, OUTB(29) => DataP_b_out_29_port
                           , OUTB(28) => DataP_b_out_28_port, OUTB(27) => 
                           DataP_b_out_27_port, OUTB(26) => DataP_b_out_26_port
                           , OUTB(25) => DataP_b_out_25_port, OUTB(24) => 
                           DataP_b_out_24_port, OUTB(23) => DataP_b_out_23_port
                           , OUTB(22) => DataP_b_out_22_port, OUTB(21) => 
                           DataP_b_out_21_port, OUTB(20) => DataP_b_out_20_port
                           , OUTB(19) => DataP_b_out_19_port, OUTB(18) => 
                           DataP_b_out_18_port, OUTB(17) => DataP_b_out_17_port
                           , OUTB(16) => DataP_b_out_16_port, OUTB(15) => 
                           DataP_b_out_15_port, OUTB(14) => DataP_b_out_14_port
                           , OUTB(13) => DataP_b_out_13_port, OUTB(12) => 
                           DataP_b_out_12_port, OUTB(11) => DataP_b_out_11_port
                           , OUTB(10) => DataP_b_out_10_port, OUTB(9) => 
                           DataP_b_out_9_port, OUTB(8) => DataP_b_out_8_port, 
                           OUTB(7) => DataP_b_out_7_port, OUTB(6) => 
                           DataP_b_out_6_port, OUTB(5) => DataP_b_out_5_port, 
                           OUTB(4) => DataP_b_out_4_port, OUTB(3) => 
                           DataP_b_out_3_port, OUTB(2) => DataP_b_out_2_port, 
                           OUTB(1) => DataP_b_out_1_port, OUTB(0) => 
                           DataP_b_out_0_port);
   DataP_BR_pred : branch_predictor port map( RST => Rst, PC_IN(31) => 
                           DataP_pc_out_31_port, PC_IN(30) => 
                           DataP_pc_out_30_port, PC_IN(29) => 
                           DataP_pc_out_29_port, PC_IN(28) => 
                           DataP_pc_out_28_port, PC_IN(27) => 
                           DataP_pc_out_27_port, PC_IN(26) => 
                           DataP_pc_out_26_port, PC_IN(25) => 
                           DataP_pc_out_25_port, PC_IN(24) => 
                           DataP_pc_out_24_port, PC_IN(23) => 
                           DataP_pc_out_23_port, PC_IN(22) => 
                           DataP_pc_out_22_port, PC_IN(21) => 
                           DataP_pc_out_21_port, PC_IN(20) => 
                           DataP_pc_out_20_port, PC_IN(19) => 
                           DataP_pc_out_19_port, PC_IN(18) => 
                           DataP_pc_out_18_port, PC_IN(17) => 
                           DataP_pc_out_17_port, PC_IN(16) => 
                           DataP_pc_out_16_port, PC_IN(15) => 
                           DataP_pc_out_15_port, PC_IN(14) => 
                           DataP_pc_out_14_port, PC_IN(13) => 
                           DataP_pc_out_13_port, PC_IN(12) => 
                           DataP_pc_out_12_port, PC_IN(11) => 
                           DataP_pc_out_11_port, PC_IN(10) => 
                           DataP_pc_out_10_port, PC_IN(9) => 
                           IRAM_ADDRESS_7_port, PC_IN(8) => IRAM_ADDRESS_6_port
                           , PC_IN(7) => IRAM_ADDRESS_5_port, PC_IN(6) => 
                           IRAM_ADDRESS_4_port, PC_IN(5) => IRAM_ADDRESS_3_port
                           , PC_IN(4) => IRAM_ADDRESS_2_port, PC_IN(3) => 
                           IRAM_ADDRESS_1_port, PC_IN(2) => IRAM_ADDRESS_0_port
                           , PC_IN(1) => DataP_pc_out_1, PC_IN(0) => 
                           DataP_pc_out_0, PC_FAIL(31) => DataP_npc_M_31_port, 
                           PC_FAIL(30) => DataP_npc_M_30_port, PC_FAIL(29) => 
                           DataP_npc_M_29_port, PC_FAIL(28) => 
                           DataP_npc_M_28_port, PC_FAIL(27) => 
                           DataP_npc_M_27_port, PC_FAIL(26) => 
                           DataP_npc_M_26_port, PC_FAIL(25) => 
                           DataP_npc_M_25_port, PC_FAIL(24) => 
                           DataP_npc_M_24_port, PC_FAIL(23) => 
                           DataP_npc_M_23_port, PC_FAIL(22) => 
                           DataP_npc_M_22_port, PC_FAIL(21) => 
                           DataP_npc_M_21_port, PC_FAIL(20) => 
                           DataP_npc_M_20_port, PC_FAIL(19) => 
                           DataP_npc_M_19_port, PC_FAIL(18) => 
                           DataP_npc_M_18_port, PC_FAIL(17) => 
                           DataP_npc_M_17_port, PC_FAIL(16) => 
                           DataP_npc_M_16_port, PC_FAIL(15) => 
                           DataP_npc_M_15_port, PC_FAIL(14) => 
                           DataP_npc_M_14_port, PC_FAIL(13) => 
                           DataP_npc_M_13_port, PC_FAIL(12) => 
                           DataP_npc_M_12_port, PC_FAIL(11) => 
                           DataP_npc_M_11_port, PC_FAIL(10) => 
                           DataP_npc_M_10_port, PC_FAIL(9) => 
                           DataP_npc_M_9_port, PC_FAIL(8) => DataP_npc_M_8_port
                           , PC_FAIL(7) => DataP_npc_M_7_port, PC_FAIL(6) => 
                           DataP_npc_M_6_port, PC_FAIL(5) => DataP_npc_M_5_port
                           , PC_FAIL(4) => DataP_npc_M_4_port, PC_FAIL(3) => 
                           DataP_npc_M_3_port, PC_FAIL(2) => DataP_npc_M_2_port
                           , PC_FAIL(1) => DataP_npc_M_1_port, PC_FAIL(0) => 
                           DataP_npc_M_0_port, IR_IN(31) => IRAM_DATA_OUT(31), 
                           IR_IN(30) => IRAM_DATA_OUT(30), IR_IN(29) => 
                           IRAM_DATA_OUT(29), IR_IN(28) => IRAM_DATA_OUT(28), 
                           IR_IN(27) => IRAM_DATA_OUT(27), IR_IN(26) => n4224, 
                           IR_IN(25) => IRAM_DATA_OUT(25), IR_IN(24) => 
                           IRAM_DATA_OUT(24), IR_IN(23) => IRAM_DATA_OUT(23), 
                           IR_IN(22) => IRAM_DATA_OUT(22), IR_IN(21) => 
                           IRAM_DATA_OUT(21), IR_IN(20) => IRAM_DATA_OUT(20), 
                           IR_IN(19) => IRAM_DATA_OUT(19), IR_IN(18) => 
                           IRAM_DATA_OUT(18), IR_IN(17) => IRAM_DATA_OUT(17), 
                           IR_IN(16) => IRAM_DATA_OUT(16), IR_IN(15) => 
                           IRAM_DATA_OUT(15), IR_IN(14) => IRAM_DATA_OUT(14), 
                           IR_IN(13) => IRAM_DATA_OUT(13), IR_IN(12) => 
                           IRAM_DATA_OUT(12), IR_IN(11) => IRAM_DATA_OUT(11), 
                           IR_IN(10) => IRAM_DATA_OUT(10), IR_IN(9) => 
                           IRAM_DATA_OUT(9), IR_IN(8) => IRAM_DATA_OUT(8), 
                           IR_IN(7) => IRAM_DATA_OUT(7), IR_IN(6) => 
                           IRAM_DATA_OUT(6), IR_IN(5) => IRAM_DATA_OUT(5), 
                           IR_IN(4) => IRAM_DATA_OUT(4), IR_IN(3) => 
                           IRAM_DATA_OUT(3), IR_IN(2) => IRAM_DATA_OUT(2), 
                           IR_IN(1) => IRAM_DATA_OUT(1), IR_IN(0) => 
                           IRAM_DATA_OUT(0), IR_FAIL(15) => DataP_IMM_s_15_port
                           , IR_FAIL(14) => DataP_IMM_s_14_port, IR_FAIL(13) =>
                           DataP_IMM_s_13_port, IR_FAIL(12) => 
                           DataP_IMM_s_12_port, IR_FAIL(11) => 
                           DataP_IMM_s_11_port, IR_FAIL(10) => 
                           DataP_IMM_s_10_port, IR_FAIL(9) => 
                           DataP_IMM_s_9_port, IR_FAIL(8) => DataP_IMM_s_8_port
                           , IR_FAIL(7) => DataP_IMM_s_7_port, IR_FAIL(6) => 
                           DataP_IMM_s_6_port, IR_FAIL(5) => DataP_IMM_s_5_port
                           , IR_FAIL(4) => DataP_IMM_s_4_port, IR_FAIL(3) => 
                           DataP_IMM_s_3_port, IR_FAIL(2) => DataP_IMM_s_2_port
                           , IR_FAIL(1) => DataP_IMM_s_1_port, IR_FAIL(0) => 
                           DataP_IMM_s_0_port, WRONG_PRE => DataP_wrong_br, 
                           RIGHT_PRE => DataP_right_br, NPC_OUT(31) => 
                           DataP_npc_pre_31_port, NPC_OUT(30) => 
                           DataP_npc_pre_30_port, NPC_OUT(29) => 
                           DataP_npc_pre_29_port, NPC_OUT(28) => 
                           DataP_npc_pre_28_port, NPC_OUT(27) => 
                           DataP_npc_pre_27_port, NPC_OUT(26) => 
                           DataP_npc_pre_26_port, NPC_OUT(25) => 
                           DataP_npc_pre_25_port, NPC_OUT(24) => 
                           DataP_npc_pre_24_port, NPC_OUT(23) => 
                           DataP_npc_pre_23_port, NPC_OUT(22) => 
                           DataP_npc_pre_22_port, NPC_OUT(21) => 
                           DataP_npc_pre_21_port, NPC_OUT(20) => 
                           DataP_npc_pre_20_port, NPC_OUT(19) => 
                           DataP_npc_pre_19_port, NPC_OUT(18) => 
                           DataP_npc_pre_18_port, NPC_OUT(17) => 
                           DataP_npc_pre_17_port, NPC_OUT(16) => 
                           DataP_npc_pre_16_port, NPC_OUT(15) => 
                           DataP_npc_pre_15_port, NPC_OUT(14) => 
                           DataP_npc_pre_14_port, NPC_OUT(13) => 
                           DataP_npc_pre_13_port, NPC_OUT(12) => 
                           DataP_npc_pre_12_port, NPC_OUT(11) => 
                           DataP_npc_pre_11_port, NPC_OUT(10) => 
                           DataP_npc_pre_10_port, NPC_OUT(9) => 
                           DataP_npc_pre_9_port, NPC_OUT(8) => 
                           DataP_npc_pre_8_port, NPC_OUT(7) => 
                           DataP_npc_pre_7_port, NPC_OUT(6) => 
                           DataP_npc_pre_6_port, NPC_OUT(5) => 
                           DataP_npc_pre_5_port, NPC_OUT(4) => 
                           DataP_npc_pre_4_port, NPC_OUT(3) => 
                           DataP_npc_pre_3_port, NPC_OUT(2) => 
                           DataP_npc_pre_2_port, NPC_OUT(1) => 
                           DataP_npc_pre_1_port, NPC_OUT(0) => 
                           DataP_npc_pre_0_port, LINK_ADD(31) => 
                           DataP_link_addr_F_31_port, LINK_ADD(30) => 
                           DataP_link_addr_F_30_port, LINK_ADD(29) => 
                           DataP_link_addr_F_29_port, LINK_ADD(28) => 
                           DataP_link_addr_F_28_port, LINK_ADD(27) => 
                           DataP_link_addr_F_27_port, LINK_ADD(26) => 
                           DataP_link_addr_F_26_port, LINK_ADD(25) => 
                           DataP_link_addr_F_25_port, LINK_ADD(24) => 
                           DataP_link_addr_F_24_port, LINK_ADD(23) => 
                           DataP_link_addr_F_23_port, LINK_ADD(22) => 
                           DataP_link_addr_F_22_port, LINK_ADD(21) => 
                           DataP_link_addr_F_21_port, LINK_ADD(20) => 
                           DataP_link_addr_F_20_port, LINK_ADD(19) => 
                           DataP_link_addr_F_19_port, LINK_ADD(18) => 
                           DataP_link_addr_F_18_port, LINK_ADD(17) => 
                           DataP_link_addr_F_17_port, LINK_ADD(16) => 
                           DataP_link_addr_F_16_port, LINK_ADD(15) => 
                           DataP_link_addr_F_15_port, LINK_ADD(14) => 
                           DataP_link_addr_F_14_port, LINK_ADD(13) => 
                           DataP_link_addr_F_13_port, LINK_ADD(12) => 
                           DataP_link_addr_F_12_port, LINK_ADD(11) => 
                           DataP_link_addr_F_11_port, LINK_ADD(10) => 
                           DataP_link_addr_F_10_port, LINK_ADD(9) => 
                           DataP_link_addr_F_9_port, LINK_ADD(8) => 
                           DataP_link_addr_F_8_port, LINK_ADD(7) => 
                           DataP_link_addr_F_7_port, LINK_ADD(6) => 
                           DataP_link_addr_F_6_port, LINK_ADD(5) => 
                           DataP_link_addr_F_5_port, LINK_ADD(4) => 
                           DataP_link_addr_F_4_port, LINK_ADD(3) => 
                           DataP_link_addr_F_3_port, LINK_ADD(2) => 
                           DataP_link_addr_F_2_port, LINK_ADD(1) => 
                           DataP_link_addr_F_1_port, LINK_ADD(0) => 
                           DataP_link_addr_F_0_port, SEL => DataP_npc_mux_sel, 
                           TAKEN => DataP_prediction);
   DataP_NPC_add_outPC_reg_0_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N1, Q => DataP_npc_0_port);
   DataP_NPC_add_outPC_reg_1_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N2, Q => DataP_npc_1_port);
   DataP_NPC_add_outPC_reg_2_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N3, Q => DataP_npc_2_port);
   DataP_NPC_add_outPC_reg_3_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N4, Q => DataP_npc_3_port);
   DataP_NPC_add_outPC_reg_4_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N5, Q => DataP_npc_4_port);
   DataP_NPC_add_outPC_reg_5_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N6, Q => DataP_npc_5_port);
   DataP_NPC_add_outPC_reg_6_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N7, Q => DataP_npc_6_port);
   DataP_NPC_add_outPC_reg_7_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N8, Q => DataP_npc_7_port);
   DataP_NPC_add_outPC_reg_8_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N9, Q => DataP_npc_8_port);
   DataP_NPC_add_outPC_reg_9_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N10, Q => DataP_npc_9_port);
   DataP_NPC_add_outPC_reg_10_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N11, Q => DataP_npc_10_port);
   DataP_NPC_add_outPC_reg_11_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N12, Q => DataP_npc_11_port);
   DataP_NPC_add_outPC_reg_12_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N13, Q => DataP_npc_12_port);
   DataP_NPC_add_outPC_reg_13_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N14, Q => DataP_npc_13_port);
   DataP_NPC_add_outPC_reg_14_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N15, Q => DataP_npc_14_port);
   DataP_NPC_add_outPC_reg_15_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N16, Q => DataP_npc_15_port);
   DataP_NPC_add_outPC_reg_16_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N17, Q => DataP_npc_16_port);
   DataP_NPC_add_outPC_reg_17_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N18, Q => DataP_npc_17_port);
   DataP_NPC_add_outPC_reg_18_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N19, Q => DataP_npc_18_port);
   DataP_NPC_add_outPC_reg_19_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N20, Q => DataP_npc_19_port);
   DataP_NPC_add_outPC_reg_20_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N21, Q => DataP_npc_20_port);
   DataP_NPC_add_outPC_reg_21_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N22, Q => DataP_npc_21_port);
   DataP_NPC_add_outPC_reg_22_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N23, Q => DataP_npc_22_port);
   DataP_NPC_add_outPC_reg_23_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N24, Q => DataP_npc_23_port);
   DataP_NPC_add_outPC_reg_24_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N25, Q => DataP_npc_24_port);
   DataP_NPC_add_outPC_reg_25_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N26, Q => DataP_npc_25_port);
   DataP_NPC_add_outPC_reg_26_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N27, Q => DataP_npc_26_port);
   DataP_NPC_add_outPC_reg_27_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N28, Q => DataP_npc_27_port);
   DataP_NPC_add_outPC_reg_28_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N29, Q => DataP_npc_28_port);
   DataP_NPC_add_outPC_reg_29_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N30, Q => DataP_npc_29_port);
   DataP_NPC_add_outPC_reg_30_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N31, Q => DataP_npc_30_port);
   DataP_NPC_add_outPC_reg_31_inst : DLH_X1 port map( G => DataP_NPC_add_N0, D 
                           => DataP_NPC_add_N32, Q => DataP_npc_31_port);
   DataP_MEM_WB_s_LMD_OUT_reg_0_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(0),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_0_port, QN 
                           => n_1004);
   DataP_MEM_WB_s_LMD_OUT_reg_1_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(1),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_1_port, QN 
                           => n_1005);
   DataP_MEM_WB_s_LMD_OUT_reg_2_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(2),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_2_port, QN 
                           => n_1006);
   DataP_MEM_WB_s_LMD_OUT_reg_3_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(3),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_3_port, QN 
                           => n_1007);
   DataP_MEM_WB_s_LMD_OUT_reg_4_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(4),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_4_port, QN 
                           => n_1008);
   DataP_MEM_WB_s_LMD_OUT_reg_5_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(5),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_5_port, QN 
                           => n_1009);
   DataP_MEM_WB_s_LMD_OUT_reg_6_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(6),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_6_port, QN 
                           => n_1010);
   DataP_MEM_WB_s_LMD_OUT_reg_7_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(7),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_7_port, QN 
                           => n_1011);
   DataP_MEM_WB_s_LMD_OUT_reg_8_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(8),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_8_port, QN 
                           => n_1012);
   DataP_MEM_WB_s_LMD_OUT_reg_9_inst : DFFR_X1 port map( D => DRAM_DATA_OUT(9),
                           CK => Clk, RN => Rst, Q => DataP_LMD_out_9_port, QN 
                           => n_1013);
   DataP_MEM_WB_s_LMD_OUT_reg_10_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(10), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_10_port, QN => n_1014);
   DataP_MEM_WB_s_LMD_OUT_reg_11_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(11), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_11_port, QN => n_1015);
   DataP_MEM_WB_s_LMD_OUT_reg_12_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(12), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_12_port, QN => n_1016);
   DataP_MEM_WB_s_LMD_OUT_reg_13_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(13), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_13_port, QN => n_1017);
   DataP_MEM_WB_s_LMD_OUT_reg_14_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(14), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_14_port, QN => n_1018);
   DataP_MEM_WB_s_LMD_OUT_reg_15_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(15), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_15_port, QN => n_1019);
   DataP_MEM_WB_s_LMD_OUT_reg_16_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(16), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_16_port, QN => n_1020);
   DataP_MEM_WB_s_LMD_OUT_reg_17_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(17), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_17_port, QN => n_1021);
   DataP_MEM_WB_s_LMD_OUT_reg_18_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(18), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_18_port, QN => n_1022);
   DataP_MEM_WB_s_LMD_OUT_reg_19_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(19), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_19_port, QN => n_1023);
   DataP_MEM_WB_s_LMD_OUT_reg_20_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(20), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_20_port, QN => n_1024);
   DataP_MEM_WB_s_LMD_OUT_reg_21_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(21), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_21_port, QN => n_1025);
   DataP_MEM_WB_s_LMD_OUT_reg_22_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(22), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_22_port, QN => n_1026);
   DataP_MEM_WB_s_LMD_OUT_reg_23_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(23), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_23_port, QN => n_1027);
   DataP_MEM_WB_s_LMD_OUT_reg_24_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(24), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_24_port, QN => n_1028);
   DataP_MEM_WB_s_LMD_OUT_reg_25_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(25), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_25_port, QN => n_1029);
   DataP_MEM_WB_s_LMD_OUT_reg_26_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(26), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_26_port, QN => n_1030);
   DataP_MEM_WB_s_LMD_OUT_reg_27_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(27), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_27_port, QN => n_1031);
   DataP_MEM_WB_s_LMD_OUT_reg_28_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(28), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_28_port, QN => n_1032);
   DataP_MEM_WB_s_LMD_OUT_reg_29_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(29), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_29_port, QN => n_1033);
   DataP_MEM_WB_s_LMD_OUT_reg_30_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(30), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_30_port, QN => n_1034);
   DataP_MEM_WB_s_LMD_OUT_reg_31_inst : DFFR_X1 port map( D => 
                           DRAM_DATA_OUT(31), CK => Clk, RN => Rst, Q => 
                           DataP_LMD_out_31_port, QN => n_1035);
   DataP_EX_MEM_s_ALU_OUT_reg_31_inst : DFFS_X1 port map( D => n297, CK => Clk,
                           SN => Rst, Q => n2414, QN => DataP_alu_out_M_31_port
                           );
   DataP_PC_reg_O_reg_31_inst : DFF_X1 port map( D => DataP_PC_reg_N33, CK => 
                           Clk, Q => DataP_pc_out_31_port, QN => n_1036);
   DataP_IF_IDs_NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => n1481, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_31_port, QN => 
                           n_1037);
   DataP_EX_MEM_s_NPC_L_OUT_reg_31_inst : DFFS_X1 port map( D => n292, CK => 
                           Clk, SN => Rst, Q => n291, QN => n_1038);
   DataP_MEM_WB_s_NPC_L_OUT_reg_31_inst : DFFS_X1 port map( D => n291, CK => 
                           Clk, SN => Rst, Q => n_1039, QN => 
                           DataP_link_addr_W_31_port);
   DataP_ID_EXs_B_OUT_reg_0_inst : DFFR_X1 port map( D => DataP_b_out_0_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_0_port, QN => 
                           n290);
   DataP_EX_MEM_s_B_OUT_reg_0_inst : DFFS_X1 port map( D => n290, CK => Clk, SN
                           => Rst, Q => n_1040, QN => DRAM_DATA_IN(0));
   DataP_ID_EXs_B_OUT_reg_1_inst : DFFR_X1 port map( D => DataP_b_out_1_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_1_port, QN => 
                           n289);
   DataP_EX_MEM_s_B_OUT_reg_1_inst : DFFS_X1 port map( D => n289, CK => Clk, SN
                           => Rst, Q => n_1041, QN => DRAM_DATA_IN(1));
   DataP_ID_EXs_B_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_b_out_2_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_2_port, QN => 
                           n288);
   DataP_EX_MEM_s_B_OUT_reg_2_inst : DFFS_X1 port map( D => n288, CK => Clk, SN
                           => Rst, Q => n_1042, QN => DRAM_DATA_IN(2));
   DataP_ID_EXs_B_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_b_out_3_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_3_port, QN => 
                           n287);
   DataP_EX_MEM_s_B_OUT_reg_3_inst : DFFS_X1 port map( D => n287, CK => Clk, SN
                           => Rst, Q => n_1043, QN => DRAM_DATA_IN(3));
   DataP_ID_EXs_B_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_b_out_4_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_4_port, QN => 
                           n286);
   DataP_EX_MEM_s_B_OUT_reg_4_inst : DFFS_X1 port map( D => n286, CK => Clk, SN
                           => Rst, Q => n_1044, QN => DRAM_DATA_IN(4));
   DataP_ID_EXs_B_OUT_reg_5_inst : DFFR_X1 port map( D => DataP_b_out_5_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_5_port, QN => 
                           n285);
   DataP_EX_MEM_s_B_OUT_reg_5_inst : DFFS_X1 port map( D => n285, CK => Clk, SN
                           => Rst, Q => n_1045, QN => DRAM_DATA_IN(5));
   DataP_ID_EXs_B_OUT_reg_6_inst : DFFR_X1 port map( D => DataP_b_out_6_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_6_port, QN => 
                           n284);
   DataP_EX_MEM_s_B_OUT_reg_6_inst : DFFS_X1 port map( D => n284, CK => Clk, SN
                           => Rst, Q => n_1046, QN => DRAM_DATA_IN(6));
   DataP_ID_EXs_B_OUT_reg_7_inst : DFFR_X1 port map( D => DataP_b_out_7_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_7_port, QN => 
                           n283);
   DataP_EX_MEM_s_B_OUT_reg_7_inst : DFFS_X1 port map( D => n283, CK => Clk, SN
                           => Rst, Q => n_1047, QN => DRAM_DATA_IN(7));
   DataP_ID_EXs_B_OUT_reg_8_inst : DFFR_X1 port map( D => DataP_b_out_8_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_8_port, QN => 
                           n282);
   DataP_EX_MEM_s_B_OUT_reg_8_inst : DFFS_X1 port map( D => n282, CK => Clk, SN
                           => Rst, Q => n_1048, QN => DRAM_DATA_IN(8));
   DataP_ID_EXs_B_OUT_reg_9_inst : DFFR_X1 port map( D => DataP_b_out_9_port, 
                           CK => Clk, RN => Rst, Q => DataP_B_s_9_port, QN => 
                           n281);
   DataP_EX_MEM_s_B_OUT_reg_9_inst : DFFS_X1 port map( D => n281, CK => Clk, SN
                           => Rst, Q => n_1049, QN => DRAM_DATA_IN(9));
   DataP_ID_EXs_B_OUT_reg_10_inst : DFFR_X1 port map( D => DataP_b_out_10_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_10_port, QN => 
                           n280);
   DataP_EX_MEM_s_B_OUT_reg_10_inst : DFFS_X1 port map( D => n280, CK => Clk, 
                           SN => Rst, Q => n_1050, QN => DRAM_DATA_IN(10));
   DataP_ID_EXs_B_OUT_reg_11_inst : DFFR_X1 port map( D => DataP_b_out_11_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_11_port, QN => 
                           n279);
   DataP_EX_MEM_s_B_OUT_reg_11_inst : DFFS_X1 port map( D => n279, CK => Clk, 
                           SN => Rst, Q => n_1051, QN => DRAM_DATA_IN(11));
   DataP_ID_EXs_B_OUT_reg_12_inst : DFFR_X1 port map( D => DataP_b_out_12_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_12_port, QN => 
                           n278);
   DataP_EX_MEM_s_B_OUT_reg_12_inst : DFFS_X1 port map( D => n278, CK => Clk, 
                           SN => Rst, Q => n_1052, QN => DRAM_DATA_IN(12));
   DataP_ID_EXs_B_OUT_reg_13_inst : DFFR_X1 port map( D => DataP_b_out_13_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_13_port, QN => 
                           n277);
   DataP_EX_MEM_s_B_OUT_reg_13_inst : DFFS_X1 port map( D => n277, CK => Clk, 
                           SN => Rst, Q => n_1053, QN => DRAM_DATA_IN(13));
   DataP_ID_EXs_B_OUT_reg_14_inst : DFFR_X1 port map( D => DataP_b_out_14_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_14_port, QN => 
                           n276);
   DataP_EX_MEM_s_B_OUT_reg_14_inst : DFFS_X1 port map( D => n276, CK => Clk, 
                           SN => Rst, Q => n_1054, QN => DRAM_DATA_IN(14));
   DataP_ID_EXs_B_OUT_reg_15_inst : DFFR_X1 port map( D => DataP_b_out_15_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_15_port, QN => 
                           n275);
   DataP_EX_MEM_s_B_OUT_reg_15_inst : DFFS_X1 port map( D => n275, CK => Clk, 
                           SN => Rst, Q => n_1055, QN => DRAM_DATA_IN(15));
   DataP_ID_EXs_B_OUT_reg_16_inst : DFFR_X1 port map( D => DataP_b_out_16_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_16_port, QN => 
                           n274);
   DataP_EX_MEM_s_B_OUT_reg_16_inst : DFFS_X1 port map( D => n274, CK => Clk, 
                           SN => Rst, Q => n_1056, QN => DRAM_DATA_IN(16));
   DataP_ID_EXs_B_OUT_reg_17_inst : DFFR_X1 port map( D => DataP_b_out_17_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_17_port, QN => 
                           n273);
   DataP_EX_MEM_s_B_OUT_reg_17_inst : DFFS_X1 port map( D => n273, CK => Clk, 
                           SN => Rst, Q => n_1057, QN => DRAM_DATA_IN(17));
   DataP_ID_EXs_B_OUT_reg_18_inst : DFFR_X1 port map( D => DataP_b_out_18_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_18_port, QN => 
                           n272);
   DataP_EX_MEM_s_B_OUT_reg_18_inst : DFFS_X1 port map( D => n272, CK => Clk, 
                           SN => Rst, Q => n_1058, QN => DRAM_DATA_IN(18));
   DataP_ID_EXs_B_OUT_reg_19_inst : DFFR_X1 port map( D => DataP_b_out_19_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_19_port, QN => 
                           n271);
   DataP_EX_MEM_s_B_OUT_reg_19_inst : DFFS_X1 port map( D => n271, CK => Clk, 
                           SN => Rst, Q => n_1059, QN => DRAM_DATA_IN(19));
   DataP_ID_EXs_B_OUT_reg_20_inst : DFFR_X1 port map( D => DataP_b_out_20_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_20_port, QN => 
                           n270);
   DataP_EX_MEM_s_B_OUT_reg_20_inst : DFFS_X1 port map( D => n270, CK => Clk, 
                           SN => Rst, Q => n_1060, QN => DRAM_DATA_IN(20));
   DataP_ID_EXs_B_OUT_reg_21_inst : DFFR_X1 port map( D => DataP_b_out_21_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_21_port, QN => 
                           n269);
   DataP_EX_MEM_s_B_OUT_reg_21_inst : DFFS_X1 port map( D => n269, CK => Clk, 
                           SN => Rst, Q => n_1061, QN => DRAM_DATA_IN(21));
   DataP_ID_EXs_B_OUT_reg_22_inst : DFFR_X1 port map( D => DataP_b_out_22_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_22_port, QN => 
                           n268);
   DataP_EX_MEM_s_B_OUT_reg_22_inst : DFFS_X1 port map( D => n268, CK => Clk, 
                           SN => Rst, Q => n_1062, QN => DRAM_DATA_IN(22));
   DataP_ID_EXs_B_OUT_reg_23_inst : DFFR_X1 port map( D => DataP_b_out_23_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_23_port, QN => 
                           n267);
   DataP_EX_MEM_s_B_OUT_reg_23_inst : DFFS_X1 port map( D => n267, CK => Clk, 
                           SN => Rst, Q => n_1063, QN => DRAM_DATA_IN(23));
   DataP_ID_EXs_B_OUT_reg_24_inst : DFFR_X1 port map( D => DataP_b_out_24_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_24_port, QN => 
                           n266);
   DataP_EX_MEM_s_B_OUT_reg_24_inst : DFFS_X1 port map( D => n266, CK => Clk, 
                           SN => Rst, Q => n_1064, QN => DRAM_DATA_IN(24));
   DataP_ID_EXs_B_OUT_reg_25_inst : DFFR_X1 port map( D => DataP_b_out_25_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_25_port, QN => 
                           n265);
   DataP_EX_MEM_s_B_OUT_reg_25_inst : DFFS_X1 port map( D => n265, CK => Clk, 
                           SN => Rst, Q => n_1065, QN => DRAM_DATA_IN(25));
   DataP_ID_EXs_B_OUT_reg_26_inst : DFFR_X1 port map( D => DataP_b_out_26_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_26_port, QN => 
                           n264);
   DataP_EX_MEM_s_B_OUT_reg_26_inst : DFFS_X1 port map( D => n264, CK => Clk, 
                           SN => Rst, Q => n_1066, QN => DRAM_DATA_IN(26));
   DataP_ID_EXs_B_OUT_reg_27_inst : DFFR_X1 port map( D => DataP_b_out_27_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_27_port, QN => 
                           n263);
   DataP_EX_MEM_s_B_OUT_reg_27_inst : DFFS_X1 port map( D => n263, CK => Clk, 
                           SN => Rst, Q => n_1067, QN => DRAM_DATA_IN(27));
   DataP_ID_EXs_B_OUT_reg_28_inst : DFFR_X1 port map( D => DataP_b_out_28_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_28_port, QN => 
                           n262);
   DataP_EX_MEM_s_B_OUT_reg_28_inst : DFFS_X1 port map( D => n262, CK => Clk, 
                           SN => Rst, Q => n_1068, QN => DRAM_DATA_IN(28));
   DataP_ID_EXs_B_OUT_reg_29_inst : DFFR_X1 port map( D => DataP_b_out_29_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_29_port, QN => 
                           n261);
   DataP_EX_MEM_s_B_OUT_reg_29_inst : DFFS_X1 port map( D => n261, CK => Clk, 
                           SN => Rst, Q => n_1069, QN => DRAM_DATA_IN(29));
   DataP_ID_EXs_B_OUT_reg_30_inst : DFFR_X1 port map( D => DataP_b_out_30_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_30_port, QN => 
                           n260);
   DataP_EX_MEM_s_B_OUT_reg_30_inst : DFFS_X1 port map( D => n260, CK => Clk, 
                           SN => Rst, Q => n_1070, QN => DRAM_DATA_IN(30));
   DataP_ID_EXs_B_OUT_reg_31_inst : DFFR_X1 port map( D => DataP_b_out_31_port,
                           CK => Clk, RN => Rst, Q => DataP_B_s_31_port, QN => 
                           n259);
   DataP_EX_MEM_s_B_OUT_reg_31_inst : DFFS_X1 port map( D => n259, CK => Clk, 
                           SN => Rst, Q => n_1071, QN => DRAM_DATA_IN(31));
   DataP_ID_EXs_A_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_a_out_2_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_2_port, QN => 
                           n2459);
   DataP_ID_EXs_A_OUT_reg_8_inst : DFFR_X1 port map( D => DataP_a_out_8_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_8_port, QN => 
                           n2467);
   DataP_ID_EXs_A_OUT_reg_9_inst : DFFR_X1 port map( D => DataP_a_out_9_port, 
                           CK => Clk, RN => Rst, Q => DataP_A_s_9_port, QN => 
                           n2435);
   DataP_EX_MEM_s_ALU_OUT_reg_15_inst : DFFS_X1 port map( D => n330, CK => Clk,
                           SN => Rst, Q => n2433, QN => DataP_alu_out_M_15_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_19_inst : DFFS_X1 port map( D => n319, CK => Clk,
                           SN => Rst, Q => n2421, QN => DataP_alu_out_M_19_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_30_inst : DFFS_X1 port map( D => n2774, CK => Clk
                           , SN => Rst, Q => n2417, QN => 
                           DataP_alu_out_M_30_port);
   DataP_IF_IDs_PR_OUT_reg : DFFR_X1 port map( D => n1449, CK => Clk, RN => Rst
                           , Q => DataP_pr_D, QN => n_1072);
   DataP_IF_IDs_NPC_L_OUT_reg_30_inst : DFFR_X1 port map( D => n1450, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_30_port, QN => 
                           n257);
   DataP_ID_EXs_NPC_L_OUT_reg_30_inst : DFFS_X1 port map( D => n257, CK => Clk,
                           SN => Rst, Q => n256, QN => n_1073);
   DataP_EX_MEM_s_NPC_L_OUT_reg_30_inst : DFFS_X1 port map( D => n256, CK => 
                           Clk, SN => Rst, Q => n255, QN => n_1074);
   DataP_MEM_WB_s_NPC_L_OUT_reg_30_inst : DFFS_X1 port map( D => n255, CK => 
                           Clk, SN => Rst, Q => n_1075, QN => 
                           DataP_link_addr_W_30_port);
   DataP_IF_IDs_NPC_L_OUT_reg_29_inst : DFFR_X1 port map( D => n1451, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_29_port, QN => 
                           n254);
   DataP_ID_EXs_NPC_L_OUT_reg_29_inst : DFFS_X1 port map( D => n254, CK => Clk,
                           SN => Rst, Q => n253, QN => n_1076);
   DataP_EX_MEM_s_NPC_L_OUT_reg_29_inst : DFFS_X1 port map( D => n253, CK => 
                           Clk, SN => Rst, Q => n252, QN => n_1077);
   DataP_MEM_WB_s_NPC_L_OUT_reg_29_inst : DFFS_X1 port map( D => n252, CK => 
                           Clk, SN => Rst, Q => n_1078, QN => 
                           DataP_link_addr_W_29_port);
   DataP_IF_IDs_NPC_L_OUT_reg_28_inst : DFFR_X1 port map( D => n1452, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_28_port, QN => 
                           n251);
   DataP_ID_EXs_NPC_L_OUT_reg_28_inst : DFFS_X1 port map( D => n251, CK => Clk,
                           SN => Rst, Q => n250, QN => n_1079);
   DataP_EX_MEM_s_NPC_L_OUT_reg_28_inst : DFFS_X1 port map( D => n250, CK => 
                           Clk, SN => Rst, Q => n249, QN => n_1080);
   DataP_MEM_WB_s_NPC_L_OUT_reg_28_inst : DFFS_X1 port map( D => n249, CK => 
                           Clk, SN => Rst, Q => n_1081, QN => 
                           DataP_link_addr_W_28_port);
   DataP_IF_IDs_NPC_L_OUT_reg_27_inst : DFFR_X1 port map( D => n1453, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_27_port, QN => 
                           n248);
   DataP_ID_EXs_NPC_L_OUT_reg_27_inst : DFFS_X1 port map( D => n248, CK => Clk,
                           SN => Rst, Q => n247, QN => n_1082);
   DataP_EX_MEM_s_NPC_L_OUT_reg_27_inst : DFFS_X1 port map( D => n247, CK => 
                           Clk, SN => Rst, Q => n246, QN => n_1083);
   DataP_MEM_WB_s_NPC_L_OUT_reg_27_inst : DFFS_X1 port map( D => n246, CK => 
                           Clk, SN => Rst, Q => n_1084, QN => 
                           DataP_link_addr_W_27_port);
   DataP_IF_IDs_NPC_L_OUT_reg_26_inst : DFFR_X1 port map( D => n1454, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_26_port, QN => 
                           n245);
   DataP_ID_EXs_NPC_L_OUT_reg_26_inst : DFFS_X1 port map( D => n245, CK => Clk,
                           SN => Rst, Q => n244, QN => n_1085);
   DataP_EX_MEM_s_NPC_L_OUT_reg_26_inst : DFFS_X1 port map( D => n244, CK => 
                           Clk, SN => Rst, Q => n243, QN => n_1086);
   DataP_MEM_WB_s_NPC_L_OUT_reg_26_inst : DFFS_X1 port map( D => n243, CK => 
                           Clk, SN => Rst, Q => n_1087, QN => 
                           DataP_link_addr_W_26_port);
   DataP_IF_IDs_NPC_L_OUT_reg_25_inst : DFFR_X1 port map( D => n1455, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_25_port, QN => 
                           n242);
   DataP_ID_EXs_NPC_L_OUT_reg_25_inst : DFFS_X1 port map( D => n242, CK => Clk,
                           SN => Rst, Q => n241, QN => n_1088);
   DataP_EX_MEM_s_NPC_L_OUT_reg_25_inst : DFFS_X1 port map( D => n241, CK => 
                           Clk, SN => Rst, Q => n240, QN => n_1089);
   DataP_MEM_WB_s_NPC_L_OUT_reg_25_inst : DFFS_X1 port map( D => n240, CK => 
                           Clk, SN => Rst, Q => n_1090, QN => 
                           DataP_link_addr_W_25_port);
   DataP_IF_IDs_NPC_L_OUT_reg_24_inst : DFFR_X1 port map( D => n1456, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_24_port, QN => 
                           n239);
   DataP_ID_EXs_NPC_L_OUT_reg_24_inst : DFFS_X1 port map( D => n239, CK => Clk,
                           SN => Rst, Q => n238, QN => n_1091);
   DataP_EX_MEM_s_NPC_L_OUT_reg_24_inst : DFFS_X1 port map( D => n238, CK => 
                           Clk, SN => Rst, Q => n237, QN => n_1092);
   DataP_MEM_WB_s_NPC_L_OUT_reg_24_inst : DFFS_X1 port map( D => n237, CK => 
                           Clk, SN => Rst, Q => n_1093, QN => 
                           DataP_link_addr_W_24_port);
   DataP_IF_IDs_NPC_L_OUT_reg_23_inst : DFFR_X1 port map( D => n1457, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_23_port, QN => 
                           n236);
   DataP_ID_EXs_NPC_L_OUT_reg_23_inst : DFFS_X1 port map( D => n236, CK => Clk,
                           SN => Rst, Q => n235, QN => n_1094);
   DataP_EX_MEM_s_NPC_L_OUT_reg_23_inst : DFFS_X1 port map( D => n235, CK => 
                           Clk, SN => Rst, Q => n234, QN => n_1095);
   DataP_MEM_WB_s_NPC_L_OUT_reg_23_inst : DFFS_X1 port map( D => n234, CK => 
                           Clk, SN => Rst, Q => n_1096, QN => 
                           DataP_link_addr_W_23_port);
   DataP_IF_IDs_NPC_L_OUT_reg_22_inst : DFFR_X1 port map( D => n1458, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_22_port, QN => 
                           n233);
   DataP_ID_EXs_NPC_L_OUT_reg_22_inst : DFFS_X1 port map( D => n233, CK => Clk,
                           SN => Rst, Q => n232, QN => n_1097);
   DataP_EX_MEM_s_NPC_L_OUT_reg_22_inst : DFFS_X1 port map( D => n232, CK => 
                           Clk, SN => Rst, Q => n231, QN => n_1098);
   DataP_MEM_WB_s_NPC_L_OUT_reg_22_inst : DFFS_X1 port map( D => n231, CK => 
                           Clk, SN => Rst, Q => n_1099, QN => 
                           DataP_link_addr_W_22_port);
   DataP_IF_IDs_NPC_L_OUT_reg_21_inst : DFFR_X1 port map( D => n1459, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_21_port, QN => 
                           n230);
   DataP_ID_EXs_NPC_L_OUT_reg_21_inst : DFFS_X1 port map( D => n230, CK => Clk,
                           SN => Rst, Q => n229, QN => n_1100);
   DataP_EX_MEM_s_NPC_L_OUT_reg_21_inst : DFFS_X1 port map( D => n229, CK => 
                           Clk, SN => Rst, Q => n228, QN => n_1101);
   DataP_MEM_WB_s_NPC_L_OUT_reg_21_inst : DFFS_X1 port map( D => n228, CK => 
                           Clk, SN => Rst, Q => n_1102, QN => 
                           DataP_link_addr_W_21_port);
   DataP_IF_IDs_NPC_L_OUT_reg_20_inst : DFFR_X1 port map( D => n1460, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_20_port, QN => 
                           n227);
   DataP_ID_EXs_NPC_L_OUT_reg_20_inst : DFFS_X1 port map( D => n227, CK => Clk,
                           SN => Rst, Q => n226, QN => n_1103);
   DataP_EX_MEM_s_NPC_L_OUT_reg_20_inst : DFFS_X1 port map( D => n226, CK => 
                           Clk, SN => Rst, Q => n225, QN => n_1104);
   DataP_MEM_WB_s_NPC_L_OUT_reg_20_inst : DFFS_X1 port map( D => n225, CK => 
                           Clk, SN => Rst, Q => n_1105, QN => 
                           DataP_link_addr_W_20_port);
   DataP_IF_IDs_NPC_L_OUT_reg_19_inst : DFFR_X1 port map( D => n1461, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_19_port, QN => 
                           n224);
   DataP_ID_EXs_NPC_L_OUT_reg_19_inst : DFFS_X1 port map( D => n224, CK => Clk,
                           SN => Rst, Q => n223, QN => n_1106);
   DataP_EX_MEM_s_NPC_L_OUT_reg_19_inst : DFFS_X1 port map( D => n223, CK => 
                           Clk, SN => Rst, Q => n222, QN => n_1107);
   DataP_MEM_WB_s_NPC_L_OUT_reg_19_inst : DFFS_X1 port map( D => n222, CK => 
                           Clk, SN => Rst, Q => n_1108, QN => 
                           DataP_link_addr_W_19_port);
   DataP_IF_IDs_NPC_L_OUT_reg_18_inst : DFFR_X1 port map( D => n1462, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_18_port, QN => 
                           n221);
   DataP_ID_EXs_NPC_L_OUT_reg_18_inst : DFFS_X1 port map( D => n221, CK => Clk,
                           SN => Rst, Q => n220, QN => n_1109);
   DataP_EX_MEM_s_NPC_L_OUT_reg_18_inst : DFFS_X1 port map( D => n220, CK => 
                           Clk, SN => Rst, Q => n219, QN => n_1110);
   DataP_MEM_WB_s_NPC_L_OUT_reg_18_inst : DFFS_X1 port map( D => n219, CK => 
                           Clk, SN => Rst, Q => n_1111, QN => 
                           DataP_link_addr_W_18_port);
   DataP_IF_IDs_NPC_L_OUT_reg_17_inst : DFFR_X1 port map( D => n1463, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_17_port, QN => 
                           n218);
   DataP_ID_EXs_NPC_L_OUT_reg_17_inst : DFFS_X1 port map( D => n218, CK => Clk,
                           SN => Rst, Q => n217, QN => n_1112);
   DataP_EX_MEM_s_NPC_L_OUT_reg_17_inst : DFFS_X1 port map( D => n217, CK => 
                           Clk, SN => Rst, Q => n216, QN => n_1113);
   DataP_MEM_WB_s_NPC_L_OUT_reg_17_inst : DFFS_X1 port map( D => n216, CK => 
                           Clk, SN => Rst, Q => n_1114, QN => 
                           DataP_link_addr_W_17_port);
   DataP_IF_IDs_NPC_L_OUT_reg_16_inst : DFFR_X1 port map( D => n1464, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_16_port, QN => 
                           n215);
   DataP_ID_EXs_NPC_L_OUT_reg_16_inst : DFFS_X1 port map( D => n215, CK => Clk,
                           SN => Rst, Q => n214, QN => n_1115);
   DataP_EX_MEM_s_NPC_L_OUT_reg_16_inst : DFFS_X1 port map( D => n214, CK => 
                           Clk, SN => Rst, Q => n213, QN => n_1116);
   DataP_MEM_WB_s_NPC_L_OUT_reg_16_inst : DFFS_X1 port map( D => n213, CK => 
                           Clk, SN => Rst, Q => n_1117, QN => 
                           DataP_link_addr_W_16_port);
   DataP_IF_IDs_NPC_L_OUT_reg_15_inst : DFFR_X1 port map( D => n1465, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_15_port, QN => 
                           n212);
   DataP_ID_EXs_NPC_L_OUT_reg_15_inst : DFFS_X1 port map( D => n212, CK => Clk,
                           SN => Rst, Q => n211, QN => n_1118);
   DataP_EX_MEM_s_NPC_L_OUT_reg_15_inst : DFFS_X1 port map( D => n211, CK => 
                           Clk, SN => Rst, Q => n210, QN => n_1119);
   DataP_MEM_WB_s_NPC_L_OUT_reg_15_inst : DFFS_X1 port map( D => n210, CK => 
                           Clk, SN => Rst, Q => n_1120, QN => 
                           DataP_link_addr_W_15_port);
   DataP_IF_IDs_NPC_L_OUT_reg_14_inst : DFFR_X1 port map( D => n1466, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_14_port, QN => 
                           n209);
   DataP_ID_EXs_NPC_L_OUT_reg_14_inst : DFFS_X1 port map( D => n209, CK => Clk,
                           SN => Rst, Q => n208, QN => n_1121);
   DataP_EX_MEM_s_NPC_L_OUT_reg_14_inst : DFFS_X1 port map( D => n208, CK => 
                           Clk, SN => Rst, Q => n207, QN => n_1122);
   DataP_MEM_WB_s_NPC_L_OUT_reg_14_inst : DFFS_X1 port map( D => n207, CK => 
                           Clk, SN => Rst, Q => n_1123, QN => 
                           DataP_link_addr_W_14_port);
   DataP_IF_IDs_NPC_L_OUT_reg_13_inst : DFFR_X1 port map( D => n1467, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_13_port, QN => 
                           n206);
   DataP_ID_EXs_NPC_L_OUT_reg_13_inst : DFFS_X1 port map( D => n206, CK => Clk,
                           SN => Rst, Q => n205, QN => n_1124);
   DataP_EX_MEM_s_NPC_L_OUT_reg_13_inst : DFFS_X1 port map( D => n205, CK => 
                           Clk, SN => Rst, Q => n204, QN => n_1125);
   DataP_MEM_WB_s_NPC_L_OUT_reg_13_inst : DFFS_X1 port map( D => n204, CK => 
                           Clk, SN => Rst, Q => n_1126, QN => 
                           DataP_link_addr_W_13_port);
   DataP_IF_IDs_NPC_L_OUT_reg_12_inst : DFFR_X1 port map( D => n1468, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_12_port, QN => 
                           n203);
   DataP_ID_EXs_NPC_L_OUT_reg_12_inst : DFFS_X1 port map( D => n203, CK => Clk,
                           SN => Rst, Q => n202, QN => n_1127);
   DataP_EX_MEM_s_NPC_L_OUT_reg_12_inst : DFFS_X1 port map( D => n202, CK => 
                           Clk, SN => Rst, Q => n201, QN => n_1128);
   DataP_MEM_WB_s_NPC_L_OUT_reg_12_inst : DFFS_X1 port map( D => n201, CK => 
                           Clk, SN => Rst, Q => n_1129, QN => 
                           DataP_link_addr_W_12_port);
   DataP_IF_IDs_NPC_L_OUT_reg_11_inst : DFFR_X1 port map( D => n1469, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_11_port, QN => 
                           n200);
   DataP_ID_EXs_NPC_L_OUT_reg_11_inst : DFFS_X1 port map( D => n200, CK => Clk,
                           SN => Rst, Q => n199, QN => n_1130);
   DataP_EX_MEM_s_NPC_L_OUT_reg_11_inst : DFFS_X1 port map( D => n199, CK => 
                           Clk, SN => Rst, Q => n198, QN => n_1131);
   DataP_MEM_WB_s_NPC_L_OUT_reg_11_inst : DFFS_X1 port map( D => n198, CK => 
                           Clk, SN => Rst, Q => n_1132, QN => 
                           DataP_link_addr_W_11_port);
   DataP_IF_IDs_NPC_L_OUT_reg_10_inst : DFFR_X1 port map( D => n1470, CK => Clk
                           , RN => Rst, Q => DataP_link_addr_D_10_port, QN => 
                           n197);
   DataP_ID_EXs_NPC_L_OUT_reg_10_inst : DFFS_X1 port map( D => n197, CK => Clk,
                           SN => Rst, Q => n196, QN => n_1133);
   DataP_EX_MEM_s_NPC_L_OUT_reg_10_inst : DFFS_X1 port map( D => n196, CK => 
                           Clk, SN => Rst, Q => n195, QN => n_1134);
   DataP_MEM_WB_s_NPC_L_OUT_reg_10_inst : DFFS_X1 port map( D => n195, CK => 
                           Clk, SN => Rst, Q => n_1135, QN => 
                           DataP_link_addr_W_10_port);
   DataP_IF_IDs_NPC_L_OUT_reg_9_inst : DFFR_X1 port map( D => n1471, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_9_port, QN => n194
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_9_inst : DFFS_X1 port map( D => n194, CK => Clk, 
                           SN => Rst, Q => n193, QN => n_1136);
   DataP_EX_MEM_s_NPC_L_OUT_reg_9_inst : DFFS_X1 port map( D => n193, CK => Clk
                           , SN => Rst, Q => n192, QN => n_1137);
   DataP_MEM_WB_s_NPC_L_OUT_reg_9_inst : DFFS_X1 port map( D => n192, CK => Clk
                           , SN => Rst, Q => n_1138, QN => 
                           DataP_link_addr_W_9_port);
   DataP_IF_IDs_NPC_L_OUT_reg_8_inst : DFFR_X1 port map( D => n1472, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_8_port, QN => n191
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_8_inst : DFFS_X1 port map( D => n191, CK => Clk, 
                           SN => Rst, Q => n190, QN => n_1139);
   DataP_EX_MEM_s_NPC_L_OUT_reg_8_inst : DFFS_X1 port map( D => n190, CK => Clk
                           , SN => Rst, Q => n189, QN => n_1140);
   DataP_MEM_WB_s_NPC_L_OUT_reg_8_inst : DFFS_X1 port map( D => n189, CK => Clk
                           , SN => Rst, Q => n_1141, QN => 
                           DataP_link_addr_W_8_port);
   DataP_IF_IDs_NPC_L_OUT_reg_7_inst : DFFR_X1 port map( D => n1473, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_7_port, QN => n188
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_7_inst : DFFS_X1 port map( D => n188, CK => Clk, 
                           SN => Rst, Q => n187, QN => n_1142);
   DataP_EX_MEM_s_NPC_L_OUT_reg_7_inst : DFFS_X1 port map( D => n187, CK => Clk
                           , SN => Rst, Q => n186, QN => n_1143);
   DataP_MEM_WB_s_NPC_L_OUT_reg_7_inst : DFFS_X1 port map( D => n186, CK => Clk
                           , SN => Rst, Q => n_1144, QN => 
                           DataP_link_addr_W_7_port);
   DataP_IF_IDs_NPC_L_OUT_reg_6_inst : DFFR_X1 port map( D => n1474, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_6_port, QN => n185
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_6_inst : DFFS_X1 port map( D => n185, CK => Clk, 
                           SN => Rst, Q => n184, QN => n_1145);
   DataP_EX_MEM_s_NPC_L_OUT_reg_6_inst : DFFS_X1 port map( D => n184, CK => Clk
                           , SN => Rst, Q => n183, QN => n_1146);
   DataP_MEM_WB_s_NPC_L_OUT_reg_6_inst : DFFS_X1 port map( D => n183, CK => Clk
                           , SN => Rst, Q => n_1147, QN => 
                           DataP_link_addr_W_6_port);
   DataP_IF_IDs_NPC_L_OUT_reg_5_inst : DFFR_X1 port map( D => n1475, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_5_port, QN => n182
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_5_inst : DFFS_X1 port map( D => n182, CK => Clk, 
                           SN => Rst, Q => n181, QN => n_1148);
   DataP_EX_MEM_s_NPC_L_OUT_reg_5_inst : DFFS_X1 port map( D => n181, CK => Clk
                           , SN => Rst, Q => n180, QN => n_1149);
   DataP_MEM_WB_s_NPC_L_OUT_reg_5_inst : DFFS_X1 port map( D => n180, CK => Clk
                           , SN => Rst, Q => n_1150, QN => 
                           DataP_link_addr_W_5_port);
   DataP_IF_IDs_NPC_L_OUT_reg_4_inst : DFFR_X1 port map( D => n1476, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_4_port, QN => n179
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_4_inst : DFFS_X1 port map( D => n179, CK => Clk, 
                           SN => Rst, Q => n178, QN => n_1151);
   DataP_EX_MEM_s_NPC_L_OUT_reg_4_inst : DFFS_X1 port map( D => n178, CK => Clk
                           , SN => Rst, Q => n177, QN => n_1152);
   DataP_MEM_WB_s_NPC_L_OUT_reg_4_inst : DFFS_X1 port map( D => n177, CK => Clk
                           , SN => Rst, Q => n_1153, QN => 
                           DataP_link_addr_W_4_port);
   DataP_IF_IDs_NPC_L_OUT_reg_3_inst : DFFR_X1 port map( D => n1477, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_3_port, QN => n176
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_3_inst : DFFS_X1 port map( D => n176, CK => Clk, 
                           SN => Rst, Q => n175, QN => n_1154);
   DataP_EX_MEM_s_NPC_L_OUT_reg_3_inst : DFFS_X1 port map( D => n175, CK => Clk
                           , SN => Rst, Q => n174, QN => n_1155);
   DataP_MEM_WB_s_NPC_L_OUT_reg_3_inst : DFFS_X1 port map( D => n174, CK => Clk
                           , SN => Rst, Q => n_1156, QN => 
                           DataP_link_addr_W_3_port);
   DataP_IF_IDs_NPC_L_OUT_reg_2_inst : DFFR_X1 port map( D => n1478, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_2_port, QN => n173
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_2_inst : DFFS_X1 port map( D => n173, CK => Clk, 
                           SN => Rst, Q => n172, QN => n_1157);
   DataP_EX_MEM_s_NPC_L_OUT_reg_2_inst : DFFS_X1 port map( D => n172, CK => Clk
                           , SN => Rst, Q => n171, QN => n_1158);
   DataP_MEM_WB_s_NPC_L_OUT_reg_2_inst : DFFS_X1 port map( D => n171, CK => Clk
                           , SN => Rst, Q => n_1159, QN => 
                           DataP_link_addr_W_2_port);
   DataP_IF_IDs_NPC_L_OUT_reg_1_inst : DFFR_X1 port map( D => n1479, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_1_port, QN => n170
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_1_inst : DFFS_X1 port map( D => n170, CK => Clk, 
                           SN => Rst, Q => n169, QN => n_1160);
   DataP_EX_MEM_s_NPC_L_OUT_reg_1_inst : DFFS_X1 port map( D => n169, CK => Clk
                           , SN => Rst, Q => n168, QN => n_1161);
   DataP_MEM_WB_s_NPC_L_OUT_reg_1_inst : DFFS_X1 port map( D => n168, CK => Clk
                           , SN => Rst, Q => n_1162, QN => 
                           DataP_link_addr_W_1_port);
   DataP_IF_IDs_NPC_L_OUT_reg_0_inst : DFFR_X1 port map( D => n1480, CK => Clk,
                           RN => Rst, Q => DataP_link_addr_D_0_port, QN => n167
                           );
   DataP_ID_EXs_NPC_L_OUT_reg_0_inst : DFFS_X1 port map( D => n167, CK => Clk, 
                           SN => Rst, Q => n166, QN => n_1163);
   DataP_EX_MEM_s_NPC_L_OUT_reg_0_inst : DFFS_X1 port map( D => n166, CK => Clk
                           , SN => Rst, Q => n165, QN => n_1164);
   DataP_MEM_WB_s_NPC_L_OUT_reg_0_inst : DFFS_X1 port map( D => n165, CK => Clk
                           , SN => Rst, Q => n_1165, QN => 
                           DataP_link_addr_W_0_port);
   DataP_IF_IDs_NPC_OUT_reg_31_inst : DFFRS_X1 port map( D => DataP_npc_31_port
                           , CK => Clk, RN => n162, SN => n163, Q => n_1166, QN
                           => n164);
   DataP_ID_EXs_NPC_OUT_reg_31_inst : DFFS_X1 port map( D => n164, CK => Clk, 
                           SN => Rst, Q => n161, QN => n_1167);
   DataP_EX_MEM_s_NPC_OUT_reg_31_inst : DFFS_X1 port map( D => n161, CK => Clk,
                           SN => Rst, Q => n_1168, QN => DataP_npc_M_31_port);
   DataP_IF_IDs_NPC_OUT_reg_30_inst : DFFRS_X1 port map( D => DataP_npc_30_port
                           , CK => Clk, RN => n158, SN => n159, Q => n_1169, QN
                           => n160);
   DataP_ID_EXs_NPC_OUT_reg_30_inst : DFFS_X1 port map( D => n160, CK => Clk, 
                           SN => Rst, Q => n157, QN => n_1170);
   DataP_EX_MEM_s_NPC_OUT_reg_30_inst : DFFS_X1 port map( D => n157, CK => Clk,
                           SN => Rst, Q => n_1171, QN => DataP_npc_M_30_port);
   DataP_IF_IDs_NPC_OUT_reg_29_inst : DFFRS_X1 port map( D => DataP_npc_29_port
                           , CK => Clk, RN => n154, SN => n155, Q => n_1172, QN
                           => n156);
   DataP_ID_EXs_NPC_OUT_reg_29_inst : DFFS_X1 port map( D => n156, CK => Clk, 
                           SN => Rst, Q => n153, QN => n_1173);
   DataP_EX_MEM_s_NPC_OUT_reg_29_inst : DFFS_X1 port map( D => n153, CK => Clk,
                           SN => Rst, Q => n_1174, QN => DataP_npc_M_29_port);
   DataP_IF_IDs_NPC_OUT_reg_28_inst : DFFRS_X1 port map( D => DataP_npc_28_port
                           , CK => Clk, RN => n150, SN => n151, Q => n_1175, QN
                           => n152);
   DataP_ID_EXs_NPC_OUT_reg_28_inst : DFFS_X1 port map( D => n152, CK => Clk, 
                           SN => Rst, Q => n149, QN => n_1176);
   DataP_EX_MEM_s_NPC_OUT_reg_28_inst : DFFS_X1 port map( D => n149, CK => Clk,
                           SN => Rst, Q => n_1177, QN => DataP_npc_M_28_port);
   DataP_IF_IDs_NPC_OUT_reg_27_inst : DFFRS_X1 port map( D => DataP_npc_27_port
                           , CK => Clk, RN => n146, SN => n147, Q => n_1178, QN
                           => n148);
   DataP_ID_EXs_NPC_OUT_reg_27_inst : DFFS_X1 port map( D => n148, CK => Clk, 
                           SN => Rst, Q => n145, QN => n_1179);
   DataP_EX_MEM_s_NPC_OUT_reg_27_inst : DFFS_X1 port map( D => n145, CK => Clk,
                           SN => Rst, Q => n_1180, QN => DataP_npc_M_27_port);
   DataP_IF_IDs_NPC_OUT_reg_26_inst : DFFRS_X1 port map( D => DataP_npc_26_port
                           , CK => Clk, RN => n142, SN => n143, Q => n_1181, QN
                           => n144);
   DataP_ID_EXs_NPC_OUT_reg_26_inst : DFFS_X1 port map( D => n144, CK => Clk, 
                           SN => Rst, Q => n141, QN => n_1182);
   DataP_EX_MEM_s_NPC_OUT_reg_26_inst : DFFS_X1 port map( D => n141, CK => Clk,
                           SN => Rst, Q => n_1183, QN => DataP_npc_M_26_port);
   DataP_IF_IDs_NPC_OUT_reg_25_inst : DFFRS_X1 port map( D => DataP_npc_25_port
                           , CK => Clk, RN => n138, SN => n139, Q => n_1184, QN
                           => n140);
   DataP_ID_EXs_NPC_OUT_reg_25_inst : DFFS_X1 port map( D => n140, CK => Clk, 
                           SN => Rst, Q => n137, QN => n_1185);
   DataP_EX_MEM_s_NPC_OUT_reg_25_inst : DFFS_X1 port map( D => n137, CK => Clk,
                           SN => Rst, Q => n_1186, QN => DataP_npc_M_25_port);
   DataP_IF_IDs_NPC_OUT_reg_24_inst : DFFRS_X1 port map( D => DataP_npc_24_port
                           , CK => Clk, RN => n134, SN => n135, Q => n_1187, QN
                           => n136);
   DataP_ID_EXs_NPC_OUT_reg_24_inst : DFFS_X1 port map( D => n136, CK => Clk, 
                           SN => Rst, Q => n133, QN => n_1188);
   DataP_EX_MEM_s_NPC_OUT_reg_24_inst : DFFS_X1 port map( D => n133, CK => Clk,
                           SN => Rst, Q => n_1189, QN => DataP_npc_M_24_port);
   DataP_IF_IDs_NPC_OUT_reg_23_inst : DFFRS_X1 port map( D => DataP_npc_23_port
                           , CK => Clk, RN => n130, SN => n131, Q => n_1190, QN
                           => n132);
   DataP_ID_EXs_NPC_OUT_reg_23_inst : DFFS_X1 port map( D => n132, CK => Clk, 
                           SN => Rst, Q => n129, QN => n_1191);
   DataP_EX_MEM_s_NPC_OUT_reg_23_inst : DFFS_X1 port map( D => n129, CK => Clk,
                           SN => Rst, Q => n_1192, QN => DataP_npc_M_23_port);
   DataP_IF_IDs_NPC_OUT_reg_22_inst : DFFRS_X1 port map( D => DataP_npc_22_port
                           , CK => Clk, RN => n126, SN => n127, Q => n_1193, QN
                           => n128);
   DataP_ID_EXs_NPC_OUT_reg_22_inst : DFFS_X1 port map( D => n128, CK => Clk, 
                           SN => Rst, Q => n125, QN => n_1194);
   DataP_EX_MEM_s_NPC_OUT_reg_22_inst : DFFS_X1 port map( D => n125, CK => Clk,
                           SN => Rst, Q => n_1195, QN => DataP_npc_M_22_port);
   DataP_IF_IDs_NPC_OUT_reg_21_inst : DFFRS_X1 port map( D => DataP_npc_21_port
                           , CK => Clk, RN => n122, SN => n123, Q => n_1196, QN
                           => n124);
   DataP_ID_EXs_NPC_OUT_reg_21_inst : DFFS_X1 port map( D => n124, CK => Clk, 
                           SN => Rst, Q => n121, QN => n_1197);
   DataP_EX_MEM_s_NPC_OUT_reg_21_inst : DFFS_X1 port map( D => n121, CK => Clk,
                           SN => Rst, Q => n_1198, QN => DataP_npc_M_21_port);
   DataP_IF_IDs_NPC_OUT_reg_20_inst : DFFRS_X1 port map( D => DataP_npc_20_port
                           , CK => Clk, RN => n118, SN => n119, Q => n_1199, QN
                           => n120);
   DataP_ID_EXs_NPC_OUT_reg_20_inst : DFFS_X1 port map( D => n120, CK => Clk, 
                           SN => Rst, Q => n117, QN => n_1200);
   DataP_EX_MEM_s_NPC_OUT_reg_20_inst : DFFS_X1 port map( D => n117, CK => Clk,
                           SN => Rst, Q => n_1201, QN => DataP_npc_M_20_port);
   DataP_IF_IDs_NPC_OUT_reg_19_inst : DFFRS_X1 port map( D => DataP_npc_19_port
                           , CK => Clk, RN => n114, SN => n115, Q => n_1202, QN
                           => n116);
   DataP_ID_EXs_NPC_OUT_reg_19_inst : DFFS_X1 port map( D => n116, CK => Clk, 
                           SN => Rst, Q => n113, QN => n_1203);
   DataP_EX_MEM_s_NPC_OUT_reg_19_inst : DFFS_X1 port map( D => n113, CK => Clk,
                           SN => Rst, Q => n_1204, QN => DataP_npc_M_19_port);
   DataP_IF_IDs_NPC_OUT_reg_18_inst : DFFRS_X1 port map( D => DataP_npc_18_port
                           , CK => Clk, RN => n110, SN => n111, Q => n_1205, QN
                           => n112);
   DataP_ID_EXs_NPC_OUT_reg_18_inst : DFFS_X1 port map( D => n112, CK => Clk, 
                           SN => Rst, Q => n109, QN => n_1206);
   DataP_EX_MEM_s_NPC_OUT_reg_18_inst : DFFS_X1 port map( D => n109, CK => Clk,
                           SN => Rst, Q => n_1207, QN => DataP_npc_M_18_port);
   DataP_IF_IDs_NPC_OUT_reg_17_inst : DFFRS_X1 port map( D => DataP_npc_17_port
                           , CK => Clk, RN => n106, SN => n107, Q => n_1208, QN
                           => n108);
   DataP_ID_EXs_NPC_OUT_reg_17_inst : DFFS_X1 port map( D => n108, CK => Clk, 
                           SN => Rst, Q => n105, QN => n1606);
   DataP_EX_MEM_s_NPC_OUT_reg_17_inst : DFFS_X1 port map( D => n105, CK => Clk,
                           SN => Rst, Q => n_1209, QN => DataP_npc_M_17_port);
   DataP_IF_IDs_NPC_OUT_reg_16_inst : DFFRS_X1 port map( D => DataP_npc_16_port
                           , CK => Clk, RN => n102, SN => n103, Q => n_1210, QN
                           => n104);
   DataP_ID_EXs_NPC_OUT_reg_16_inst : DFFS_X1 port map( D => n104, CK => Clk, 
                           SN => Rst, Q => n101, QN => n_1211);
   DataP_EX_MEM_s_NPC_OUT_reg_16_inst : DFFS_X1 port map( D => n101, CK => Clk,
                           SN => Rst, Q => n_1212, QN => DataP_npc_M_16_port);
   DataP_IF_IDs_NPC_OUT_reg_15_inst : DFFRS_X1 port map( D => DataP_npc_15_port
                           , CK => Clk, RN => n98, SN => n99, Q => n_1213, QN 
                           => n100);
   DataP_ID_EXs_NPC_OUT_reg_15_inst : DFFS_X1 port map( D => n100, CK => Clk, 
                           SN => Rst, Q => n97, QN => n_1214);
   DataP_EX_MEM_s_NPC_OUT_reg_15_inst : DFFS_X1 port map( D => n97, CK => Clk, 
                           SN => Rst, Q => n_1215, QN => DataP_npc_M_15_port);
   DataP_IF_IDs_NPC_OUT_reg_14_inst : DFFRS_X1 port map( D => DataP_npc_14_port
                           , CK => Clk, RN => n94, SN => n95, Q => n_1216, QN 
                           => n96);
   DataP_ID_EXs_NPC_OUT_reg_14_inst : DFFS_X1 port map( D => n96, CK => Clk, SN
                           => Rst, Q => n93, QN => n_1217);
   DataP_EX_MEM_s_NPC_OUT_reg_14_inst : DFFS_X1 port map( D => n93, CK => Clk, 
                           SN => Rst, Q => n_1218, QN => DataP_npc_M_14_port);
   DataP_IF_IDs_NPC_OUT_reg_13_inst : DFFRS_X1 port map( D => DataP_npc_13_port
                           , CK => Clk, RN => n90, SN => n91, Q => n_1219, QN 
                           => n92);
   DataP_ID_EXs_NPC_OUT_reg_13_inst : DFFS_X1 port map( D => n92, CK => Clk, SN
                           => Rst, Q => n89, QN => n_1220);
   DataP_EX_MEM_s_NPC_OUT_reg_13_inst : DFFS_X1 port map( D => n89, CK => Clk, 
                           SN => Rst, Q => n_1221, QN => DataP_npc_M_13_port);
   DataP_IF_IDs_NPC_OUT_reg_12_inst : DFFRS_X1 port map( D => DataP_npc_12_port
                           , CK => Clk, RN => n86, SN => n87, Q => n_1222, QN 
                           => n88);
   DataP_ID_EXs_NPC_OUT_reg_12_inst : DFFS_X1 port map( D => n88, CK => Clk, SN
                           => Rst, Q => n85, QN => n1969);
   DataP_EX_MEM_s_NPC_OUT_reg_12_inst : DFFS_X1 port map( D => n85, CK => Clk, 
                           SN => Rst, Q => n_1223, QN => DataP_npc_M_12_port);
   DataP_IF_IDs_NPC_OUT_reg_11_inst : DFFRS_X1 port map( D => DataP_npc_11_port
                           , CK => Clk, RN => n82, SN => n83, Q => n_1224, QN 
                           => n84);
   DataP_ID_EXs_NPC_OUT_reg_11_inst : DFFS_X1 port map( D => n84, CK => Clk, SN
                           => Rst, Q => n81, QN => n_1225);
   DataP_EX_MEM_s_NPC_OUT_reg_11_inst : DFFS_X1 port map( D => n81, CK => Clk, 
                           SN => Rst, Q => n_1226, QN => DataP_npc_M_11_port);
   DataP_IF_IDs_NPC_OUT_reg_10_inst : DFFRS_X1 port map( D => DataP_npc_10_port
                           , CK => Clk, RN => n78, SN => n79, Q => n_1227, QN 
                           => n80);
   DataP_ID_EXs_NPC_OUT_reg_10_inst : DFFS_X1 port map( D => n80, CK => Clk, SN
                           => Rst, Q => n77, QN => n_1228);
   DataP_EX_MEM_s_NPC_OUT_reg_10_inst : DFFS_X1 port map( D => n77, CK => Clk, 
                           SN => Rst, Q => n_1229, QN => DataP_npc_M_10_port);
   DataP_IF_IDs_NPC_OUT_reg_9_inst : DFFRS_X1 port map( D => DataP_npc_9_port, 
                           CK => Clk, RN => n74, SN => n75, Q => n_1230, QN => 
                           n76);
   DataP_ID_EXs_NPC_OUT_reg_9_inst : DFFS_X1 port map( D => n76, CK => Clk, SN 
                           => Rst, Q => n73, QN => DataP_npc_E_9_port);
   DataP_EX_MEM_s_NPC_OUT_reg_9_inst : DFFS_X1 port map( D => n73, CK => Clk, 
                           SN => Rst, Q => n_1231, QN => DataP_npc_M_9_port);
   DataP_IF_IDs_NPC_OUT_reg_8_inst : DFFRS_X1 port map( D => DataP_npc_8_port, 
                           CK => Clk, RN => n70, SN => n71, Q => n_1232, QN => 
                           n72);
   DataP_ID_EXs_NPC_OUT_reg_8_inst : DFFS_X1 port map( D => n72, CK => Clk, SN 
                           => Rst, Q => n69, QN => n_1233);
   DataP_EX_MEM_s_NPC_OUT_reg_8_inst : DFFS_X1 port map( D => n69, CK => Clk, 
                           SN => Rst, Q => n_1234, QN => DataP_npc_M_8_port);
   DataP_IF_IDs_NPC_OUT_reg_7_inst : DFFRS_X1 port map( D => DataP_npc_7_port, 
                           CK => Clk, RN => n66, SN => n67, Q => n_1235, QN => 
                           n68);
   DataP_ID_EXs_NPC_OUT_reg_7_inst : DFFS_X1 port map( D => n68, CK => Clk, SN 
                           => Rst, Q => n65, QN => n_1236);
   DataP_EX_MEM_s_NPC_OUT_reg_7_inst : DFFS_X1 port map( D => n65, CK => Clk, 
                           SN => Rst, Q => n_1237, QN => DataP_npc_M_7_port);
   DataP_IF_IDs_NPC_OUT_reg_6_inst : DFFRS_X1 port map( D => DataP_npc_6_port, 
                           CK => Clk, RN => n62, SN => n63, Q => n_1238, QN => 
                           n64);
   DataP_ID_EXs_NPC_OUT_reg_6_inst : DFFS_X1 port map( D => n64, CK => Clk, SN 
                           => Rst, Q => n61, QN => n_1239);
   DataP_EX_MEM_s_NPC_OUT_reg_6_inst : DFFS_X1 port map( D => n61, CK => Clk, 
                           SN => Rst, Q => n_1240, QN => DataP_npc_M_6_port);
   DataP_IF_IDs_NPC_OUT_reg_5_inst : DFFRS_X1 port map( D => DataP_npc_5_port, 
                           CK => Clk, RN => n58, SN => n59, Q => n_1241, QN => 
                           n60);
   DataP_ID_EXs_NPC_OUT_reg_5_inst : DFFS_X1 port map( D => n60, CK => Clk, SN 
                           => Rst, Q => n57, QN => n_1242);
   DataP_EX_MEM_s_NPC_OUT_reg_5_inst : DFFS_X1 port map( D => n57, CK => Clk, 
                           SN => Rst, Q => n_1243, QN => DataP_npc_M_5_port);
   DataP_IF_IDs_NPC_OUT_reg_4_inst : DFFRS_X1 port map( D => DataP_npc_4_port, 
                           CK => Clk, RN => n54, SN => n55, Q => n_1244, QN => 
                           n56);
   DataP_ID_EXs_NPC_OUT_reg_4_inst : DFFS_X1 port map( D => n56, CK => Clk, SN 
                           => Rst, Q => n53, QN => n_1245);
   DataP_EX_MEM_s_NPC_OUT_reg_4_inst : DFFS_X1 port map( D => n53, CK => Clk, 
                           SN => Rst, Q => n_1246, QN => DataP_npc_M_4_port);
   DataP_IF_IDs_NPC_OUT_reg_3_inst : DFFRS_X1 port map( D => DataP_npc_3_port, 
                           CK => Clk, RN => n50, SN => n51, Q => n_1247, QN => 
                           n52);
   DataP_ID_EXs_NPC_OUT_reg_3_inst : DFFS_X1 port map( D => n52, CK => Clk, SN 
                           => Rst, Q => n49, QN => n_1248);
   DataP_EX_MEM_s_NPC_OUT_reg_3_inst : DFFS_X1 port map( D => n49, CK => Clk, 
                           SN => Rst, Q => n_1249, QN => DataP_npc_M_3_port);
   DataP_IF_IDs_NPC_OUT_reg_2_inst : DFFRS_X1 port map( D => DataP_npc_2_port, 
                           CK => Clk, RN => n46, SN => n47, Q => n_1250, QN => 
                           n48);
   DataP_ID_EXs_NPC_OUT_reg_2_inst : DFFS_X1 port map( D => n48, CK => Clk, SN 
                           => Rst, Q => n45, QN => n_1251);
   DataP_EX_MEM_s_NPC_OUT_reg_2_inst : DFFS_X1 port map( D => n45, CK => Clk, 
                           SN => Rst, Q => n_1252, QN => DataP_npc_M_2_port);
   DataP_IF_IDs_NPC_OUT_reg_1_inst : DFFRS_X1 port map( D => DataP_npc_1_port, 
                           CK => Clk, RN => n42, SN => n43, Q => n_1253, QN => 
                           n44);
   DataP_ID_EXs_NPC_OUT_reg_1_inst : DFFS_X1 port map( D => n44, CK => Clk, SN 
                           => Rst, Q => n41, QN => n_1254);
   DataP_EX_MEM_s_NPC_OUT_reg_1_inst : DFFS_X1 port map( D => n41, CK => Clk, 
                           SN => Rst, Q => n_1255, QN => DataP_npc_M_1_port);
   DataP_IF_IDs_NPC_OUT_reg_0_inst : DFFRS_X1 port map( D => DataP_npc_0_port, 
                           CK => Clk, RN => n38, SN => n39, Q => n_1256, QN => 
                           n40);
   DataP_ID_EXs_NPC_OUT_reg_0_inst : DFFS_X1 port map( D => n40, CK => Clk, SN 
                           => Rst, Q => n37, QN => n_1257);
   DataP_EX_MEM_s_NPC_OUT_reg_0_inst : DFFS_X1 port map( D => n37, CK => Clk, 
                           SN => Rst, Q => n_1258, QN => DataP_npc_M_0_port);
   DataP_IF_IDs_IR_OUT_reg_0_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(0), CK
                           => Clk, RN => n36, Q => IR_CU_0_port, QN => n476);
   DataP_ID_EXs_IMM_OUT_reg_0_inst : DFFS_X1 port map( D => n476, CK => Clk, SN
                           => Rst, Q => n_1259, QN => DataP_IMM_s_0_port);
   DataP_IF_IDs_IR_OUT_reg_1_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(1), CK
                           => Clk, RN => n36, Q => IR_CU_1_port, QN => n477);
   DataP_ID_EXs_IMM_OUT_reg_1_inst : DFFS_X1 port map( D => n477, CK => Clk, SN
                           => Rst, Q => n_1260, QN => DataP_IMM_s_1_port);
   DataP_IF_IDs_IR_OUT_reg_2_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(2), CK
                           => Clk, RN => n36, Q => n2375, QN => n478);
   DataP_ID_EXs_IMM_OUT_reg_2_inst : DFFS_X1 port map( D => n478, CK => Clk, SN
                           => Rst, Q => n_1261, QN => DataP_IMM_s_2_port);
   DataP_IF_IDs_IR_OUT_reg_3_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(3), CK
                           => Clk, RN => n36, Q => n2399, QN => n479);
   DataP_ID_EXs_IMM_OUT_reg_3_inst : DFFS_X1 port map( D => n479, CK => Clk, SN
                           => Rst, Q => n_1262, QN => DataP_IMM_s_3_port);
   DataP_IF_IDs_IR_OUT_reg_4_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(4), CK
                           => Clk, RN => n36, Q => IR_CU_4_port, QN => n480);
   DataP_ID_EXs_IMM_OUT_reg_4_inst : DFFS_X1 port map( D => n480, CK => Clk, SN
                           => Rst, Q => n_1263, QN => DataP_IMM_s_4_port);
   DataP_IF_IDs_IR_OUT_reg_5_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(5), CK
                           => Clk, RN => n36, Q => IR_CU_5_port, QN => n482);
   DataP_ID_EXs_IMM_OUT_reg_5_inst : DFFS_X1 port map( D => n482, CK => Clk, SN
                           => Rst, Q => n_1264, QN => DataP_IMM_s_5_port);
   DataP_IF_IDs_IR_OUT_reg_6_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(6), CK
                           => Clk, RN => n36, Q => IR_CU_6_port, QN => n35);
   DataP_ID_EXs_IMM_OUT_reg_6_inst : DFFS_X1 port map( D => n35, CK => Clk, SN 
                           => Rst, Q => n_1265, QN => DataP_IMM_s_6_port);
   DataP_IF_IDs_IR_OUT_reg_7_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(7), CK
                           => Clk, RN => n36, Q => IR_CU_7_port, QN => n34);
   DataP_ID_EXs_IMM_OUT_reg_7_inst : DFFS_X1 port map( D => n34, CK => Clk, SN 
                           => Rst, Q => n_1266, QN => DataP_IMM_s_7_port);
   DataP_IF_IDs_IR_OUT_reg_8_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(8), CK
                           => Clk, RN => n36, Q => IR_CU_8_port, QN => n33);
   DataP_ID_EXs_IMM_OUT_reg_8_inst : DFFS_X1 port map( D => n33, CK => Clk, SN 
                           => Rst, Q => n_1267, QN => DataP_IMM_s_8_port);
   DataP_IF_IDs_IR_OUT_reg_9_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(9), CK
                           => Clk, RN => n36, Q => IR_CU_9_port, QN => n32);
   DataP_ID_EXs_IMM_OUT_reg_9_inst : DFFS_X1 port map( D => n32, CK => Clk, SN 
                           => Rst, Q => n_1268, QN => DataP_IMM_s_9_port);
   DataP_IF_IDs_IR_OUT_reg_10_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(10), 
                           CK => Clk, RN => n36, Q => n_1269, QN => n484);
   DataP_ID_EXs_IMM_OUT_reg_10_inst : DFFS_X1 port map( D => n484, CK => Clk, 
                           SN => Rst, Q => n_1270, QN => DataP_IMM_s_10_port);
   DataP_IF_IDs_IR_OUT_reg_11_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(11), 
                           CK => Clk, RN => n36, Q => DataP_IR1_11_port, QN => 
                           n31);
   DataP_ID_EXs_IMM_OUT_reg_11_inst : DFFS_X1 port map( D => n31, CK => Clk, SN
                           => Rst, Q => n_1271, QN => DataP_IMM_s_11_port);
   DataP_IF_IDs_IR_OUT_reg_12_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(12), 
                           CK => Clk, RN => n36, Q => DataP_IR1_12_port, QN => 
                           n30);
   DataP_ID_EXs_IMM_OUT_reg_12_inst : DFFS_X1 port map( D => n30, CK => Clk, SN
                           => Rst, Q => n_1272, QN => DataP_IMM_s_12_port);
   DataP_IF_IDs_IR_OUT_reg_13_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(13), 
                           CK => Clk, RN => n36, Q => DataP_IR1_13_port, QN => 
                           n29);
   DataP_ID_EXs_IMM_OUT_reg_13_inst : DFFS_X1 port map( D => n29, CK => Clk, SN
                           => Rst, Q => n_1273, QN => DataP_IMM_s_13_port);
   DataP_IF_IDs_IR_OUT_reg_14_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(14), 
                           CK => Clk, RN => n36, Q => DataP_IR1_14_port, QN => 
                           n28);
   DataP_ID_EXs_IMM_OUT_reg_14_inst : DFFS_X1 port map( D => n28, CK => Clk, SN
                           => Rst, Q => n_1274, QN => DataP_IMM_s_14_port);
   DataP_IF_IDs_IR_OUT_reg_15_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(15), 
                           CK => Clk, RN => n36, Q => DataP_IR1_15_port, QN => 
                           n27);
   DataP_ID_EXs_IMM_OUT_reg_15_inst : DFFS_X1 port map( D => n27, CK => Clk, SN
                           => Rst, Q => n_1275, QN => DataP_IMM_s_15_port);
   DataP_IF_IDs_IR_OUT_reg_16_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(16), 
                           CK => Clk, RN => n36, Q => n_1276, QN => n485);
   DataP_IF_IDs_IR_OUT_reg_17_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(17), 
                           CK => Clk, RN => n36, Q => n_1277, QN => n486);
   DataP_IF_IDs_IR_OUT_reg_18_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(18), 
                           CK => Clk, RN => n36, Q => n_1278, QN => n487);
   DataP_IF_IDs_IR_OUT_reg_19_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(19), 
                           CK => Clk, RN => n36, Q => n_1279, QN => n488);
   DataP_IF_IDs_IR_OUT_reg_20_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(20), 
                           CK => Clk, RN => n36, Q => n_1280, QN => n489);
   DataP_IF_IDs_IR_OUT_reg_21_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(21), 
                           CK => Clk, RN => n36, Q => DataP_IR1_21_port, QN => 
                           n26);
   DataP_ID_EXs_RS1_OUT_reg_0_inst : DFFS_X1 port map( D => n26, CK => Clk, SN 
                           => Rst, Q => n2392, QN => n_1281);
   DataP_IF_IDs_IR_OUT_reg_22_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(22), 
                           CK => Clk, RN => n36, Q => DataP_IR1_22_port, QN => 
                           n25);
   DataP_ID_EXs_RS1_OUT_reg_1_inst : DFFS_X1 port map( D => n25, CK => Clk, SN 
                           => Rst, Q => n2429, QN => DataP_Rs1_1_port);
   DataP_IF_IDs_IR_OUT_reg_23_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(23), 
                           CK => Clk, RN => n36, Q => DataP_IR1_23_port, QN => 
                           n24);
   DataP_ID_EXs_RS1_OUT_reg_2_inst : DFFS_X1 port map( D => n24, CK => Clk, SN 
                           => Rst, Q => n2407, QN => DataP_Rs1_2_port);
   DataP_IF_IDs_IR_OUT_reg_24_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(24), 
                           CK => Clk, RN => n36, Q => DataP_IR1_24_port, QN => 
                           n_1282);
   DataP_ID_EXs_RS1_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_IR1_24_port, 
                           CK => Clk, RN => Rst, Q => n_1283, QN => n523);
   DataP_IF_IDs_IR_OUT_reg_25_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(25), 
                           CK => Clk, RN => n36, Q => DataP_IR1_25_port, QN => 
                           n_1284);
   DataP_ID_EXs_RS1_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_IR1_25_port, 
                           CK => Clk, RN => Rst, Q => n_1285, QN => n524);
   DataP_IF_IDs_IR_OUT_reg_26_inst : DFFS_X1 port map( D => IRAM_DATA_OUT(26), 
                           CK => Clk, SN => n36, Q => IR_CU_26, QN => n497);
   DataP_ID_EXs_OPCODE_OUT_reg_0_inst : DFFS_X1 port map( D => n497, CK => Clk,
                           SN => Rst, Q => n23, QN => DataP_opcode_E_0_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_0_inst : DFFS_X1 port map( D => n23, CK => Clk
                           , SN => Rst, Q => n22, QN => DataP_opcode_M_0_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_0_inst : DFFS_X1 port map( D => n22, CK => Clk
                           , SN => Rst, Q => n2403, QN => DataP_opcode_W_0_port
                           );
   DataP_ID_EXs_OPCODE_OUT_reg_1_inst : DFFS_X1 port map( D => n504, CK => Clk,
                           SN => Rst, Q => n520, QN => DataP_opcode_E_1_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_1_inst : DFFS_X1 port map( D => n520, CK => 
                           Clk, SN => Rst, Q => n2249, QN => 
                           DataP_opcode_M_1_port);
   DataP_IF_IDs_IR_OUT_reg_28_inst : DFFS_X1 port map( D => IRAM_DATA_OUT(28), 
                           CK => Clk, SN => n36, Q => IR_CU_28, QN => n1960);
   DataP_IF_IDs_IR_OUT_reg_29_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(29), 
                           CK => Clk, RN => n36, Q => n2374, QN => n514);
   DataP_ID_EXs_OPCODE_OUT_reg_3_inst : DFFS_X1 port map( D => n514, CK => Clk,
                           SN => Rst, Q => n21, QN => DataP_opcode_E_3_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_3_inst : DFFS_X1 port map( D => n21, CK => Clk
                           , SN => Rst, Q => n20, QN => DataP_opcode_M_3_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_3_inst : DFFS_X1 port map( D => n20, CK => Clk
                           , SN => Rst, Q => n2401, QN => DataP_opcode_W_3_port
                           );
   DataP_ID_EXs_OPCODE_OUT_reg_4_inst : DFFS_X1 port map( D => n515, CK => Clk,
                           SN => Rst, Q => n19, QN => DataP_opcode_E_4_port);
   DataP_EX_MEM_s_OPCODE_OUT_reg_4_inst : DFFS_X1 port map( D => n19, CK => Clk
                           , SN => Rst, Q => n18, QN => DataP_opcode_M_4_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_4_inst : DFFS_X1 port map( D => n18, CK => Clk
                           , SN => Rst, Q => n2383, QN => DataP_opcode_W_4_port
                           );
   DataP_IF_IDs_IR_OUT_reg_31_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(31), 
                           CK => Clk, RN => n36, Q => IR_CU_31, QN => n516);
   DataP_EX_MEM_s_OPCODE_OUT_reg_5_inst : DFFS_X1 port map( D => n17, CK => Clk
                           , SN => Rst, Q => n2387, QN => n_1286);
   DataP_FORWARDING_BR_SEL_reg_1_inst : DLH_X1 port map( G => 
                           DataP_FORWARDING_BR_N12, D => n3910, Q => 
                           DataP_FWD_MUX_BR_S_1_port);
   CU_I_cw1_reg_8_inst : SDFFR_X1 port map( D => n16, SI => n607, SE => n504, 
                           CK => Clk, RN => Rst, Q => BR_EN_i, QN => n_1287);
   CU_I_cw1_reg_7_inst : DFFR_X1 port map( D => CU_I_cw_7_port, CK => Clk, RN 
                           => Rst, Q => n_1288, QN => n15);
   CU_I_cw2_reg_7_inst : DFFS_X1 port map( D => n15, CK => Clk, SN => Rst, Q =>
                           n_1289, QN => DRAM_RW);
   DataP_ID_EXs_RD_OUT_reg_4_inst : DFFR_X1 port map( D => DataP_dest_D_4_port,
                           CK => Clk, RN => Rst, Q => n_1290, QN => n14);
   DataP_ID_EXs_RD_OUT_reg_3_inst : DFFR_X1 port map( D => DataP_dest_D_3_port,
                           CK => Clk, RN => Rst, Q => n_1291, QN => n13);
   DataP_ID_EXs_RD_OUT_reg_2_inst : DFFR_X1 port map( D => DataP_dest_D_2_port,
                           CK => Clk, RN => Rst, Q => n_1292, QN => n12);
   DataP_EX_MEM_s_RD_OUT_reg_2_inst : DFFS_X1 port map( D => n12, CK => Clk, SN
                           => Rst, Q => n530, QN => DataP_dest_M_2_port);
   DataP_MEM_WB_s_RD_OUT_reg_2_inst : DFFR_X1 port map( D => 
                           DataP_dest_M_2_port, CK => Clk, RN => Rst, Q => 
                           DataP_add_D_2_port, QN => n538);
   DataP_ID_EXs_RD_OUT_reg_1_inst : DFFR_X1 port map( D => DataP_dest_D_1_port,
                           CK => Clk, RN => Rst, Q => n_1293, QN => n11);
   DataP_ID_EXs_RD_OUT_reg_0_inst : DFFR_X1 port map( D => DataP_dest_D_0_port,
                           CK => Clk, RN => Rst, Q => n_1294, QN => n10);
   DataP_EX_MEM_s_RD_OUT_reg_0_inst : DFFS_X1 port map( D => n10, CK => Clk, SN
                           => Rst, Q => n528, QN => DataP_dest_M_0_port);
   DataP_MEM_WB_s_RD_OUT_reg_0_inst : DFFR_X1 port map( D => 
                           DataP_dest_M_0_port, CK => Clk, RN => Rst, Q => 
                           DataP_add_D_0_port, QN => n536);
   DataP_FORWARDING_BR_SEL_reg_0_inst : DLH_X1 port map( G => 
                           DataP_FORWARDING_BR_N12, D => n3909, Q => 
                           DataP_FWD_MUX_BR_S_0_port);
   CU_I_aluOpcode1_reg_2_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_2_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_2_port, QN 
                           => n2391);
   CU_I_cw1_reg_5_inst : DFFS_X1 port map( D => n1358, CK => Clk, SN => Rst, Q 
                           => n9, QN => n_1295);
   CU_I_cw2_reg_5_inst : DFFS_X1 port map( D => n9, CK => Clk, SN => Rst, Q => 
                           n_1296, QN => DRAM_SEL(2));
   CU_I_cw1_reg_0_inst : DFFR_X1 port map( D => CU_I_cw_0_port, CK => Clk, RN 
                           => Rst, Q => n_1297, QN => n8);
   CU_I_cw2_reg_0_inst : DFFS_X1 port map( D => n8, CK => Clk, SN => Rst, Q => 
                           n7, QN => n_1298);
   CU_I_cw3_reg_0_inst : DFFS_X1 port map( D => n7, CK => Clk, SN => Rst, Q => 
                           n_1299, QN => RF_WE_i);
   CU_I_cw1_reg_2_inst : DFFS_X1 port map( D => n1372, CK => Clk, SN => Rst, Q 
                           => n6, QN => n_1300);
   CU_I_cw2_reg_2_inst : DFFS_X1 port map( D => n6, CK => Clk, SN => Rst, Q => 
                           n5, QN => n_1301);
   CU_I_cw3_reg_2_inst : DFFS_X1 port map( D => n5, CK => Clk, SN => Rst, Q => 
                           n_1302, QN => WB_MUX_SEL_i_1_port);
   CU_I_cw1_reg_4_inst : DFFR_X1 port map( D => CU_I_cw_4_port, CK => Clk, RN 
                           => Rst, Q => n_1303, QN => n4);
   CU_I_cw2_reg_4_inst : DFFS_X1 port map( D => n4, CK => Clk, SN => Rst, Q => 
                           n_1304, QN => DRAM_SEL(1));
   CU_I_cw1_reg_3_inst : DFFR_X1 port map( D => CU_I_cw_3_port, CK => Clk, RN 
                           => Rst, Q => n_1305, QN => n3);
   CU_I_cw2_reg_3_inst : DFFS_X1 port map( D => n3, CK => Clk, SN => Rst, Q => 
                           n_1306, QN => DRAM_SEL(0));
   CU_I_cw1_reg_6_inst : DFFR_X1 port map( D => CU_I_cw_6_port, CK => Clk, RN 
                           => Rst, Q => n_1307, QN => n2);
   CU_I_cw2_reg_6_inst : DFFS_X1 port map( D => n2, CK => Clk, SN => Rst, Q => 
                           n_1308, QN => DRAM_ENABLE);
   DataP_EX_MEM_s_ALU_OUT_reg_12_inst : DFFS_X1 port map( D => n337, CK => Clk,
                           SN => Rst, Q => n2424, QN => DataP_alu_out_M_12_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_13_inst : DFFS_X1 port map( D => n333, CK => Clk,
                           SN => Rst, Q => n2423, QN => DataP_alu_out_M_13_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_14_inst : DFFS_X1 port map( D => n332, CK => Clk,
                           SN => Rst, Q => n2418, QN => DataP_alu_out_M_14_port
                           );
   DataP_PC_reg_O_reg_14_inst : DFF_X1 port map( D => DataP_PC_reg_N16, CK => 
                           Clk, Q => DataP_pc_out_14_port, QN => n_1309);
   DataP_PC_reg_O_reg_13_inst : DFF_X1 port map( D => DataP_PC_reg_N15, CK => 
                           Clk, Q => DataP_pc_out_13_port, QN => n_1310);
   DataP_PC_reg_O_reg_12_inst : DFF_X1 port map( D => DataP_PC_reg_N14, CK => 
                           Clk, Q => DataP_pc_out_12_port, QN => n_1311);
   DataP_EX_MEM_s_ALU_OUT_reg_4_inst : DFFS_X1 port map( D => n355, CK => Clk, 
                           SN => Rst, Q => n2466, QN => DRAM_ADDRESS_4_port);
   DataP_EX_MEM_s_ALU_OUT_reg_5_inst : DFFS_X1 port map( D => n354, CK => Clk, 
                           SN => Rst, Q => n2450, QN => DRAM_ADDRESS_5_port);
   DataP_EX_MEM_s_ALU_OUT_reg_6_inst : DFFS_X1 port map( D => n353, CK => Clk, 
                           SN => Rst, Q => n2410, QN => DRAM_ADDRESS_6_port);
   DataP_PC_reg_O_reg_6_inst : DFF_X1 port map( D => DataP_PC_reg_N8, CK => Clk
                           , Q => IRAM_ADDRESS_4_port, QN => n_1312);
   DataP_PC_reg_O_reg_5_inst : DFF_X1 port map( D => DataP_PC_reg_N7, CK => Clk
                           , Q => IRAM_ADDRESS_3_port, QN => n_1313);
   DataP_PC_reg_O_reg_4_inst : DFF_X1 port map( D => DataP_PC_reg_N6, CK => Clk
                           , Q => IRAM_ADDRESS_2_port, QN => n_1314);
   DataP_EX_MEM_s_ALU_OUT_reg_1_inst : DFFS_X1 port map( D => n358, CK => Clk, 
                           SN => Rst, Q => n2469, QN => DRAM_ADDRESS_1_port);
   DataP_PC_reg_O_reg_1_inst : DFF_X1 port map( D => DataP_PC_reg_N3, CK => Clk
                           , Q => DataP_pc_out_1, QN => n_1315);
   DataP_EX_MEM_s_ALU_OUT_reg_2_inst : DFFS_X1 port map( D => n357, CK => Clk, 
                           SN => Rst, Q => n2471, QN => DRAM_ADDRESS_2_port);
   DataP_PC_reg_O_reg_2_inst : DFF_X1 port map( D => DataP_PC_reg_N4, CK => Clk
                           , Q => IRAM_ADDRESS_0_port, QN => n_1316);
   DataP_EX_MEM_s_ALU_OUT_reg_3_inst : DFFS_X1 port map( D => n356, CK => Clk, 
                           SN => Rst, Q => n2478, QN => DRAM_ADDRESS_3_port);
   DataP_PC_reg_O_reg_3_inst : DFF_X1 port map( D => DataP_PC_reg_N5, CK => Clk
                           , Q => IRAM_ADDRESS_1_port, QN => n_1317);
   DataP_EX_MEM_s_ALU_OUT_reg_8_inst : DFFS_X1 port map( D => n345, CK => Clk, 
                           SN => Rst, Q => n2408, QN => DRAM_ADDRESS_8_port);
   DataP_EX_MEM_s_ALU_OUT_reg_9_inst : DFFS_X1 port map( D => n341, CK => Clk, 
                           SN => Rst, Q => n2477, QN => DRAM_ADDRESS_9_port);
   DataP_EX_MEM_s_ALU_OUT_reg_10_inst : DFFS_X1 port map( D => n340, CK => Clk,
                           SN => Rst, Q => n2409, QN => DRAM_ADDRESS_10_port);
   DataP_PC_reg_O_reg_10_inst : DFF_X1 port map( D => DataP_PC_reg_N12, CK => 
                           Clk, Q => DataP_pc_out_10_port, QN => n_1318);
   DataP_EX_MEM_s_ALU_OUT_reg_11_inst : DFFS_X1 port map( D => n2386, CK => Clk
                           , SN => Rst, Q => n2431, QN => DRAM_ADDRESS_11_port)
                           ;
   DataP_PC_reg_O_reg_9_inst : DFF_X1 port map( D => DataP_PC_reg_N11, CK => 
                           Clk, Q => IRAM_ADDRESS_7_port, QN => n_1319);
   DataP_PC_reg_O_reg_8_inst : DFF_X1 port map( D => DataP_PC_reg_N10, CK => 
                           Clk, Q => IRAM_ADDRESS_6_port, QN => n_1320);
   CU_I_cw1_reg_1_inst : DFFR_X1 port map( D => CU_I_cw_1_port, CK => Clk, RN 
                           => Rst, Q => n_1321, QN => n1);
   CU_I_cw2_reg_1_inst : DFFS_X1 port map( D => n1, CK => Clk, SN => Rst, Q => 
                           n_1322, QN => CU_I_cw2_1_port);
   CU_I_cw3_reg_1_inst : DFFR_X1 port map( D => CU_I_cw2_1_port, CK => Clk, RN 
                           => Rst, Q => n_1323, QN => n294);
   DataP_EX_MEM_s_ALU_OUT_reg_28_inst : DFFS_X1 port map( D => n300, CK => Clk,
                           SN => Rst, Q => n2426, QN => DataP_alu_out_M_28_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_24_inst : DFFS_X1 port map( D => n1759, CK => Clk
                           , SN => Rst, Q => n2427, QN => 
                           DataP_alu_out_M_24_port);
   DataP_EX_MEM_s_ALU_OUT_reg_25_inst : DFFS_X1 port map( D => n1624, CK => Clk
                           , SN => Rst, Q => n2422, QN => 
                           DataP_alu_out_M_25_port);
   DataP_EX_MEM_s_ALU_OUT_reg_20_inst : DFFS_X1 port map( D => n317, CK => Clk,
                           SN => Rst, Q => n2420, QN => DataP_alu_out_M_20_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_21_inst : DFFS_X1 port map( D => n313, CK => Clk,
                           SN => Rst, Q => n2419, QN => DataP_alu_out_M_21_port
                           );
   DataP_PC_reg_O_reg_22_inst : DFF_X1 port map( D => DataP_PC_reg_N24, CK => 
                           Clk, Q => DataP_pc_out_22_port, QN => n_1324);
   DataP_EX_MEM_s_ALU_OUT_reg_16_inst : DFFS_X1 port map( D => n326, CK => Clk,
                           SN => Rst, Q => n2412, QN => DataP_alu_out_M_16_port
                           );
   DataP_EX_MEM_s_ALU_OUT_reg_18_inst : DFFS_X1 port map( D => n322, CK => Clk,
                           SN => Rst, Q => n2425, QN => DataP_alu_out_M_18_port
                           );
   DataP_PC_reg_O_reg_18_inst : DFF_X1 port map( D => DataP_PC_reg_N20, CK => 
                           Clk, Q => DataP_pc_out_18_port, QN => n_1325);
   DataP_PC_reg_O_reg_16_inst : DFF_X1 port map( D => DataP_PC_reg_N18, CK => 
                           Clk, Q => DataP_pc_out_16_port, QN => n_1326);
   DataP_PC_reg_O_reg_27_inst : DFF_X1 port map( D => DataP_PC_reg_N29, CK => 
                           Clk, Q => DataP_pc_out_27_port, QN => n_1327);
   DataP_PC_reg_O_reg_23_inst : DFF_X1 port map( D => DataP_PC_reg_N25, CK => 
                           Clk, Q => DataP_pc_out_23_port, QN => n_1328);
   DataP_PC_reg_O_reg_19_inst : DFF_X1 port map( D => DataP_PC_reg_N21, CK => 
                           Clk, Q => DataP_pc_out_19_port, QN => n_1329);
   DataP_PC_reg_O_reg_7_inst : DFF_X1 port map( D => DataP_PC_reg_N9, CK => Clk
                           , Q => IRAM_ADDRESS_5_port, QN => n_1330);
   DataP_EX_MEM_s_RD_OUT_reg_4_inst : DFFS_X1 port map( D => n14, CK => Clk, SN
                           => Rst, Q => n2778, QN => DataP_dest_M_4_port);
   DataP_EX_MEM_s_RD_OUT_reg_3_inst : DFFS_X1 port map( D => n13, CK => Clk, SN
                           => Rst, Q => n2777, QN => DataP_dest_M_3_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_5_inst : DFFS_X1 port map( D => n2387, CK => 
                           Clk, SN => Rst, Q => n3264, QN => 
                           DataP_opcode_W_5_port);
   DataP_ID_EXs_RS2_OUT_reg_0_inst : DFFS_X1 port map( D => n2768, CK => Clk, 
                           SN => Rst, Q => n1965, QN => DataP_Rs2_0_port);
   DataP_ID_EXs_RS2_OUT_reg_3_inst : DFFS_X1 port map( D => n2767, CK => Clk, 
                           SN => Rst, Q => n_1331, QN => DataP_Rs2_3_port);
   DataP_MEM_WB_s_RD_OUT_reg_1_inst : DFFS_X1 port map( D => n1637, CK => Clk, 
                           SN => Rst, Q => n2228, QN => DataP_add_D_1_port);
   DataP_MEM_WB_s_RD_OUT_reg_3_inst : DFFS_X1 port map( D => n2777, CK => Clk, 
                           SN => Rst, Q => n2775, QN => DataP_add_D_3_port);
   DataP_EX_MEM_s_RD_OUT_reg_1_inst : DFFS_X1 port map( D => n11, CK => Clk, SN
                           => Rst, Q => n529, QN => DataP_dest_M_1_port);
   DataP_IF_IDs_IR_OUT_reg_30_inst : DFFS_X1 port map( D => IRAM_DATA_OUT(30), 
                           CK => Clk, SN => n36, Q => n2377, QN => n515);
   CU_I_aluOpcode1_reg_0_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_0_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_0_port, QN 
                           => n2395);
   CU_I_aluOpcode1_reg_1_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_1_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_1_port, QN 
                           => n2379);
   DataP_PC_reg_O_reg_30_inst : DFF_X2 port map( D => DataP_PC_reg_N32, CK => 
                           Clk, Q => DataP_pc_out_30_port, QN => n_1332);
   DataP_EX_MEM_s_ALU_OUT_reg_23_inst : DFFS_X2 port map( D => n2217, CK => Clk
                           , SN => Rst, Q => n2413, QN => 
                           DataP_alu_out_M_23_port);
   DataP_PC_reg_O_reg_26_inst : DFF_X2 port map( D => DataP_PC_reg_N28, CK => 
                           Clk, Q => DataP_pc_out_26_port, QN => n_1333);
   DataP_PC_reg_O_reg_21_inst : DFF_X2 port map( D => DataP_PC_reg_N23, CK => 
                           Clk, Q => DataP_pc_out_21_port, QN => n_1334);
   DataP_EX_MEM_s_OPCODE_OUT_reg_2_inst : DFFS_X1 port map( D => n521, CK => 
                           Clk, SN => Rst, Q => n2147, QN => 
                           DataP_opcode_M_2_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_1_inst : DFFS_X1 port map( D => n2249, CK => 
                           Clk, SN => Rst, Q => n2776, QN => 
                           DataP_opcode_W_1_port);
   DataP_MEM_WB_s_OPCODE_OUT_reg_2_inst : DFFS_X1 port map( D => n1643, CK => 
                           Clk, SN => Rst, Q => n2779, QN => 
                           DataP_opcode_W_2_port);
   DataP_ID_EXs_PR_OUT_reg : DFFR_X1 port map( D => DataP_pr_D, CK => Clk, RN 
                           => Rst, Q => DataP_pr_E, QN => n_1335);
   DataP_ID_EXs_IMM_OUT_reg_30_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_31_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_30_port, QN => n_1336);
   DataP_ID_EXs_IMM_OUT_reg_24_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_24_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_24_port, QN => n_1337);
   DataP_ID_EXs_IMM_OUT_reg_23_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_23_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_23_port, QN => n_1338);
   DataP_ID_EXs_IMM_OUT_reg_22_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_22_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_22_port, QN => n_1339);
   DataP_ID_EXs_IMM_OUT_reg_21_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_21_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_21_port, QN => n_1340);
   DataP_ID_EXs_IMM_OUT_reg_20_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_20_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_20_port, QN => n_1341);
   DataP_ID_EXs_IMM_OUT_reg_19_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_19_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_19_port, QN => n_1342);
   DataP_ID_EXs_IMM_OUT_reg_18_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_18_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_18_port, QN => n_1343);
   DataP_ID_EXs_IMM_OUT_reg_17_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_17_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_17_port, QN => n_1344);
   DataP_ID_EXs_IMM_OUT_reg_16_inst : DFFR_X1 port map( D => 
                           DataP_imm_out_16_port, CK => Clk, RN => Rst, Q => 
                           DataP_IMM_s_16_port, QN => n_1345);
   CU_I_aluOpcode1_reg_3_inst : DFFR_X1 port map( D => CU_I_aluOpcode_i_3_port,
                           CK => Clk, RN => Rst, Q => ALU_OPCODE_i_3_port, QN 
                           => n2672);
   DataP_MEM_WB_s_ALU_OUT_reg_31_inst : DFFS_X1 port map( D => n2414, CK => Clk
                           , SN => Rst, Q => n2517, QN => 
                           DataP_alu_out_W_31_port);
   DataP_MEM_WB_s_ALU_OUT_reg_15_inst : DFFS_X1 port map( D => n2433, CK => Clk
                           , SN => Rst, Q => n2516, QN => 
                           DataP_alu_out_W_15_port);
   DataP_MEM_WB_s_ALU_OUT_reg_28_inst : DFFS_X1 port map( D => n2426, CK => Clk
                           , SN => Rst, Q => n2508, QN => 
                           DataP_alu_out_W_28_port);
   DataP_MEM_WB_s_ALU_OUT_reg_24_inst : DFFS_X1 port map( D => n2427, CK => Clk
                           , SN => Rst, Q => n2513, QN => 
                           DataP_alu_out_W_24_port);
   DataP_MEM_WB_s_ALU_OUT_reg_22_inst : DFFS_X1 port map( D => n2428, CK => Clk
                           , SN => Rst, Q => n2512, QN => 
                           DataP_alu_out_W_22_port);
   DataP_MEM_WB_s_ALU_OUT_reg_18_inst : DFFS_X1 port map( D => n2425, CK => Clk
                           , SN => Rst, Q => n2505, QN => 
                           DataP_alu_out_W_18_port);
   DataP_MEM_WB_s_ALU_OUT_reg_12_inst : DFFS_X1 port map( D => n2424, CK => Clk
                           , SN => Rst, Q => n2492, QN => 
                           DataP_alu_out_W_12_port);
   DataP_MEM_WB_s_ALU_OUT_reg_25_inst : DFFS_X1 port map( D => n2422, CK => Clk
                           , SN => Rst, Q => n2507, QN => 
                           DataP_alu_out_W_25_port);
   DataP_MEM_WB_s_ALU_OUT_reg_20_inst : DFFS_X1 port map( D => n2420, CK => Clk
                           , SN => Rst, Q => n2506, QN => 
                           DataP_alu_out_W_20_port);
   DataP_MEM_WB_s_ALU_OUT_reg_19_inst : DFFS_X1 port map( D => n2421, CK => Clk
                           , SN => Rst, Q => n2498, QN => 
                           DataP_alu_out_W_19_port);
   DataP_MEM_WB_s_ALU_OUT_reg_13_inst : DFFS_X1 port map( D => n2423, CK => Clk
                           , SN => Rst, Q => n2504, QN => 
                           DataP_alu_out_W_13_port);
   DataP_MEM_WB_s_ALU_OUT_reg_30_inst : DFFS_X1 port map( D => n2417, CK => Clk
                           , SN => Rst, Q => n2496, QN => 
                           DataP_alu_out_W_30_port);
   DataP_MEM_WB_s_ALU_OUT_reg_26_inst : DFFS_X1 port map( D => n2415, CK => Clk
                           , SN => Rst, Q => n2500, QN => 
                           DataP_alu_out_W_26_port);
   DataP_MEM_WB_s_ALU_OUT_reg_21_inst : DFFS_X1 port map( D => n2419, CK => Clk
                           , SN => Rst, Q => n2499, QN => 
                           DataP_alu_out_W_21_port);
   DataP_MEM_WB_s_ALU_OUT_reg_17_inst : DFFS_X1 port map( D => n2416, CK => Clk
                           , SN => Rst, Q => n2493, QN => 
                           DataP_alu_out_W_17_port);
   DataP_MEM_WB_s_ALU_OUT_reg_14_inst : DFFS_X1 port map( D => n2418, CK => Clk
                           , SN => Rst, Q => n2497, QN => 
                           DataP_alu_out_W_14_port);
   DataP_MEM_WB_s_ALU_OUT_reg_16_inst : DFFS_X1 port map( D => n2412, CK => Clk
                           , SN => Rst, Q => n2511, QN => 
                           DataP_alu_out_W_16_port);
   DataP_MEM_WB_s_ALU_OUT_reg_6_inst : DFFS_X1 port map( D => n2410, CK => Clk,
                           SN => Rst, Q => n2515, QN => DataP_alu_out_W_6_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_2_inst : DFFS_X1 port map( D => n2471, CK => Clk,
                           SN => Rst, Q => n2514, QN => DataP_alu_out_W_2_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_1_inst : DFFS_X1 port map( D => n2469, CK => Clk,
                           SN => Rst, Q => n2522, QN => DataP_alu_out_W_1_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_7_inst : DFFS_X1 port map( D => n2468, CK => Clk,
                           SN => Rst, Q => n2510, QN => DataP_alu_out_W_7_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_3_inst : DFFS_X1 port map( D => n2478, CK => Clk,
                           SN => Rst, Q => n2523, QN => DataP_alu_out_W_3_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_10_inst : DFFS_X1 port map( D => n2409, CK => Clk
                           , SN => Rst, Q => n2503, QN => 
                           DataP_alu_out_W_10_port);
   DataP_MEM_WB_s_ALU_OUT_reg_8_inst : DFFS_X1 port map( D => n2408, CK => Clk,
                           SN => Rst, Q => n2502, QN => DataP_alu_out_W_8_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_4_inst : DFFS_X1 port map( D => n2466, CK => Clk,
                           SN => Rst, Q => n2509, QN => DataP_alu_out_W_4_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_11_inst : DFFS_X1 port map( D => n2431, CK => Clk
                           , SN => Rst, Q => n2518, QN => 
                           DataP_alu_out_W_11_port);
   DataP_MEM_WB_s_ALU_OUT_reg_9_inst : DFFS_X1 port map( D => n2477, CK => Clk,
                           SN => Rst, Q => n2519, QN => DataP_alu_out_W_9_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_5_inst : DFFS_X1 port map( D => n2450, CK => Clk,
                           SN => Rst, Q => n2520, QN => DataP_alu_out_W_5_port)
                           ;
   DataP_MEM_WB_s_ALU_OUT_reg_29_inst : DFFS_X1 port map( D => n2008, CK => Clk
                           , SN => Rst, Q => n2501, QN => 
                           DataP_alu_out_W_29_port);
   DataP_MEM_WB_s_ALU_OUT_reg_27_inst : DFFS_X1 port map( D => n2411, CK => Clk
                           , SN => Rst, Q => n2495, QN => 
                           DataP_alu_out_W_27_port);
   DataP_MEM_WB_s_ALU_OUT_reg_23_inst : DFFS_X1 port map( D => n2413, CK => Clk
                           , SN => Rst, Q => n2494, QN => 
                           DataP_alu_out_W_23_port);
   DataP_MEM_WB_s_ALU_OUT_reg_0_inst : DFFS_X1 port map( D => n2472, CK => Clk,
                           SN => Rst, Q => n2521, QN => DataP_alu_out_W_0_port)
                           ;
   CU_I_cw1_reg_10_inst : DFFS_X1 port map( D => n2007, CK => Clk, SN => Rst, Q
                           => n432, QN => n2475);
   CU_I_cw1_reg_9_inst : DFFS_X1 port map( D => n1961, CK => Clk, SN => Rst, Q 
                           => n399, QN => n2481);
   DataP_ID_EXs_A_OUT_reg_31_inst : DFFS_X1 port map( D => n2006, CK => Clk, SN
                           => Rst, Q => n2436, QN => DataP_A_s_31_port);
   DataP_ID_EXs_A_OUT_reg_6_inst : DFFS_X1 port map( D => n2005, CK => Clk, SN 
                           => Rst, Q => n2462, QN => DataP_A_s_6_port);
   DataP_ID_EXs_A_OUT_reg_5_inst : DFFS_X1 port map( D => n2004, CK => Clk, SN 
                           => Rst, Q => n2443, QN => DataP_A_s_5_port);
   DataP_ID_EXs_A_OUT_reg_4_inst : DFFS_X1 port map( D => n2003, CK => Clk, SN 
                           => Rst, Q => n2470, QN => DataP_A_s_4_port);
   DataP_ID_EXs_A_OUT_reg_3_inst : DFFS_X1 port map( D => n2002, CK => Clk, SN 
                           => Rst, Q => n2458, QN => DataP_A_s_3_port);
   DataP_ID_EXs_A_OUT_reg_30_inst : DFFS_X1 port map( D => n2001, CK => Clk, SN
                           => Rst, Q => n2437, QN => DataP_A_s_30_port);
   CU_I_aluOpcode1_reg_4_inst : DFFS_X1 port map( D => n2000, CK => Clk, SN => 
                           Rst, Q => n443, QN => n2491);
   DataP_ID_EXs_A_OUT_reg_0_inst : DFFS_X1 port map( D => n1999, CK => Clk, SN 
                           => Rst, Q => n2460, QN => DataP_A_s_0_port);
   DataP_ID_EXs_A_OUT_reg_25_inst : DFFS_X1 port map( D => n1998, CK => Clk, SN
                           => Rst, Q => n2453, QN => DataP_A_s_25_port);
   DataP_ID_EXs_A_OUT_reg_24_inst : DFFS_X1 port map( D => n1997, CK => Clk, SN
                           => Rst, Q => n2463, QN => DataP_A_s_24_port);
   DataP_ID_EXs_A_OUT_reg_23_inst : DFFS_X1 port map( D => n1996, CK => Clk, SN
                           => Rst, Q => n2439, QN => DataP_A_s_23_port);
   DataP_ID_EXs_A_OUT_reg_22_inst : DFFS_X1 port map( D => n1995, CK => Clk, SN
                           => Rst, Q => n2464, QN => DataP_A_s_22_port);
   DataP_ID_EXs_A_OUT_reg_21_inst : DFFS_X1 port map( D => n1994, CK => Clk, SN
                           => Rst, Q => n2446, QN => DataP_A_s_21_port);
   DataP_ID_EXs_A_OUT_reg_20_inst : DFFS_X1 port map( D => n1993, CK => Clk, SN
                           => Rst, Q => n2454, QN => DataP_A_s_20_port);
   DataP_ID_EXs_A_OUT_reg_19_inst : DFFS_X1 port map( D => n1992, CK => Clk, SN
                           => Rst, Q => n2447, QN => DataP_A_s_19_port);
   DataP_ID_EXs_A_OUT_reg_18_inst : DFFS_X1 port map( D => n1991, CK => Clk, SN
                           => Rst, Q => n2455, QN => DataP_A_s_18_port);
   DataP_ID_EXs_A_OUT_reg_17_inst : DFFS_X1 port map( D => n1990, CK => Clk, SN
                           => Rst, Q => n2440, QN => DataP_A_s_17_port);
   DataP_ID_EXs_A_OUT_reg_16_inst : DFFS_X1 port map( D => n1989, CK => Clk, SN
                           => Rst, Q => n2465, QN => DataP_A_s_16_port);
   DataP_ID_EXs_A_OUT_reg_15_inst : DFFS_X1 port map( D => n1988, CK => Clk, SN
                           => Rst, Q => n2441, QN => DataP_A_s_15_port);
   DataP_ID_EXs_A_OUT_reg_14_inst : DFFS_X1 port map( D => n1987, CK => Clk, SN
                           => Rst, Q => n2448, QN => DataP_A_s_14_port);
   DataP_ID_EXs_A_OUT_reg_13_inst : DFFS_X1 port map( D => n1986, CK => Clk, SN
                           => Rst, Q => n2456, QN => DataP_A_s_13_port);
   DataP_ID_EXs_A_OUT_reg_12_inst : DFFS_X1 port map( D => n1985, CK => Clk, SN
                           => Rst, Q => n2442, QN => DataP_A_s_12_port);
   DataP_ID_EXs_A_OUT_reg_11_inst : DFFS_X1 port map( D => n1984, CK => Clk, SN
                           => Rst, Q => n2449, QN => DataP_A_s_11_port);
   DataP_ID_EXs_A_OUT_reg_10_inst : DFFS_X1 port map( D => n1983, CK => Clk, SN
                           => Rst, Q => n2457, QN => DataP_A_s_10_port);
   DataP_ID_EXs_A_OUT_reg_7_inst : DFFS_X1 port map( D => n1982, CK => Clk, SN 
                           => Rst, Q => n2451, QN => DataP_A_s_7_port);
   DataP_ID_EXs_A_OUT_reg_1_inst : DFFS_X1 port map( D => n1981, CK => Clk, SN 
                           => Rst, Q => n2461, QN => DataP_A_s_1_port);
   DataP_ID_EXs_A_OUT_reg_28_inst : DFFS_X1 port map( D => n1980, CK => Clk, SN
                           => Rst, Q => n2452, QN => DataP_A_s_28_port);
   DataP_ID_EXs_A_OUT_reg_26_inst : DFFS_X1 port map( D => n1979, CK => Clk, SN
                           => Rst, Q => n2445, QN => DataP_A_s_26_port);
   DataP_ID_EXs_A_OUT_reg_29_inst : DFFS_X1 port map( D => n1978, CK => Clk, SN
                           => Rst, Q => n2444, QN => DataP_A_s_29_port);
   DataP_ID_EXs_A_OUT_reg_27_inst : DFFS_X1 port map( D => n1977, CK => Clk, SN
                           => Rst, Q => n2438, QN => DataP_A_s_27_port);
   DataP_PC_reg_O_reg_11_inst : DFFRS_X1 port map( D => DataP_PC_reg_N13, CK =>
                           Clk, RN => n1976, SN => n1976, Q => 
                           DataP_pc_out_11_port, QN => n_1346);
   DataP_ID_EXs_NPC_L_OUT_reg_31_inst : DFFR_X1 port map( D => 
                           DataP_link_addr_D_31_port, CK => Clk, RN => Rst, Q 
                           => n_1347, QN => n292);
   DataP_PC_reg_O_reg_20_inst : DFFRS_X1 port map( D => DataP_PC_reg_N22, CK =>
                           Clk, RN => n1975, SN => n1975, Q => 
                           DataP_pc_out_20_port, QN => n_1348);
   DataP_ID_EXs_RS2_OUT_reg_1_inst : DFFS_X1 port map( D => n2770, CK => Clk, 
                           SN => Rst, Q => n_1349, QN => DataP_Rs2_1_port);
   DataP_EX_MEM_s_ALU_OUT_reg_29_inst : DFFS_X1 port map( D => n299, CK => Clk,
                           SN => Rst, Q => n2008, QN => DataP_alu_out_M_29_port
                           );
   DataP_ID_EXs_RS2_OUT_reg_4_inst : DFFS_X1 port map( D => n2769, CK => Clk, 
                           SN => Rst, Q => n2029, QN => DataP_Rs2_4_port);
   DataP_ID_EXs_RS2_OUT_reg_2_inst : DFFS_X1 port map( D => n1974, CK => Clk, 
                           SN => Rst, Q => n1603, QN => DataP_Rs2_2_port);
   DataP_MEM_WB_s_RD_OUT_reg_4_inst : DFFR_X1 port map( D => n1720, CK => Clk, 
                           RN => Rst, Q => DataP_add_D_4_port, QN => n540);
   DataP_ID_EXs_OPCODE_OUT_reg_5_inst : DFFR_X1 port map( D => IR_CU_31, CK => 
                           Clk, RN => Rst, Q => n_1350, QN => n17);
   DataP_IF_IDs_IR_OUT_reg_27_inst : DFFR_X1 port map( D => IRAM_DATA_OUT(27), 
                           CK => Clk, RN => n36, Q => IR_CU_27, QN => n504);
   DataP_EX_MEM_s_ALU_OUT_reg_0_inst : DFFS_X1 port map( D => n2243, CK => Clk,
                           SN => Rst, Q => n2472, QN => DRAM_ADDRESS_0_port);
   DataP_PC_reg_O_reg_28_inst : DFF_X1 port map( D => DataP_PC_reg_N30, CK => 
                           Clk, Q => DataP_pc_out_28_port, QN => n_1351);
   DataP_EX_MEM_s_ALU_OUT_reg_27_inst : DFFS_X1 port map( D => n301, CK => Clk,
                           SN => Rst, Q => n2411, QN => DataP_alu_out_M_27_port
                           );
   DataP_PC_reg_O_reg_15_inst : DFF_X1 port map( D => DataP_PC_reg_N17, CK => 
                           Clk, Q => DataP_pc_out_15_port, QN => n_1352);
   DataP_EX_MEM_s_ALU_OUT_reg_22_inst : DFFS_X2 port map( D => n1708, CK => Clk
                           , SN => Rst, Q => n2428, QN => 
                           DataP_alu_out_M_22_port);
   DataP_ID_EXs_OPCODE_OUT_reg_2_inst : DFFR_X1 port map( D => IR_CU_28, CK => 
                           Clk, RN => Rst, Q => n_1353, QN => n521);
   DataP_PC_reg_O_reg_25_inst : DFF_X2 port map( D => DataP_PC_reg_N27, CK => 
                           Clk, Q => DataP_pc_out_25_port, QN => n_1354);
   DataP_PC_reg_O_reg_24_inst : DFF_X1 port map( D => DataP_PC_reg_N26, CK => 
                           Clk, Q => DataP_pc_out_24_port, QN => n_1355);
   DataP_PC_reg_O_reg_17_inst : DFF_X1 port map( D => DataP_PC_reg_N19, CK => 
                           Clk, Q => DataP_pc_out_17_port, QN => n_1356);
   DataP_EX_MEM_s_ALU_OUT_reg_26_inst : DFFS_X2 port map( D => n1598, CK => Clk
                           , SN => Rst, Q => n2415, QN => 
                           DataP_alu_out_M_26_port);
   DataP_EX_MEM_s_ALU_OUT_reg_17_inst : DFFS_X2 port map( D => n1611, CK => Clk
                           , SN => Rst, Q => n2416, QN => 
                           DataP_alu_out_M_17_port);
   DataP_PC_reg_O_reg_0_inst : DFF_X1 port map( D => DataP_PC_reg_N2, CK => Clk
                           , Q => DataP_pc_out_0, QN => n_1357);
   DataP_EX_MEM_s_ALU_OUT_reg_7_inst : DFFS_X2 port map( D => n1569, CK => Clk,
                           SN => Rst, Q => n2468, QN => DRAM_ADDRESS_7_port);
   DataP_PC_reg_O_reg_29_inst : DFF_X1 port map( D => DataP_PC_reg_N31, CK => 
                           Clk, Q => DataP_pc_out_29_port, QN => n_1358);
   U1484 : NOR2_X1 port map( A1 => n3294, A2 => n3234, ZN => n3909);
   U1485 : INV_X2 port map( A => n3880, ZN => n2129);
   U1486 : NAND2_X1 port map( A1 => n3689, A2 => DataP_alu_a_in_23_port, ZN => 
                           n1548);
   U1487 : NOR2_X1 port map( A1 => DataP_alu_b_in_8_port, A2 => n1577, ZN => 
                           n1549);
   U1488 : NAND4_X1 port map( A1 => n3527, A2 => n3526, A3 => n3525, A4 => 
                           n3524, ZN => n1550);
   U1489 : OAI211_X1 port map( C1 => n3662, C2 => n3682, A => n1566, B => n2169
                           , ZN => n1551);
   U1490 : AND2_X2 port map( A1 => n2527, A2 => n1570, ZN => n3662);
   U1491 : NAND2_X1 port map( A1 => n2667, A2 => n2665, ZN => n1552);
   U1492 : NAND2_X1 port map( A1 => n2532, A2 => n3730, ZN => n2531);
   U1493 : NAND2_X1 port map( A1 => n1553, A2 => n1554, ZN => 
                           DataP_alu_a_in_0_port);
   U1494 : INV_X1 port map( A => n3331, ZN => n1553);
   U1495 : INV_X1 port map( A => n3332, ZN => n1554);
   U1496 : AND2_X1 port map( A1 => n3661, A2 => n3660, ZN => n2219);
   U1497 : AOI21_X1 port map( B1 => DataP_alu_a_in_4_port, B2 => n2380, A => 
                           n1922, ZN => n2256);
   U1498 : NAND2_X1 port map( A1 => n2727, A2 => n3797, ZN => n2718);
   U1499 : NAND3_X1 port map( A1 => n1552, A2 => n2718, A3 => n2713, ZN => 
                           n1555);
   U1500 : AND2_X2 port map( A1 => n2727, A2 => n3797, ZN => n2382);
   U1501 : NAND2_X1 port map( A1 => n2745, A2 => n2071, ZN => n1556);
   U1502 : NOR2_X1 port map( A1 => n2746, A2 => n3826, ZN => n1557);
   U1503 : XNOR2_X1 port map( A => n1556, B => n1557, ZN => n1558);
   U1504 : AOI21_X1 port map( B1 => n1558, B2 => n2129, A => n3833, ZN => n299)
                           ;
   U1505 : NAND2_X1 port map( A1 => n1558, A2 => n1607, ZN => n1659);
   U1506 : NOR2_X1 port map( A1 => n1559, A2 => n1838, ZN => n3423);
   U1507 : NAND4_X1 port map( A1 => n2658, A2 => n1587, A3 => n2660, A4 => 
                           n1595, ZN => n1559);
   U1508 : NOR2_X1 port map( A1 => sra_131_SH_4_port, A2 => n1559, ZN => n1704)
                           ;
   U1509 : AND4_X1 port map( A1 => n1560, A2 => n1561, A3 => n1562, A4 => n1563
                           , ZN => n4103);
   U1510 : AND3_X1 port map( A1 => n3707, A2 => n3898, A3 => n3875, ZN => n1560
                           );
   U1511 : AND4_X1 port map( A1 => n3741, A2 => n3731, A3 => n3872, A4 => n3613
                           , ZN => n1561);
   U1512 : AND4_X1 port map( A1 => n3859, A2 => n3853, A3 => n3603, A4 => n3536
                           , ZN => n1562);
   U1513 : AND3_X1 port map( A1 => n3542, A2 => n3541, A3 => n3848, ZN => n1563
                           );
   U1514 : OAI211_X1 port map( C1 => n2728, C2 => n2382, A => n1555, B => n2712
                           , ZN => n1564);
   U1515 : NAND3_X1 port map( A1 => n2192, A2 => n3690, A3 => n2193, ZN => 
                           n1565);
   U1516 : BUF_X2 port map( A => n2233, Z => n2226);
   U1517 : CLKBUF_X3 port map( A => n3401, Z => n3213);
   U1518 : AOI211_X4 port map( C1 => n2299, C2 => n2289, A => n2287, B => n2288
                           , ZN => n2290);
   U1519 : MUX2_X2 port map( A => n3413, B => n3200, S => n3886, Z => n3414);
   U1520 : AND2_X1 port map( A1 => n3685, A2 => n3649, ZN => n1566);
   U1521 : AND2_X1 port map( A1 => n3685, A2 => n3649, ZN => n3684);
   U1522 : NAND2_X1 port map( A1 => n2077, A2 => n1593, ZN => n1567);
   U1523 : INV_X2 port map( A => n2072, ZN => n3207);
   U1524 : NOR2_X1 port map( A1 => n2659, A2 => n2090, ZN => n1568);
   U1525 : AOI211_X1 port map( C1 => n3228, C2 => n1909, A => n1914, B => n1918
                           , ZN => n1569);
   U1526 : AOI211_X1 port map( C1 => n3228, C2 => n1909, A => n1914, B => n1918
                           , ZN => n350);
   U1527 : NAND2_X1 port map( A1 => n2173, A2 => n2528, ZN => n1570);
   U1528 : AND3_X1 port map( A1 => n1636, A2 => n3681, A3 => n3686, ZN => n1571
                           );
   U1529 : AND3_X1 port map( A1 => n1636, A2 => n3681, A3 => n3686, ZN => n3712
                           );
   U1530 : BUF_X1 port map( A => n3221, Z => n1572);
   U1531 : AND4_X1 port map( A1 => n3478, A2 => n3477, A3 => n3475, A4 => n3476
                           , ZN => n1573);
   U1532 : AND2_X2 port map( A1 => n2723, A2 => n1599, ZN => n1574);
   U1533 : AND2_X1 port map( A1 => n2723, A2 => n1599, ZN => n3709);
   U1534 : BUF_X2 port map( A => DataP_alu_b_in_11_port, Z => n2151);
   U1535 : BUF_X1 port map( A => DataP_alu_b_in_8_port, Z => n1575);
   U1536 : INV_X2 port map( A => n1753, ZN => DataP_alu_b_in_17_port);
   U1537 : BUF_X1 port map( A => n2188, Z => n1576);
   U1538 : BUF_X1 port map( A => DataP_alu_b_in_9_port, Z => n1577);
   U1539 : OAI211_X1 port map( C1 => n2772, C2 => n2478, A => n2661, B => n2662
                           , ZN => n1578);
   U1540 : BUF_X2 port map( A => DataP_alu_b_in_10_port, Z => n2165);
   U1541 : AND2_X1 port map( A1 => n2657, A2 => n2656, ZN => n1579);
   U1542 : AND4_X1 port map( A1 => n3317, A2 => n3318, A3 => n3316, A4 => n3315
                           , ZN => n2380);
   U1543 : NAND2_X1 port map( A1 => n1709, A2 => n1580, ZN => n3694);
   U1544 : NOR2_X1 port map( A1 => n3641, A2 => n3640, ZN => n1580);
   U1545 : NAND2_X1 port map( A1 => n2076, A2 => n1580, ZN => n1760);
   U1546 : OAI211_X2 port map( C1 => n2427, C2 => n2771, A => n1841, B => n1842
                           , ZN => DataP_alu_b_in_24_port);
   U1547 : BUF_X2 port map( A => n3548, Z => n1581);
   U1548 : AND2_X1 port map( A1 => DataP_alu_b_in_18_port, A2 => n1694, ZN => 
                           n2731);
   U1549 : INV_X2 port map( A => n3201, ZN => n3048);
   U1550 : AOI21_X1 port map( B1 => n3635, B2 => n3636, A => n2715, ZN => n1582
                           );
   U1551 : NAND2_X1 port map( A1 => n2246, A2 => DataP_IMM_s_1_port, ZN => 
                           n1583);
   U1552 : NAND2_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n2535, ZN => 
                           n2534);
   U1553 : NAND2_X1 port map( A1 => n1644, A2 => n1662, ZN => n1584);
   U1554 : AND2_X1 port map( A1 => n3449, A2 => DataP_alu_a_in_10_port, ZN => 
                           n3489);
   U1555 : NAND4_X1 port map( A1 => n1568, A2 => n1587, A3 => n1595, A4 => 
                           n1586, ZN => n1585);
   U1556 : INV_X1 port map( A => n1578, ZN => n1586);
   U1557 : AND2_X1 port map( A1 => n2656, A2 => n2657, ZN => n1587);
   U1558 : NAND2_X1 port map( A1 => n3666, A2 => DataP_alu_a_in_20_port, ZN => 
                           n1588);
   U1559 : AND2_X1 port map( A1 => n2154, A2 => n2153, ZN => n1589);
   U1560 : OAI211_X1 port map( C1 => n2604, C2 => n2607, A => n2603, B => n3686
                           , ZN => n1590);
   U1561 : OR2_X1 port map( A1 => n3295, A2 => n1718, ZN => n1673);
   U1562 : INV_X1 port map( A => n3429, ZN => n1591);
   U1563 : OAI211_X1 port map( C1 => n2728, C2 => n2382, A => n2711, B => n2712
                           , ZN => n1592);
   U1564 : AND2_X1 port map( A1 => n3308, A2 => n3309, ZN => n1593);
   U1565 : OAI21_X1 port map( B1 => n2596, B2 => n2535, A => n2701, ZN => n1594
                           );
   U1566 : AND4_X1 port map( A1 => n3314, A2 => n3313, A3 => n3312, A4 => n3311
                           , ZN => n1595);
   U1567 : AND4_X1 port map( A1 => n3314, A2 => n3313, A3 => n3312, A4 => n3311
                           , ZN => n2240);
   U1568 : CLKBUF_X3 port map( A => n2773, Z => n1627);
   U1569 : AND2_X1 port map( A1 => n3683, A2 => n1663, ZN => n1596);
   U1570 : NAND2_X1 port map( A1 => n1683, A2 => n3721, ZN => n2583);
   U1571 : XNOR2_X1 port map( A => DataP_Rs2_3_port, B => DataP_add_D_3_port, 
                           ZN => n1962);
   U1572 : XOR2_X1 port map( A => lt_x_135_B_12_port, B => n1941, Z => n1597);
   U1573 : NOR2_X2 port map( A1 => n2068, A2 => n3480, ZN => n1941);
   U1574 : BUF_X1 port map( A => n303, Z => n1598);
   U1575 : NOR2_X1 port map( A1 => n3659, A2 => n1737, ZN => n1599);
   U1576 : BUF_X1 port map( A => DataP_alu_b_in_19_port, Z => n1600);
   U1577 : CLKBUF_X3 port map( A => n3401, Z => n3214);
   U1578 : BUF_X1 port map( A => n2250, Z => n1601);
   U1579 : INV_X1 port map( A => n2074, ZN => lt_x_135_B_5_port);
   U1580 : INV_X2 port map( A => n3886, ZN => n2108);
   U1581 : OR2_X1 port map( A1 => n1732, A2 => n2322, ZN => n1602);
   U1582 : INV_X1 port map( A => n3886, ZN => n1694);
   U1583 : AND2_X1 port map( A1 => DataP_alu_a_in_24_port, A2 => n1691, ZN => 
                           n1604);
   U1584 : AND2_X1 port map( A1 => n1904, A2 => n3717, ZN => n1605);
   U1585 : AND2_X1 port map( A1 => n2129, A2 => n1656, ZN => n1607);
   U1586 : NAND2_X1 port map( A1 => n3540, A2 => n1696, ZN => n1608);
   U1587 : NAND2_X1 port map( A1 => n1904, A2 => n2727, ZN => n1609);
   U1588 : XOR2_X1 port map( A => n1830, B => n2030, Z => n1610);
   U1589 : BUF_X1 port map( A => n323, Z => n1611);
   U1590 : XNOR2_X1 port map( A => n1612, B => n2404, ZN => n3796);
   U1591 : NAND2_X1 port map( A1 => n1626, A2 => n1548, ZN => n1612);
   U1592 : NAND2_X1 port map( A1 => n2697, A2 => n2696, ZN => n1613);
   U1593 : NAND2_X1 port map( A1 => n2697, A2 => n2696, ZN => n3777);
   U1594 : BUF_X1 port map( A => n1581, Z => n1614);
   U1595 : OAI21_X1 port map( B1 => n2681, B2 => n2128, A => n2680, ZN => n1615
                           );
   U1596 : OR2_X4 port map( A1 => n3343, A2 => n3342, ZN => 
                           DataP_alu_a_in_6_port);
   U1597 : NAND2_X1 port map( A1 => n1615, A2 => DataP_alu_a_in_6_port, ZN => 
                           n1616);
   U1598 : NAND2_X1 port map( A1 => n3609, A2 => n1616, ZN => n3855);
   U1599 : INV_X1 port map( A => DataP_alu_a_in_6_port, ZN => n3857);
   U1600 : AND2_X1 port map( A1 => n3884, A2 => n2489, ZN => n1617);
   U1601 : AND2_X1 port map( A1 => n3884, A2 => n2489, ZN => n1618);
   U1602 : AND2_X1 port map( A1 => n1571, A2 => n1582, ZN => n1619);
   U1603 : BUF_X1 port map( A => n3221, Z => n1620);
   U1604 : NAND2_X1 port map( A1 => n1679, A2 => n3718, ZN => n3799);
   U1605 : BUF_X1 port map( A => DataP_dest_M_3_port, Z => n1621);
   U1606 : BUF_X1 port map( A => n3575, Z => n1622);
   U1607 : BUF_X1 port map( A => n1581, Z => n1623);
   U1608 : BUF_X1 port map( A => n304, Z => n1624);
   U1609 : BUF_X1 port map( A => DataP_dest_M_4_port, Z => n1625);
   U1610 : NAND3_X1 port map( A1 => n2192, A2 => n3690, A3 => n2133, ZN => 
                           n1626);
   U1611 : BUF_X2 port map( A => n2781, Z => n2773);
   U1612 : BUF_X1 port map( A => n540, Z => n1628);
   U1613 : INV_X1 port map( A => n1628, ZN => n1629);
   U1614 : BUF_X1 port map( A => n536, Z => n1630);
   U1615 : BUF_X1 port map( A => n3221, Z => n1631);
   U1616 : BUF_X1 port map( A => n3796, Z => n1632);
   U1617 : NAND2_X1 port map( A1 => n1590, A2 => n2608, ZN => n1633);
   U1618 : NOR2_X1 port map( A1 => n3861, A2 => n3868, ZN => n1634);
   U1619 : BUF_X1 port map( A => n2241, Z => n1635);
   U1620 : BUF_X1 port map( A => n1551, Z => n1636);
   U1621 : INV_X1 port map( A => DataP_dest_M_1_port, ZN => n1637);
   U1622 : OR2_X1 port map( A1 => n2190, A2 => DataP_alu_a_in_26_port, ZN => 
                           n3719);
   U1623 : INV_X1 port map( A => DataP_dest_M_2_port, ZN => n1638);
   U1624 : NAND2_X1 port map( A1 => DataP_Rs2_4_port, A2 => DataP_add_D_4_port,
                           ZN => n1641);
   U1625 : NAND2_X1 port map( A1 => n1639, A2 => n1640, ZN => n1642);
   U1626 : NAND2_X1 port map( A1 => n1641, A2 => n1642, ZN => n3245);
   U1627 : INV_X1 port map( A => DataP_Rs2_4_port, ZN => n1639);
   U1628 : INV_X1 port map( A => DataP_add_D_4_port, ZN => n1640);
   U1629 : INV_X1 port map( A => DataP_opcode_M_2_port, ZN => n1643);
   U1630 : BUF_X1 port map( A => n3845, Z => n1644);
   U1631 : BUF_X1 port map( A => n3221, Z => n1645);
   U1632 : BUF_X1 port map( A => n1571, Z => n1646);
   U1633 : BUF_X1 port map( A => n3642, Z => n1647);
   U1634 : BUF_X1 port map( A => n3609, Z => n1648);
   U1635 : AND2_X1 port map( A1 => n538, A2 => n540, ZN => n1649);
   U1636 : NAND4_X1 port map( A1 => n1757, A2 => n1649, A3 => n2228, A4 => 
                           n1630, ZN => n1650);
   U1637 : AND2_X1 port map( A1 => n3289, A2 => n1650, ZN => n1651);
   U1638 : NAND3_X1 port map( A1 => n1742, A2 => n3290, A3 => n1651, ZN => 
                           n3293);
   U1639 : NAND2_X1 port map( A1 => n3245, A2 => n1650, ZN => n2637);
   U1640 : INV_X1 port map( A => n1650, ZN => n1671);
   U1641 : INV_X1 port map( A => n2228, ZN => n2229);
   U1642 : XNOR2_X1 port map( A => n2249, B => n2147, ZN => n1652);
   U1643 : NOR2_X1 port map( A1 => n1652, A2 => n18, ZN => n1653);
   U1644 : AND2_X1 port map( A1 => n2195, A2 => n2387, ZN => n1654);
   U1645 : OAI21_X1 port map( B1 => n1653, B2 => n1654, A => 
                           DataP_opcode_M_3_port, ZN => n3250);
   U1646 : NAND2_X1 port map( A1 => n2040, A2 => n1968, ZN => n1655);
   U1647 : NAND2_X1 port map( A1 => n1659, A2 => n1658, ZN => DataP_PC_reg_N31)
                           ;
   U1648 : INV_X2 port map( A => n4111, ZN => n1656);
   U1649 : NOR2_X2 port map( A1 => n4110, A2 => n4193, ZN => n1657);
   U1650 : AOI21_X2 port map( B1 => n3833, B2 => n2131, A => n1657, ZN => n1658
                           );
   U1651 : NAND2_X1 port map( A1 => n1661, A2 => n1660, ZN => n3629);
   U1652 : AND2_X1 port map( A1 => n2109, A2 => n2740, ZN => n1660);
   U1653 : NAND2_X1 port map( A1 => n3619, A2 => n2108, ZN => n1661);
   U1654 : BUF_X1 port map( A => n3548, Z => n3222);
   U1655 : AND3_X1 port map( A1 => n2194, A2 => n2094, A3 => n1579, ZN => n1755
                           );
   U1656 : BUF_X1 port map( A => n3844, Z => n1662);
   U1657 : NAND2_X4 port map( A1 => n3908, A2 => Rst, ZN => n4111);
   U1658 : BUF_X1 port map( A => n2239, Z => n1663);
   U1659 : OAI21_X1 port map( B1 => n313, B2 => n4111, A => n1664, ZN => 
                           DataP_PC_reg_N23);
   U1660 : OR2_X1 port map( A1 => n4110, A2 => n4201, ZN => n1664);
   U1661 : OAI22_X1 port map( A1 => n2678, A2 => n2677, B1 => 
                           DataP_alu_a_in_21_port, B2 => n2679, ZN => n2653);
   U1662 : NAND2_X1 port map( A1 => n2599, A2 => n2630, ZN => n2678);
   U1663 : NAND2_X1 port map( A1 => n2745, A2 => n2071, ZN => n2083);
   U1664 : NAND2_X1 port map( A1 => n1592, A2 => n2717, ZN => n2745);
   U1665 : OAI211_X1 port map( C1 => n3214, C2 => n37, A => n1666, B => n1665, 
                           ZN => n3332);
   U1666 : NAND2_X1 port map( A1 => n3209, A2 => DataP_alu_out_W_0_port, ZN => 
                           n1665);
   U1667 : NAND2_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_0_port, ZN => 
                           n1666);
   U1668 : XNOR2_X1 port map( A => n3423, B => n1748, ZN => n2681);
   U1669 : NAND2_X1 port map( A1 => n1668, A2 => n1667, ZN => n2430);
   U1670 : NOR2_X1 port map( A1 => n3885, A2 => n2385, ZN => n1667);
   U1671 : INV_X1 port map( A => n3722, ZN => n1668);
   U1672 : XNOR2_X1 port map( A => n1603, B => n538, ZN => n2143);
   U1673 : NAND3_X1 port map( A1 => n3294, A2 => n3290, A3 => n1669, ZN => 
                           n3279);
   U1674 : OR2_X1 port map( A1 => n3279, A2 => n1743, ZN => n2634);
   U1675 : NAND4_X1 port map( A1 => n3292, A2 => n1673, A3 => n1672, A4 => 
                           n2634, ZN => n3401);
   U1676 : NOR2_X2 port map( A1 => n1671, A2 => n1670, ZN => n1669);
   U1677 : INV_X2 port map( A => Rst, ZN => n1670);
   U1678 : AOI21_X1 port map( B1 => n3909, B2 => n2619, A => n432, ZN => n1672)
                           ;
   U1679 : NAND2_X1 port map( A1 => n2663, A2 => n2564, ZN => n2590);
   U1680 : XNOR2_X1 port map( A => n1675, B => n1674, ZN => n2663);
   U1681 : INV_X1 port map( A => n1576, ZN => n1674);
   U1682 : AOI21_X1 port map( B1 => n1565, B2 => n1677, A => n1676, ZN => n1675
                           );
   U1683 : INV_X1 port map( A => n3719, ZN => n1676);
   U1684 : AND2_X1 port map( A1 => n2705, A2 => n2584, ZN => n1677);
   U1685 : NAND2_X1 port map( A1 => n2664, A2 => n2720, ZN => n2595);
   U1686 : AND2_X2 port map( A1 => n1609, A2 => n1678, ZN => n2664);
   U1687 : NAND3_X1 port map( A1 => n1605, A2 => n1744, A3 => n2729, ZN => 
                           n1678);
   U1688 : NAND3_X1 port map( A1 => n2729, A2 => n1744, A3 => n3717, ZN => 
                           n1679);
   U1689 : NAND2_X1 port map( A1 => n2188, A2 => n1680, ZN => n1683);
   U1690 : OR2_X1 port map( A1 => n2096, A2 => n3719, ZN => n1680);
   U1691 : AOI21_X1 port map( B1 => n1681, B2 => n2582, A => n2746, ZN => n1682
                           );
   U1692 : NAND2_X1 port map( A1 => n1683, A2 => n3721, ZN => n1681);
   U1693 : NAND2_X1 port map( A1 => n2748, A2 => n1682, ZN => n2021);
   U1694 : NAND2_X2 port map( A1 => n2583, A2 => n2582, ZN => n2766);
   U1695 : NAND2_X2 port map( A1 => n1686, A2 => n2535, ZN => n2585);
   U1696 : NAND2_X2 port map( A1 => DataP_alu_a_in_25_port, A2 => n1684, ZN => 
                           n1821);
   U1697 : NOR2_X2 port map( A1 => n2588, A2 => n3851, ZN => n1684);
   U1698 : OAI21_X2 port map( B1 => DataP_alu_a_in_25_port, B2 => n1686, A => 
                           n3894, ZN => n1820);
   U1699 : XNOR2_X2 port map( A => DataP_alu_a_in_25_port, B => n1686, ZN => 
                           n3800);
   U1700 : NOR2_X2 port map( A1 => n2137, A2 => n1686, ZN => n2282);
   U1701 : AOI21_X2 port map( B1 => n2283, B2 => DataP_alu_b_in_24_port, A => 
                           n1685, ZN => n2356);
   U1702 : AND2_X2 port map( A1 => n2137, A2 => n1686, ZN => n1685);
   U1703 : INV_X2 port map( A => n2588, ZN => n1686);
   U1704 : NOR2_X2 port map( A1 => n1688, A2 => n1687, ZN => n2588);
   U1705 : NAND2_X2 port map( A1 => n3504, A2 => n3505, ZN => n1687);
   U1706 : NAND2_X2 port map( A1 => n3506, A2 => n3523, ZN => n1688);
   U1707 : OAI21_X1 port map( B1 => n3695, B2 => n1692, A => n1604, ZN => n3718
                           );
   U1708 : AOI21_X2 port map( B1 => n3695, B2 => n1694, A => n1689, ZN => n3788
                           );
   U1709 : NAND2_X2 port map( A1 => n1690, A2 => n1693, ZN => n1689);
   U1710 : INV_X2 port map( A => DataP_alu_a_in_24_port, ZN => n1690);
   U1711 : NAND2_X2 port map( A1 => n1693, A2 => n1698, ZN => n1691);
   U1712 : INV_X2 port map( A => n1693, ZN => n1692);
   U1713 : NAND2_X2 port map( A1 => DataP_alu_b_in_24_port, A2 => n3886, ZN => 
                           n1693);
   U1714 : OAI211_X1 port map( C1 => n3462, C2 => n1696, A => n1695, B => n1608
                           , ZN => n3464);
   U1715 : OR2_X2 port map( A1 => n3467, A2 => n1696, ZN => n1695);
   U1716 : AND2_X2 port map( A1 => n3464, A2 => n3491, ZN => n3488);
   U1717 : NAND2_X1 port map( A1 => n3488, A2 => n3489, ZN => n2612);
   U1718 : INV_X2 port map( A => n2108, ZN => n1696);
   U1719 : OAI21_X1 port map( B1 => n3448, B2 => n1698, A => n1697, ZN => n3449
                           );
   U1720 : NAND2_X1 port map( A1 => n2165, A2 => n1698, ZN => n1697);
   U1721 : INV_X1 port map( A => n2108, ZN => n1698);
   U1722 : XNOR2_X1 port map( A => n3460, B => n3459, ZN => n3448);
   U1723 : AND2_X1 port map( A1 => n2076, A2 => n1549, ZN => n3460);
   U1724 : OAI21_X1 port map( B1 => n2083, B2 => n1699, A => n2552, ZN => n2551
                           );
   U1725 : NAND2_X1 port map( A1 => n1701, A2 => n1700, ZN => n1699);
   U1726 : INV_X1 port map( A => n4111, ZN => n1700);
   U1727 : INV_X1 port map( A => n2752, ZN => n1701);
   U1728 : NAND2_X1 port map( A1 => n1703, A2 => n1702, ZN => n2752);
   U1729 : INV_X1 port map( A => n2704, ZN => n1702);
   U1730 : NAND2_X1 port map( A1 => n1617, A2 => n3826, ZN => n1703);
   U1731 : OAI21_X1 port map( B1 => n2044, B2 => n2128, A => n2163, ZN => n3421
                           );
   U1732 : XNOR2_X1 port map( A => n1704, B => lt_x_135_B_5_port, ZN => n2044);
   U1733 : NAND2_X1 port map( A1 => n2687, A2 => n2686, ZN => n3836);
   U1734 : NAND2_X1 port map( A1 => n1705, A2 => n2108, ZN => n2687);
   U1735 : XNOR2_X1 port map( A => n3642, B => n3841, ZN => n1705);
   U1736 : INV_X1 port map( A => n3642, ZN => n3480);
   U1737 : XNOR2_X1 port map( A => n1613, B => n3776, ZN => n1706);
   U1738 : BUF_X1 port map( A => n3662, Z => n1707);
   U1739 : AOI21_X1 port map( B1 => n1706, B2 => n2129, A => n3786, ZN => n1708
                           );
   U1740 : AND2_X1 port map( A1 => n1755, A2 => n2093, ZN => n1709);
   U1741 : AND2_X2 port map( A1 => n2075, A2 => n2027, ZN => n2245);
   U1742 : BUF_X1 port map( A => n3864, Z => n1710);
   U1743 : AND2_X2 port map( A1 => n2093, A2 => n2092, ZN => n2075);
   U1744 : NAND2_X1 port map( A1 => n2191, A2 => n2705, ZN => n1711);
   U1745 : AND2_X1 port map( A1 => n1730, A2 => n1758, ZN => n1712);
   U1746 : XNOR2_X1 port map( A => n3618, B => n2106, ZN => n1713);
   U1747 : XOR2_X1 port map( A => n3461, B => n2151, Z => n1714);
   U1748 : BUF_X1 port map( A => n2242, Z => n1748);
   U1749 : AND4_X2 port map( A1 => n2660, A2 => n2242, A3 => n2372, A4 => n2240
                           , ZN => n2093);
   U1750 : INV_X1 port map( A => n2232, ZN => n1715);
   U1751 : BUF_X1 port map( A => n2240, Z => n1716);
   U1752 : OR2_X1 port map( A1 => n3669, A2 => n2631, ZN => n2599);
   U1753 : NAND2_X1 port map( A1 => n2568, A2 => n2487, ZN => n1717);
   U1754 : OR2_X1 port map( A1 => n3294, A2 => n3234, ZN => n1718);
   U1755 : NOR2_X2 port map( A1 => n3330, A2 => n3329, ZN => n1719);
   U1756 : BUF_X2 port map( A => n3548, Z => n3223);
   U1757 : NAND4_X4 port map( A1 => n3500, A2 => n3499, A3 => n3498, A4 => 
                           n3497, ZN => DataP_alu_b_in_20_port);
   U1758 : INV_X1 port map( A => n2778, ZN => n1720);
   U1759 : CLKBUF_X3 port map( A => n3402, Z => n3216);
   U1760 : AOI21_X1 port map( B1 => n1617, B2 => n3826, A => n2704, ZN => n1721
                           );
   U1761 : INV_X1 port map( A => n2732, ZN => n1722);
   U1762 : BUF_X1 port map( A => n3763, Z => n1723);
   U1763 : OAI211_X1 port map( C1 => n2421, C2 => n2771, A => n1928, B => n1929
                           , ZN => DataP_alu_b_in_19_port);
   U1764 : OAI211_X1 port map( C1 => n2598, C2 => n2599, A => n2530, B => n2490
                           , ZN => n3763);
   U1765 : AND2_X1 port map( A1 => n3601, A2 => n2082, ZN => n1724);
   U1766 : AND2_X1 port map( A1 => n3601, A2 => n2082, ZN => n1725);
   U1767 : AND2_X1 port map( A1 => n3601, A2 => n2082, ZN => n2194);
   U1768 : BUF_X1 port map( A => n2735, Z => n1726);
   U1769 : AND4_X2 port map( A1 => n3321, A2 => n3322, A3 => n3319, A4 => n3320
                           , ZN => n3601);
   U1770 : NAND2_X1 port map( A1 => n1727, A2 => n3585, ZN => n3844);
   U1771 : NAND2_X1 port map( A1 => n3588, A2 => n3586, ZN => n1727);
   U1772 : NAND2_X1 port map( A1 => n1719, A2 => n3417, ZN => n3586);
   U1773 : NAND2_X1 port map( A1 => n1729, A2 => n3575, ZN => n3588);
   U1774 : XNOR2_X1 port map( A => n1926, B => n1728, ZN => n3417);
   U1775 : INV_X1 port map( A => n1716, ZN => n1728);
   U1776 : NAND2_X1 port map( A1 => n3574, A2 => n3577, ZN => n1729);
   U1777 : NAND2_X1 port map( A1 => n3415, A2 => n2232, ZN => n3575);
   U1778 : NAND2_X1 port map( A1 => n1730, A2 => n1758, ZN => n3849);
   U1779 : NAND2_X1 port map( A1 => n1731, A2 => n2108, ZN => n1730);
   U1780 : XNOR2_X1 port map( A => n1585, B => sra_131_SH_4_port, ZN => n1731);
   U1781 : AND2_X1 port map( A1 => n3459, A2 => DataP_alu_a_in_10_port, ZN => 
                           n1732);
   U1782 : BUF_X1 port map( A => n3572, Z => n1733);
   U1783 : OR2_X4 port map( A1 => n3404, A2 => n3403, ZN => 
                           DataP_alu_a_in_10_port);
   U1784 : INV_X4 port map( A => n2138, ZN => n2102);
   U1785 : BUF_X4 port map( A => sra_131_SH_4_port, Z => n2138);
   U1786 : NAND2_X1 port map( A1 => n2549, A2 => n2547, ZN => n1734);
   U1787 : NOR2_X1 port map( A1 => n3659, A2 => n1737, ZN => n1735);
   U1788 : INV_X1 port map( A => n2123, ZN => n1736);
   U1789 : NOR2_X1 port map( A1 => n3659, A2 => n1737, ZN => n3691);
   U1790 : OAI211_X1 port map( C1 => n2425, C2 => n1627, A => n1901, B => n1900
                           , ZN => DataP_alu_b_in_18_port);
   U1791 : OR2_X1 port map( A1 => DataP_alu_b_in_19_port, A2 => 
                           DataP_alu_b_in_18_port, ZN => n1737);
   U1792 : AND2_X1 port map( A1 => n2075, A2 => n2027, ZN => n1738);
   U1793 : NAND2_X1 port map( A1 => n3488, A2 => n3489, ZN => n1739);
   U1794 : BUF_X1 port map( A => n3588, Z => n1740);
   U1795 : INV_X1 port map( A => n3539, ZN => n1741);
   U1796 : INV_X1 port map( A => n3288, ZN => n1742);
   U1797 : NAND2_X1 port map( A1 => n2619, A2 => n1742, ZN => n1743);
   U1798 : AND2_X1 port map( A1 => DataP_alu_a_in_0_port, A2 => n2226, ZN => 
                           n3577);
   U1799 : NAND2_X1 port map( A1 => n1633, A2 => n2726, ZN => n1744);
   U1800 : AND2_X1 port map( A1 => n2612, A2 => n3632, ZN => n1745);
   U1801 : AND2_X1 port map( A1 => n3648, A2 => DataP_alu_a_in_19_port, ZN => 
                           n1746);
   U1802 : OAI21_X1 port map( B1 => n2044, B2 => n2128, A => n2163, ZN => n1747
                           );
   U1803 : NOR2_X1 port map( A1 => n3334, A2 => n3333, ZN => n2206);
   U1804 : BUF_X1 port map( A => n3834, Z => n1749);
   U1805 : INV_X1 port map( A => n1595, ZN => DataP_alu_b_in_2_port);
   U1806 : OR2_X4 port map( A1 => n3365, A2 => n3364, ZN => 
                           DataP_alu_a_in_25_port);
   U1807 : AND4_X2 port map( A1 => n3318, A2 => n3317, A3 => n3316, A4 => n3315
                           , ZN => n2082);
   U1808 : INV_X1 port map( A => DataP_alu_a_in_17_port, ZN => n1750);
   U1809 : BUF_X2 port map( A => DataP_alu_a_in_17_port, Z => n1751);
   U1810 : OAI21_X1 port map( B1 => n3216, B2 => n2440, A => n1840, ZN => 
                           DataP_alu_a_in_17_port);
   U1811 : INV_X1 port map( A => n3841, ZN => n1752);
   U1812 : NAND4_X1 port map( A1 => n3350, A2 => n3349, A3 => n3348, A4 => 
                           n3347, ZN => DataP_alu_b_in_8_port);
   U1813 : AND4_X2 port map( A1 => n3522, A2 => n3521, A3 => n3520, A4 => n3519
                           , ZN => n1753);
   U1814 : BUF_X1 port map( A => n3574, Z => n1754);
   U1815 : AND3_X1 port map( A1 => n1724, A2 => n2094, A3 => n1579, ZN => n2092
                           );
   U1816 : AND4_X2 port map( A1 => n2176, A2 => n2178, A3 => n2621, A4 => n2175
                           , ZN => n2780);
   U1817 : NAND2_X1 port map( A1 => n2615, A2 => n1756, ZN => n3649);
   U1818 : AND2_X1 port map( A1 => n2733, A2 => n2202, ZN => n1756);
   U1819 : INV_X1 port map( A => DataP_add_D_3_port, ZN => n1757);
   U1820 : NAND4_X1 port map( A1 => n3457, A2 => n3456, A3 => n3454, A4 => 
                           n3455, ZN => DataP_alu_b_in_11_port);
   U1821 : NAND2_X1 port map( A1 => n2380, A2 => n1698, ZN => n1758);
   U1822 : AOI21_X1 port map( B1 => n1632, B2 => n2129, A => n3795, ZN => n1759
                           );
   U1823 : OR2_X1 port map( A1 => n2141, A2 => n1762, ZN => n1761);
   U1824 : INV_X1 port map( A => n1573, ZN => n1762);
   U1825 : NOR2_X1 port map( A1 => n2371, A2 => n2108, ZN => n2390);
   U1826 : NAND4_X1 port map( A1 => n3325, A2 => n3326, A3 => n3324, A4 => 
                           n3323, ZN => DataP_alu_b_in_6_port);
   U1827 : OAI21_X1 port map( B1 => n3624, B2 => DataP_alu_b_in_15_port, A => 
                           n2145, ZN => n2329);
   U1828 : INV_X1 port map( A => n2068, ZN => n2043);
   U1829 : NOR2_X1 port map( A1 => n1761, A2 => n2145, ZN => n2675);
   U1830 : AOI211_X1 port map( C1 => n2279, C2 => n2278, A => n2277, B => n2348
                           , ZN => n2291);
   U1831 : NOR2_X1 port map( A1 => n2379, A2 => n2395, ZN => n2033);
   U1832 : AND3_X2 port map( A1 => n3531, A2 => n3530, A3 => n1963, ZN => n2371
                           );
   U1833 : NOR2_X1 port map( A1 => n2068, A2 => lt_x_135_B_12_port, ZN => n2042
                           );
   U1834 : XNOR2_X1 port map( A => n3620, B => n2145, ZN => n2685);
   U1835 : NAND2_X1 port map( A1 => n1647, A2 => n2041, ZN => n3620);
   U1836 : NOR2_X1 port map( A1 => n2068, A2 => n1761, ZN => n2041);
   U1837 : INV_X1 port map( A => n2108, ZN => n2128);
   U1838 : INV_X1 port map( A => n2016, ZN => n2014);
   U1839 : OR2_X2 port map( A1 => n3340, A2 => n3339, ZN => 
                           DataP_alu_a_in_5_port);
   U1840 : OR2_X2 port map( A1 => n3398, A2 => n3397, ZN => 
                           DataP_alu_a_in_12_port);
   U1841 : BUF_X1 port map( A => n1734, Z => n2167);
   U1842 : NAND2_X1 port map( A1 => n2040, A2 => n1968, ZN => n3608);
   U1843 : NAND2_X1 port map( A1 => n2680, A2 => n3886, ZN => n2039);
   U1844 : INV_X1 port map( A => n2052, ZN => n2048);
   U1845 : BUF_X1 port map( A => n3606, Z => n2156);
   U1846 : INV_X1 port map( A => DataP_a_out_27_port, ZN => n1977);
   U1847 : INV_X1 port map( A => DataP_a_out_29_port, ZN => n1978);
   U1848 : INV_X1 port map( A => DataP_a_out_26_port, ZN => n1979);
   U1849 : INV_X1 port map( A => DataP_a_out_28_port, ZN => n1980);
   U1850 : INV_X1 port map( A => DataP_a_out_1_port, ZN => n1981);
   U1851 : INV_X1 port map( A => DataP_a_out_7_port, ZN => n1982);
   U1852 : INV_X1 port map( A => DataP_a_out_10_port, ZN => n1983);
   U1853 : INV_X1 port map( A => DataP_a_out_11_port, ZN => n1984);
   U1854 : INV_X1 port map( A => DataP_a_out_12_port, ZN => n1985);
   U1855 : INV_X1 port map( A => DataP_a_out_13_port, ZN => n1986);
   U1856 : INV_X1 port map( A => DataP_a_out_14_port, ZN => n1987);
   U1857 : INV_X1 port map( A => DataP_a_out_15_port, ZN => n1988);
   U1858 : INV_X1 port map( A => DataP_a_out_30_port, ZN => n2001);
   U1859 : INV_X1 port map( A => DataP_a_out_3_port, ZN => n2002);
   U1860 : INV_X1 port map( A => DataP_a_out_4_port, ZN => n2003);
   U1861 : INV_X1 port map( A => DataP_a_out_5_port, ZN => n2004);
   U1862 : INV_X1 port map( A => DataP_a_out_6_port, ZN => n2005);
   U1863 : INV_X1 port map( A => CU_I_cw_10_port, ZN => n2007);
   U1864 : NAND2_X1 port map( A1 => n2063, A2 => n2065, ZN => n2560);
   U1865 : NAND2_X1 port map( A1 => n3777, A2 => n2066, ZN => n2065);
   U1866 : NAND3_X1 port map( A1 => n2034, A2 => n3432, A3 => n2290, ZN => 
                           n1763);
   U1867 : OAI211_X1 port map( C1 => n3562, C2 => n2391, A => n2016, B => n1763
                           , ZN => n2013);
   U1868 : AOI22_X1 port map( A1 => n3051, A2 => n2856, B1 => n2919, B2 => 
                           n2879, ZN => n1764);
   U1869 : AOI22_X1 port map( A1 => n2115, A2 => n2857, B1 => n2101, B2 => 
                           n1764, ZN => n1765);
   U1870 : MUX2_X1 port map( A => n1765, B => n2901, S => n2138, Z => 
                           DataP_ALU_C_shifter_N43);
   U1871 : INV_X1 port map( A => DataP_a_out_16_port, ZN => n1989);
   U1872 : NOR2_X1 port map( A1 => n3055, A2 => n2902, ZN => n1766);
   U1873 : OAI21_X1 port map( B1 => n3897, B2 => n3495, A => n3453, ZN => n1767
                           );
   U1874 : NOR2_X1 port map( A1 => n3450, A2 => n3489, ZN => n1768);
   U1875 : XNOR2_X1 port map( A => n1768, B => n3458, ZN => n1769);
   U1876 : OAI221_X1 port map( B1 => n2102, B2 => n3132, C1 => n1866, C2 => 
                           n3071, A => n3877, ZN => n1770);
   U1877 : INV_X1 port map( A => n3055, ZN => n1771);
   U1878 : OAI221_X1 port map( B1 => n3055, B2 => n2935, C1 => n1771, C2 => 
                           n2995, A => n3227, ZN => n1772);
   U1879 : OAI211_X1 port map( C1 => n3880, C2 => n1769, A => n1770, B => n1772
                           , ZN => n1773);
   U1880 : AOI211_X1 port map( C1 => n3228, C2 => n1766, A => n1767, B => n1773
                           , ZN => n340);
   U1881 : AOI211_X1 port map( C1 => n2301, C2 => DataP_alu_a_in_16_port, A => 
                           n2298, B => n2274, ZN => n1774);
   U1882 : AOI221_X1 port map( B1 => n2320, B2 => n2257, C1 => n2256, C2 => 
                           n2257, A => n2255, ZN => n1775);
   U1883 : AOI211_X1 port map( C1 => n2266, C2 => n2267, A => n2264, B => n2265
                           , ZN => n1776);
   U1884 : OAI21_X1 port map( B1 => n1775, B2 => n2268, A => n1776, ZN => n1777
                           );
   U1885 : NAND3_X1 port map( A1 => n2369, A2 => n1774, A3 => n1777, ZN => 
                           n2292);
   U1886 : AOI22_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_30_port, B1 =>
                           DataP_B_s_30_port, B2 => n2227, ZN => n1778);
   U1887 : OAI211_X1 port map( C1 => n2417, C2 => n2772, A => n3523, B => n1778
                           , ZN => DataP_alu_b_in_30_port);
   U1888 : OAI21_X1 port map( B1 => n2135, B2 => n3851, A => n3891, ZN => n1779
                           );
   U1889 : AOI22_X1 port map( A1 => DataP_alu_a_in_18_port, A2 => n3894, B1 => 
                           n1736, B2 => n1779, ZN => n1780);
   U1890 : NAND3_X1 port map( A1 => n3227, A2 => n3006, A3 => n2102, ZN => 
                           n1781);
   U1891 : OAI211_X1 port map( C1 => n3897, C2 => n3747, A => n1780, B => n1781
                           , ZN => n3748);
   U1892 : AOI22_X1 port map( A1 => n3052, A2 => n3033, B1 => n3034, B2 => 
                           n3051, ZN => n1782);
   U1893 : AOI22_X1 port map( A1 => n1782, A2 => n2101, B1 => n3035, B2 => 
                           n2112, ZN => n3037);
   U1894 : INV_X1 port map( A => DataP_a_out_17_port, ZN => n1990);
   U1895 : OAI21_X1 port map( B1 => n2102, B2 => n3198, A => n3194, ZN => n1783
                           );
   U1896 : AOI21_X1 port map( B1 => n2221, B2 => n3837, A => n3428, ZN => n1784
                           );
   U1897 : NAND2_X1 port map( A1 => n3443, A2 => n3483, ZN => n1785);
   U1898 : NOR2_X1 port map( A1 => n1784, A2 => n1785, ZN => n1786);
   U1899 : AOI211_X1 port map( C1 => n1784, C2 => n1785, A => n3880, B => n1786
                           , ZN => n1787);
   U1900 : NOR2_X1 port map( A1 => n3055, A2 => n2915, ZN => n1788);
   U1901 : AOI22_X1 port map( A1 => DataP_ALU_C_shifter_N59, A2 => n3227, B1 =>
                           n3228, B2 => n1788, ZN => n1789);
   U1902 : OAI211_X1 port map( C1 => n3897, C2 => n3494, A => n3437, B => n1789
                           , ZN => n1790);
   U1903 : AOI211_X1 port map( C1 => n3877, C2 => n1783, A => n1787, B => n1790
                           , ZN => n341);
   U1904 : NAND2_X1 port map( A1 => n3569, A2 => ALU_OPCODE_i_0_port, ZN => 
                           n1791);
   U1905 : AOI21_X1 port map( B1 => n2034, B2 => n2290, A => n1791, ZN => n1792
                           );
   U1906 : NOR3_X1 port map( A1 => n1792, A2 => n1964, A3 => n2033, ZN => n2032
                           );
   U1907 : INV_X1 port map( A => DataP_a_out_18_port, ZN => n1991);
   U1908 : OAI21_X1 port map( B1 => n3206, B2 => n3197, A => n3190, ZN => n1793
                           );
   U1909 : OAI22_X1 port map( A1 => n3841, A2 => n3842, B1 => n2110, B2 => 
                           n3840, ZN => n1794);
   U1910 : INV_X1 port map( A => n3055, ZN => n1795);
   U1911 : OAI221_X1 port map( B1 => n3055, B2 => n3041, C1 => n1795, C2 => 
                           n3040, A => n3900, ZN => n1796);
   U1912 : NOR2_X1 port map( A1 => n2138, A2 => n2914, ZN => n1797);
   U1913 : XNOR2_X1 port map( A => DataP_alu_a_in_8_port, B => n2204, ZN => 
                           n1798);
   U1914 : AOI21_X1 port map( B1 => n3835, B2 => n2221, A => n3837, ZN => n1799
                           );
   U1915 : AOI211_X1 port map( C1 => n3837, C2 => n1798, A => n1799, B => n3880
                           , ZN => n1800);
   U1916 : AOI21_X1 port map( B1 => n3228, B2 => n1797, A => n1800, ZN => n1801
                           );
   U1917 : NAND2_X1 port map( A1 => n1796, A2 => n1801, ZN => n1802);
   U1918 : AOI211_X1 port map( C1 => n3877, C2 => n1793, A => n1794, B => n1802
                           , ZN => n345);
   U1919 : AOI22_X1 port map( A1 => n3697, A2 => DataP_alu_b_in_27_port, B1 => 
                           n2354, B2 => DataP_alu_b_in_26_port, ZN => n1803);
   U1920 : INV_X1 port map( A => n2355, ZN => n1804);
   U1921 : AOI221_X1 port map( B1 => n2356, B2 => n1803, C1 => n2367, C2 => 
                           n1803, A => n1804, ZN => n2359);
   U1922 : OAI21_X1 port map( B1 => DataP_alu_a_in_16_port, B2 => 
                           DataP_alu_b_in_16_port, A => n3894, ZN => n1805);
   U1923 : NAND3_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => 
                           DataP_alu_b_in_16_port, A3 => n3890, ZN => n1806);
   U1924 : OAI211_X1 port map( C1 => n3731, C2 => n3897, A => n1805, B => n1806
                           , ZN => n3732);
   U1925 : AOI22_X1 port map( A1 => n3189, A2 => n3205, B1 => n2101, B2 => 
                           n3188, ZN => n1807);
   U1926 : NAND2_X1 port map( A1 => n3206, A2 => n1807, ZN => n3190);
   U1927 : INV_X1 port map( A => DataP_a_out_19_port, ZN => n1992);
   U1928 : XOR2_X1 port map( A => n3854, B => n2203, Z => n1808);
   U1929 : INV_X1 port map( A => n3055, ZN => n1809);
   U1930 : OAI221_X1 port map( B1 => n3055, B2 => n3032, C1 => n1809, C2 => 
                           n3031, A => n3900, ZN => n1810);
   U1931 : OAI21_X1 port map( B1 => n2102, B2 => n3181, A => n3180, ZN => n1811
                           );
   U1932 : NAND2_X1 port map( A1 => n1811, A2 => n3877, ZN => n1812);
   U1933 : OAI211_X1 port map( C1 => n1808, C2 => n3880, A => n1810, B => n1812
                           , ZN => n1813);
   U1934 : AOI21_X1 port map( B1 => n3894, B2 => DataP_alu_a_in_6_port, A => 
                           n3858, ZN => n1814);
   U1935 : NAND3_X1 port map( A1 => n3228, A2 => n2898, A3 => n1809, ZN => 
                           n1815);
   U1936 : OAI211_X1 port map( C1 => n3897, C2 => n3859, A => n1814, B => n1815
                           , ZN => n1816);
   U1937 : NOR2_X1 port map( A1 => n1813, A2 => n1816, ZN => n353);
   U1938 : NOR2_X1 port map( A1 => DataP_alu_a_in_18_port, A2 => n2341, ZN => 
                           n1817);
   U1939 : AOI22_X1 port map( A1 => n1722, A2 => n2202, B1 => n1736, B2 => 
                           n1817, ZN => n2346);
   U1940 : NAND3_X1 port map( A1 => n1574, A2 => n2120, A3 => n3726, ZN => 
                           n1818);
   U1941 : NAND2_X1 port map( A1 => n1818, A2 => n1694, ZN => n1819);
   U1942 : XNOR2_X1 port map( A => n1819, B => n2125, ZN => n3728);
   U1943 : OAI211_X1 port map( C1 => n3800, C2 => n3897, A => n1820, B => n1821
                           , ZN => n3801);
   U1944 : INV_X1 port map( A => DataP_a_out_20_port, ZN => n1993);
   U1945 : NOR2_X1 port map( A1 => n3055, A2 => n2912, ZN => n1822);
   U1946 : NAND2_X1 port map( A1 => n2215, A2 => n2156, ZN => n1823);
   U1947 : XNOR2_X1 port map( A => n1823, B => n3607, ZN => n1824);
   U1948 : OAI21_X1 port map( B1 => n3206, B2 => n3174, A => n3173, ZN => n1825
                           );
   U1949 : NAND2_X1 port map( A1 => n1825, A2 => n3877, ZN => n1826);
   U1950 : OAI21_X1 port map( B1 => n3880, B2 => n1824, A => n1826, ZN => n1827
                           );
   U1951 : OAI221_X1 port map( B1 => n2138, B2 => n3026, C1 => n1908, C2 => 
                           n3025, A => n3227, ZN => n1828);
   U1952 : OAI211_X1 port map( C1 => n3603, C2 => n3897, A => n3602, B => n1828
                           , ZN => n1829);
   U1953 : AOI211_X1 port map( C1 => n3228, C2 => n1822, A => n1827, B => n1829
                           , ZN => n354);
   U1954 : NAND2_X1 port map( A1 => n1694, A2 => n2031, ZN => n1830);
   U1955 : XNOR2_X1 port map( A => n1830, B => n2030, ZN => n3427);
   U1956 : AOI22_X1 port map( A1 => DataP_alu_out_W_27_port, A2 => n3207, B1 =>
                           DataP_alu_out_M_27_port, B2 => n3211, ZN => n1831);
   U1957 : OAI21_X1 port map( B1 => n3213, B2 => n145, A => n1831, ZN => n1832)
                           ;
   U1958 : NOR2_X1 port map( A1 => n3217, A2 => n2438, ZN => n1833);
   U1959 : NOR2_X2 port map( A1 => n1832, A2 => n1833, ZN => n3697);
   U1960 : AOI22_X1 port map( A1 => n3219, A2 => DataP_B_s_22_port, B1 => n1581
                           , B2 => DataP_IMM_s_22_port, ZN => n1834);
   U1961 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_22_port, ZN =>
                           n1835);
   U1962 : OAI211_X1 port map( C1 => n2428, C2 => n2772, A => n1834, B => n1835
                           , ZN => DataP_alu_b_in_22_port);
   U1963 : AOI21_X1 port map( B1 => n3890, B2 => n3048, A => n3894, ZN => n1836
                           );
   U1964 : OAI22_X1 port map( A1 => n3891, A2 => n3047, B1 => n1715, B2 => 
                           n1836, ZN => n3578);
   U1965 : INV_X1 port map( A => DataP_a_out_21_port, ZN => n1994);
   U1966 : OAI21_X1 port map( B1 => DataP_alu_b_in_15_port, B2 => n2210, A => 
                           n2145, ZN => n1837);
   U1967 : OAI22_X1 port map( A1 => DataP_alu_a_in_14_port, A2 => n1837, B1 => 
                           DataP_alu_a_in_15_port, B2 => n2230, ZN => n2264);
   U1968 : INV_X1 port map( A => n1725, ZN => n1838);
   U1969 : INV_X1 port map( A => n3214, ZN => n1839);
   U1970 : AOI222_X1 port map( A1 => n1606, A2 => n1839, B1 => 
                           DataP_alu_out_M_17_port, B2 => n2209, C1 => n3207, 
                           C2 => DataP_alu_out_W_17_port, ZN => n1840);
   U1971 : AOI22_X1 port map( A1 => n3219, A2 => DataP_B_s_24_port, B1 => n1581
                           , B2 => DataP_IMM_s_24_port, ZN => n1841);
   U1972 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_24_port, ZN =>
                           n1842);
   U1973 : NAND2_X1 port map( A1 => n2026, A2 => n1694, ZN => n1843);
   U1974 : XNOR2_X1 port map( A => n3429, B => n1843, ZN => n2011);
   U1975 : INV_X1 port map( A => DataP_a_out_22_port, ZN => n1995);
   U1976 : NOR2_X1 port map( A1 => n2138, A2 => n2911, ZN => n1844);
   U1977 : XNOR2_X1 port map( A => DataP_alu_a_in_4_port, B => n3849, ZN => 
                           n1845);
   U1978 : XNOR2_X1 port map( A => n1845, B => n3850, ZN => n1846);
   U1979 : OAI21_X1 port map( B1 => n2102, B2 => n3167, A => n3166, ZN => n1847
                           );
   U1980 : NAND2_X1 port map( A1 => n1847, A2 => n3877, ZN => n1848);
   U1981 : OAI21_X1 port map( B1 => n3880, B2 => n1846, A => n1848, ZN => n1849
                           );
   U1982 : AOI22_X1 port map( A1 => n2138, A2 => n3894, B1 => 
                           DataP_alu_a_in_4_port, B2 => n3852, ZN => n1850);
   U1983 : INV_X1 port map( A => n3055, ZN => n1851);
   U1984 : OAI221_X1 port map( B1 => n3055, B2 => n3020, C1 => n1851, C2 => 
                           n3019, A => n3900, ZN => n1852);
   U1985 : OAI211_X1 port map( C1 => n3853, C2 => n3897, A => n1850, B => n1852
                           , ZN => n1853);
   U1986 : AOI211_X1 port map( C1 => n3228, C2 => n1844, A => n1849, B => n1853
                           , ZN => n355);
   U1987 : AND3_X1 port map( A1 => n2123, A2 => n1722, A3 => n2108, ZN => n2617
                           );
   U1988 : NAND3_X1 port map( A1 => n1647, A2 => n2043, A3 => n2675, ZN => 
                           n1854);
   U1989 : XNOR2_X1 port map( A => n1854, B => n2230, ZN => n3616);
   U1990 : INV_X1 port map( A => n2535, ZN => n1855);
   U1991 : NAND2_X1 port map( A1 => n2213, A2 => n1855, ZN => n1856);
   U1992 : XNOR2_X1 port map( A => DataP_alu_b_in_20_port, B => n1856, ZN => 
                           n3666);
   U1993 : AOI22_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_29_port, B1 =>
                           n2782, B2 => DataP_alu_out_M_29_port, ZN => n1857);
   U1994 : NAND2_X1 port map( A1 => DataP_B_s_29_port, A2 => n2227, ZN => n1858
                           );
   U1995 : NAND3_X1 port map( A1 => n1858, A2 => n1857, A3 => n3523, ZN => 
                           DataP_alu_b_in_29_port);
   U1996 : OAI21_X1 port map( B1 => n2074, B2 => n3851, A => n3891, ZN => n1859
                           );
   U1997 : AOI22_X1 port map( A1 => lt_x_135_B_5_port, A2 => n3894, B1 => 
                           DataP_alu_a_in_5_port, B2 => n1859, ZN => n3602);
   U1998 : INV_X1 port map( A => DataP_a_out_23_port, ZN => n1996);
   U1999 : OAI211_X1 port map( C1 => n3872, C2 => n3897, A => n3871, B => n3870
                           , ZN => n1860);
   U2000 : NOR2_X1 port map( A1 => n3055, A2 => n2905, ZN => n1861);
   U2001 : AOI21_X1 port map( B1 => n1861, B2 => n3228, A => n1860, ZN => n1862
                           );
   U2002 : NOR2_X1 port map( A1 => n3861, A2 => n3862, ZN => n1863);
   U2003 : OAI211_X1 port map( C1 => n3868, C2 => n3867, A => n3866, B => n2208
                           , ZN => n1864);
   U2004 : OAI211_X1 port map( C1 => n1863, C2 => n2214, A => n2129, B => n1864
                           , ZN => n1865);
   U2005 : INV_X1 port map( A => n2102, ZN => n1866);
   U2006 : OAI221_X1 port map( B1 => n2102, B2 => n3138, C1 => n1866, C2 => 
                           n3088, A => n3877, ZN => n1867);
   U2007 : OAI221_X1 port map( B1 => n2138, B2 => n2953, C1 => n1888, C2 => 
                           n2998, A => n3227, ZN => n1868);
   U2008 : AND4_X1 port map( A1 => n1862, A2 => n1865, A3 => n1867, A4 => n1868
                           , ZN => n333);
   U2009 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_19_port, B1 =>
                           DataP_alu_out_W_19_port, B2 => n3207, ZN => n1869);
   U2010 : OAI21_X1 port map( B1 => n113, B2 => n3213, A => n1869, ZN => n3382)
                           ;
   U2011 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_30_port, B1 => 
                           DataP_alu_a_in_31_port, B2 => n2916, ZN => n1870);
   U2012 : AOI22_X1 port map( A1 => n2105, A2 => n1870, B1 => n2891, B2 => 
                           n2917, ZN => n1871);
   U2013 : AOI22_X1 port map( A1 => n3202, A2 => n2892, B1 => n1871, B2 => 
                           n3053, ZN => n1872);
   U2014 : AOI22_X1 port map( A1 => n2115, A2 => n2893, B1 => n2101, B2 => 
                           n1872, ZN => n1873);
   U2015 : MUX2_X1 port map( A => n1873, B => n2894, S => n3055, Z => 
                           DataP_ALU_C_shifter_N49);
   U2016 : INV_X1 port map( A => n3055, ZN => n1874);
   U2017 : NAND3_X1 port map( A1 => n3904, A2 => n2810, A3 => n1874, ZN => 
                           n3558);
   U2018 : AOI22_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_28_port, B1 =>
                           DataP_B_s_28_port, B2 => n2227, ZN => n1875);
   U2019 : OAI211_X1 port map( C1 => n2426, C2 => n1627, A => n3523, B => n1875
                           , ZN => DataP_alu_b_in_28_port);
   U2020 : AOI22_X1 port map( A1 => n3052, A2 => n3016, B1 => n3017, B2 => 
                           n3202, ZN => n1876);
   U2021 : AOI22_X1 port map( A1 => n1876, A2 => n2101, B1 => n3018, B2 => 
                           n2112, ZN => n3020);
   U2022 : NAND3_X1 port map( A1 => DataP_alu_a_in_14_port, A2 => n2145, A3 => 
                           n3890, ZN => n1877);
   U2023 : OAI21_X1 port map( B1 => DataP_alu_a_in_14_port, B2 => n2145, A => 
                           n3894, ZN => n1878);
   U2024 : OAI211_X1 port map( C1 => n3875, C2 => n3897, A => n1877, B => n1878
                           , ZN => n3876);
   U2025 : INV_X1 port map( A => DataP_a_out_24_port, ZN => n1997);
   U2026 : OAI21_X1 port map( B1 => n2102, B2 => n3160, A => n3159, ZN => n1879
                           );
   U2027 : INV_X1 port map( A => n3228, ZN => n1880);
   U2028 : NOR3_X1 port map( A1 => n3055, A2 => n2910, A3 => n1880, ZN => n1881
                           );
   U2029 : AOI22_X1 port map( A1 => n1973, A2 => n3846, B1 => 
                           DataP_alu_b_in_3_port, B2 => n3894, ZN => n1882);
   U2030 : OAI211_X1 port map( C1 => n3897, C2 => n3848, A => n3847, B => n1882
                           , ZN => n1883);
   U2031 : AOI211_X1 port map( C1 => n3877, C2 => n1879, A => n1881, B => n1883
                           , ZN => n1884);
   U2032 : AOI22_X1 port map( A1 => n3049, A2 => n3013, B1 => n3047, B2 => 
                           n3012, ZN => n1885);
   U2033 : AOI22_X1 port map( A1 => n3202, A2 => n3033, B1 => n3052, B2 => 
                           n1885, ZN => n1886);
   U2034 : AOI22_X1 port map( A1 => n2101, A2 => n1886, B1 => n3014, B2 => 
                           n3204, ZN => n1887);
   U2035 : INV_X1 port map( A => n3055, ZN => n1888);
   U2036 : OAI221_X1 port map( B1 => n3055, B2 => n1887, C1 => n1888, C2 => 
                           n3015, A => n3227, ZN => n1889);
   U2037 : AND2_X1 port map( A1 => n1884, A2 => n1889, ZN => n356);
   U2038 : NAND2_X1 port map( A1 => n2208, A2 => n3863, ZN => n1890);
   U2039 : XOR2_X1 port map( A => n1710, B => n1890, Z => n1891);
   U2040 : OAI21_X1 port map( B1 => n3206, B2 => n2997, A => n2942, ZN => n1892
                           );
   U2041 : OAI211_X1 port map( C1 => n3496, C2 => n3897, A => n3493, B => n3492
                           , ZN => n1893);
   U2042 : AOI21_X1 port map( B1 => n3227, B2 => n1892, A => n1893, ZN => n1894
                           );
   U2043 : OAI221_X1 port map( B1 => n2102, B2 => n3136, C1 => n1866, C2 => 
                           n3078, A => n3877, ZN => n1895);
   U2044 : OAI211_X1 port map( C1 => n3880, C2 => n1891, A => n1894, B => n1895
                           , ZN => n1896);
   U2045 : NOR2_X1 port map( A1 => n3055, A2 => n2904, ZN => n1897);
   U2046 : AOI21_X1 port map( B1 => n1897, B2 => n3228, A => n1896, ZN => n337)
                           ;
   U2047 : INV_X1 port map( A => n2381, ZN => n1898);
   U2048 : NAND2_X1 port map( A1 => n2614, A2 => n1898, ZN => n2385);
   U2049 : INV_X1 port map( A => n2209, ZN => n1899);
   U2050 : OAI222_X1 port map( A1 => n2433, A2 => n1899, B1 => n3213, B2 => n97
                           , C1 => n2072, C2 => n2516, ZN => n2693);
   U2051 : AOI22_X1 port map( A1 => n1631, A2 => DataP_B_s_18_port, B1 => n1623
                           , B2 => DataP_IMM_s_18_port, ZN => n1900);
   U2052 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_18_port, ZN =>
                           n1901);
   U2053 : OAI211_X1 port map( C1 => n2772, C2 => n2478, A => n2661, B => n2662
                           , ZN => n1902);
   U2054 : INV_X1 port map( A => n1902, ZN => n2660);
   U2055 : NAND2_X1 port map( A1 => n1597, A2 => n2108, ZN => n1903);
   U2056 : NAND3_X1 port map( A1 => n1903, A2 => DataP_alu_a_in_12_port, A3 => 
                           n2739, ZN => n3865);
   U2057 : NOR2_X1 port map( A1 => n2744, A2 => n3826, ZN => n1904);
   U2058 : INV_X1 port map( A => n4183, ZN => n1905);
   U2059 : AOI221_X1 port map( B1 => n4184, B2 => n4183, C1 => n3907, C2 => 
                           n1905, A => n4182, ZN => DataP_wrong_br);
   U2060 : OAI21_X1 port map( B1 => n1613, B2 => n2067, A => n2064, ZN => n1906
                           );
   U2061 : INV_X1 port map( A => n1906, ZN => n2063);
   U2062 : AOI22_X1 port map( A1 => n2101, A2 => n2857, B1 => n2858, B2 => 
                           n2115, ZN => n1907);
   U2063 : INV_X1 port map( A => n3055, ZN => n1908);
   U2064 : OAI221_X1 port map( B1 => n3055, B2 => n1907, C1 => n1908, C2 => 
                           n2827, A => n3228, ZN => n3743);
   U2065 : INV_X1 port map( A => DataP_a_out_25_port, ZN => n1998);
   U2066 : NOR2_X1 port map( A1 => n3055, A2 => n2913, ZN => n1909);
   U2067 : OAI21_X1 port map( B1 => n3854, B2 => n3610, A => n1648, ZN => n1910
                           );
   U2068 : OAI21_X1 port map( B1 => n2102, B2 => n3196, A => n3187, ZN => n1911
                           );
   U2069 : NAND2_X1 port map( A1 => n1911, A2 => n3877, ZN => n1912);
   U2070 : XOR2_X1 port map( A => n1910, B => n2211, Z => n1913);
   U2071 : OAI21_X1 port map( B1 => n1913, B2 => n3880, A => n1912, ZN => n1914
                           );
   U2072 : AOI22_X1 port map( A1 => DataP_alu_a_in_7_port, A2 => n3894, B1 => 
                           DataP_alu_b_in_7_port, B2 => n3612, ZN => n1915);
   U2073 : INV_X1 port map( A => n3055, ZN => n1916);
   U2074 : OAI221_X1 port map( B1 => n3055, B2 => n3037, C1 => n1916, C2 => 
                           n3036, A => n3227, ZN => n1917);
   U2075 : OAI211_X1 port map( C1 => n3897, C2 => n3613, A => n1915, B => n1917
                           , ZN => n1918);
   U2076 : NOR2_X1 port map( A1 => n2119, A2 => n1973, ZN => n1919);
   U2077 : NAND3_X1 port map( A1 => n2254, A2 => n2080, A3 => n2081, ZN => 
                           n1920);
   U2078 : OAI21_X1 port map( B1 => DataP_alu_a_in_2_port, B2 => n2315, A => 
                           n1920, ZN => n1921);
   U2079 : OAI22_X1 port map( A1 => n1919, A2 => n1921, B1 => lt_x_135_B_5_port
                           , B2 => n2113, ZN => n1922);
   U2080 : NAND2_X1 port map( A1 => DataP_alu_a_in_26_port, A2 => n2127, ZN => 
                           n1923);
   U2081 : OAI21_X1 port map( B1 => n3697, B2 => DataP_alu_b_in_27_port, A => 
                           n1923, ZN => n2297);
   U2082 : NAND4_X1 port map( A1 => n4108, A2 => n3782, A3 => n3771, A4 => 
                           n4109, ZN => n2743);
   U2083 : INV_X1 port map( A => DataP_alu_a_in_25_port, ZN => n1924);
   U2084 : AOI21_X1 port map( B1 => n2586, B2 => n2585, A => n1924, ZN => n3798
                           );
   U2085 : INV_X1 port map( A => n2108, ZN => n1925);
   U2086 : NOR2_X1 port map( A1 => n1925, A2 => n3416, ZN => n1926);
   U2087 : AOI21_X1 port map( B1 => n2128, B2 => n2739, A => 
                           DataP_alu_a_in_12_port, ZN => n2735);
   U2088 : INV_X1 port map( A => n2241, ZN => n1927);
   U2089 : NOR2_X1 port map( A1 => n3725, A2 => n1927, ZN => n2432);
   U2090 : AOI22_X1 port map( A1 => n1631, A2 => DataP_B_s_19_port, B1 => n1623
                           , B2 => DataP_IMM_s_19_port, ZN => n1928);
   U2091 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_19_port, ZN =>
                           n1929);
   U2092 : INV_X1 port map( A => n3680, ZN => n1930);
   U2093 : AOI21_X1 port map( B1 => n2378, B2 => n1930, A => n1707, ZN => n2674
                           );
   U2094 : INV_X1 port map( A => n3688, ZN => n1931);
   U2095 : NOR2_X1 port map( A1 => n1931, A2 => n2133, ZN => n1932);
   U2096 : AOI22_X1 port map( A1 => n1931, A2 => n2133, B1 => n3672, B2 => 
                           n1932, ZN => n2064);
   U2097 : AOI21_X1 port map( B1 => n2102, B2 => n3150, A => n3195, ZN => n1933
                           );
   U2098 : OAI211_X1 port map( C1 => n3707, C2 => n3897, A => n3706, B => n3705
                           , ZN => n1934);
   U2099 : AOI21_X1 port map( B1 => n3227, B2 => DataP_ALU_C_shifter_N80, A => 
                           n1934, ZN => n1935);
   U2100 : AOI22_X1 port map( A1 => n3202, A2 => n2888, B1 => n2918, B2 => 
                           n2887, ZN => n1936);
   U2101 : AOI22_X1 port map( A1 => n2115, A2 => n2889, B1 => n2101, B2 => 
                           n1936, ZN => n1937);
   U2102 : OAI221_X1 port map( B1 => n2138, B2 => n1937, C1 => n1916, C2 => 
                           n2890, A => n3904, ZN => n1938);
   U2103 : OAI211_X1 port map( C1 => n3892, C2 => n1933, A => n1935, B => n1938
                           , ZN => n2756);
   U2104 : INV_X1 port map( A => DataP_a_out_0_port, ZN => n1999);
   U2105 : NOR2_X1 port map( A1 => n3788, A2 => n2744, ZN => n2389);
   U2106 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_9_port, B1 => 
                           n3207, B2 => DataP_alu_out_W_9_port, ZN => n1939);
   U2107 : NAND2_X1 port map( A1 => n2139, A2 => DataP_npc_E_9_port, ZN => 
                           n1940);
   U2108 : OAI211_X1 port map( C1 => n3216, C2 => n2435, A => n1939, B => n1940
                           , ZN => DataP_alu_a_in_9_port);
   U2109 : XOR2_X1 port map( A => lt_x_135_B_12_port, B => n1941, Z => n3481);
   U2110 : OAI211_X1 port map( C1 => n2685, C2 => n2128, A => n2651, B => n2652
                           , ZN => n3631);
   U2111 : OAI221_X1 port map( B1 => n3195, B2 => n3101, C1 => n3195, C2 => 
                           n2102, A => n3877, ZN => n3734);
   U2112 : AOI22_X1 port map( A1 => n3051, A2 => n2861, B1 => n2918, B2 => 
                           n2888, ZN => n1942);
   U2113 : AOI22_X1 port map( A1 => n2101, A2 => n1942, B1 => n2862, B2 => 
                           n2115, ZN => n1943);
   U2114 : INV_X1 port map( A => n3055, ZN => n1944);
   U2115 : OAI221_X1 port map( B1 => n3055, B2 => n1943, C1 => n1944, C2 => 
                           n2863, A => n3228, ZN => n3814);
   U2116 : INV_X1 port map( A => n3417, ZN => n1945);
   U2117 : NAND2_X1 port map( A1 => DataP_alu_a_in_2_port, A2 => n1945, ZN => 
                           n3585);
   U2118 : NOR3_X1 port map( A1 => n4005, A2 => IR_CU_4_port, A3 => 
                           IR_CU_5_port, ZN => n1946);
   U2119 : AOI21_X1 port map( B1 => n3996, B2 => n607, A => n1946, ZN => n1947)
                           ;
   U2120 : OAI221_X1 port map( B1 => n4036, B2 => n4027, C1 => n4036, C2 => 
                           n4016, A => n1947, ZN => n4006);
   U2121 : AOI21_X1 port map( B1 => n2432, B2 => n2766, A => n2765, ZN => n1948
                           );
   U2122 : NOR2_X1 port map( A1 => n2746, A2 => n1948, ZN => n2719);
   U2123 : OAI21_X1 port map( B1 => n2234, B2 => n2673, A => n2674, ZN => n1949
                           );
   U2124 : OAI21_X1 port map( B1 => n3682, B2 => n1949, A => n2167, ZN => n3650
                           );
   U2125 : INV_X1 port map( A => DataP_a_out_31_port, ZN => n2006);
   U2126 : NAND2_X1 port map( A1 => n3964, A2 => n3965, ZN => n1950);
   U2127 : NOR3_X1 port map( A1 => n3969, A2 => n3970, A3 => n3971, ZN => n1951
                           );
   U2128 : NAND4_X1 port map( A1 => n3972, A2 => n3973, A3 => n3968, A4 => 
                           n1951, ZN => n1952);
   U2129 : NOR4_X1 port map( A1 => n3966, A2 => n3967, A3 => n1950, A4 => n1952
                           , ZN => n1953);
   U2130 : INV_X1 port map( A => n3956, ZN => n1954);
   U2131 : NAND4_X1 port map( A1 => n3957, A2 => n3958, A3 => n3959, A4 => 
                           n1954, ZN => n1955);
   U2132 : NOR2_X1 port map( A1 => n3954, A2 => n3955, ZN => n1956);
   U2133 : NAND3_X1 port map( A1 => n3953, A2 => n3952, A3 => n1956, ZN => 
                           n1957);
   U2134 : NOR4_X1 port map( A1 => n3960, A2 => n3961, A3 => n1955, A4 => n1957
                           , ZN => n1958);
   U2135 : NAND4_X1 port map( A1 => n3962, A2 => n3963, A3 => n1953, A4 => 
                           n1958, ZN => n1959);
   U2136 : NAND2_X1 port map( A1 => n3974, A2 => n1959, ZN => DataP_NPC_add_N0)
                           ;
   U2137 : INV_X1 port map( A => n2108, ZN => n2535);
   U2138 : INV_X2 port map( A => n3051, ZN => n2919);
   U2139 : INV_X2 port map( A => n3051, ZN => n2918);
   U2140 : INV_X1 port map( A => n2073, ZN => DataP_alu_a_in_31_port);
   U2141 : INV_X1 port map( A => n2380, ZN => sra_131_SH_4_port);
   U2142 : INV_X2 port map( A => n2138, ZN => n3206);
   U2143 : AND3_X1 port map( A1 => n4061, A2 => n4060, A3 => n4059, ZN => n1961
                           );
   U2144 : BUF_X4 port map( A => DataP_alu_b_in_2_port, Z => n3202);
   U2145 : CLKBUF_X3 port map( A => n3203, Z => n3051);
   U2146 : INV_X4 port map( A => n3046, ZN => n2103);
   U2147 : OR2_X1 port map( A1 => n2578, A2 => n3327, ZN => 
                           DataP_alu_a_in_3_port);
   U2148 : OR2_X4 port map( A1 => n3356, A2 => n3355, ZN => 
                           DataP_alu_a_in_29_port);
   U2149 : AND2_X1 port map( A1 => n3529, A2 => n3528, ZN => n1963);
   U2150 : OR2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => n2672, ZN => n1964
                           );
   U2151 : OR2_X2 port map( A1 => n3385, A2 => n3384, ZN => 
                           DataP_alu_a_in_18_port);
   U2152 : OR2_X2 port map( A1 => n3377, A2 => n3376, ZN => 
                           DataP_alu_a_in_21_port);
   U2153 : OR2_X1 port map( A1 => n4110, A2 => n4199, ZN => n1966);
   U2154 : NAND2_X2 port map( A1 => n3433, A2 => n3561, ZN => n3886);
   U2155 : AND2_X1 port map( A1 => n2355, A2 => n2306, ZN => n1967);
   U2156 : AND2_X1 port map( A1 => DataP_alu_a_in_6_port, A2 => n2039, ZN => 
                           n1968);
   U2157 : OR2_X1 port map( A1 => n3269, A2 => n3270, ZN => n1970);
   U2158 : AND2_X1 port map( A1 => n2066, A2 => n2062, ZN => n1971);
   U2159 : OR2_X1 port map( A1 => n2067, A2 => n2708, ZN => n1972);
   U2160 : NOR2_X4 port map( A1 => n3235, A2 => n2104, ZN => n36);
   U2161 : INV_X1 port map( A => CU_I_aluOpcode_i_4_port, ZN => n2000);
   U2162 : BUF_X2 port map( A => DataP_alu_a_in_3_port, Z => n1973);
   U2163 : INV_X1 port map( A => DataP_add_S2_2_port, ZN => n1974);
   n1975 <= '1';
   n1976 <= '1';
   U2166 : NAND2_X1 port map( A1 => n2009, A2 => n3479, ZN => n3641);
   U2167 : NOR2_X1 port map( A1 => DataP_alu_b_in_8_port, A2 => 
                           DataP_alu_b_in_9_port, ZN => n2009);
   U2168 : NAND2_X1 port map( A1 => n2010, A2 => n3483, ZN => n3485);
   U2169 : OR2_X2 port map( A1 => n2011, A2 => n2099, ZN => n3483);
   U2170 : NAND2_X1 port map( A1 => n3834, A2 => n3443, ZN => n2010);
   U2171 : NAND2_X1 port map( A1 => n2011, A2 => n2099, ZN => n3443);
   U2172 : NAND2_X1 port map( A1 => n3836, A2 => n2110, ZN => n3834);
   U2173 : NAND2_X1 port map( A1 => DataP_ALU_C_comp_N24, A2 => n2012, ZN => 
                           n2016);
   U2174 : AND2_X1 port map( A1 => n3561, A2 => n2391, ZN => n2012);
   U2175 : OAI211_X1 port map( C1 => n2017, C2 => n2014, A => n2013, B => n2015
                           , ZN => n3567);
   U2176 : NOR2_X1 port map( A1 => n3571, A2 => n2379, ZN => n2015);
   U2177 : NAND2_X1 port map( A1 => DataP_ALU_C_comp_N50, A2 => 
                           ALU_OPCODE_i_2_port, ZN => n2017);
   U2178 : NAND2_X1 port map( A1 => n2018, A2 => n2361, ZN => 
                           DataP_ALU_C_comp_N50);
   U2179 : NAND2_X1 port map( A1 => n2019, A2 => n1967, ZN => n2018);
   U2180 : NAND2_X1 port map( A1 => n2363, A2 => n2362, ZN => n2019);
   U2181 : AND2_X1 port map( A1 => n2594, A2 => n2593, ZN => n2576);
   U2182 : NAND2_X1 port map( A1 => n2664, A2 => n2020, ZN => n2594);
   U2183 : AND2_X1 port map( A1 => n2710, A2 => n2720, ZN => n2020);
   U2184 : NAND2_X1 port map( A1 => n2021, A2 => n2750, ZN => n2720);
   U2185 : OAI211_X1 port map( C1 => n2025, C2 => n1574, A => n2024, B => n2022
                           , ZN => n2190);
   U2186 : INV_X1 port map( A => n2023, ZN => n2022);
   U2187 : OAI21_X1 port map( B1 => n2485, B2 => n2025, A => n2722, ZN => n2023
                           );
   U2188 : NAND4_X1 port map( A1 => n3709, A2 => n2485, A3 => 
                           DataP_alu_b_in_26_port, A4 => n2108, ZN => n2024);
   U2189 : NAND2_X1 port map( A1 => n2127, A2 => n2108, ZN => n2025);
   U2190 : NAND2_X1 port map( A1 => n2075, A2 => n3841, ZN => n2026);
   U2191 : NAND2_X1 port map( A1 => n2245, A2 => n1735, ZN => n3669);
   U2192 : NOR2_X1 port map( A1 => n3640, A2 => n3641, ZN => n2027);
   U2193 : XNOR2_X1 port map( A => n1965, B => n536, ZN => n2144);
   U2194 : NAND2_X1 port map( A1 => n2028, A2 => Rst, ZN => n2097);
   U2195 : XNOR2_X1 port map( A => n2778, B => n2029, ZN => n2028);
   U2196 : INV_X1 port map( A => DataP_alu_b_in_7_port, ZN => n2030);
   U2197 : NAND2_X1 port map( A1 => n3423, A2 => n1748, ZN => n2031);
   U2198 : AOI21_X1 port map( B1 => n2037, B2 => n2032, A => n2671, ZN => n2670
                           );
   U2199 : NAND2_X1 port map( A1 => n2036, A2 => n2035, ZN => n2034);
   U2200 : INV_X1 port map( A => n2293, ZN => n2035);
   U2201 : NAND2_X1 port map( A1 => n2291, A2 => n2292, ZN => n2036);
   U2202 : NAND2_X1 port map( A1 => n2038, A2 => n2395, ZN => n2037);
   U2203 : OAI21_X1 port map( B1 => n3571, B2 => DataP_ALU_C_comp_N24, A => 
                           ALU_OPCODE_i_1_port, ZN => n2038);
   U2204 : OAI211_X1 port map( C1 => n2681, C2 => n3886, A => n2680, B => n3857
                           , ZN => n3609);
   U2205 : NAND2_X1 port map( A1 => n2681, A2 => n2680, ZN => n2040);
   U2206 : NAND2_X1 port map( A1 => n2042, A2 => n1647, ZN => n3618);
   U2207 : NAND2_X1 port map( A1 => n3421, A2 => n2113, ZN => n3604);
   U2208 : INV_X1 port map( A => n2371, ZN => n2145);
   U2209 : NAND2_X1 port map( A1 => n2581, A2 => n2052, ZN => n2045);
   U2210 : OAI211_X1 port map( C1 => n2581, C2 => n2053, A => n2049, B => n2045
                           , ZN => n2654);
   U2211 : OAI211_X1 port map( C1 => n2581, C2 => n2047, A => n2046, B => n2564
                           , ZN => n2055);
   U2212 : NAND3_X1 port map( A1 => n2048, A2 => n2581, A3 => n2049, ZN => 
                           n2046);
   U2213 : NAND2_X1 port map( A1 => n2049, A2 => n2053, ZN => n2047);
   U2214 : OAI21_X1 port map( B1 => n2051, B2 => n2236, A => n2050, ZN => n2049
                           );
   U2215 : NAND2_X1 port map( A1 => n2236, A2 => n2400, ZN => n2050);
   U2216 : NOR2_X1 port map( A1 => n2054, A2 => n2580, ZN => n2051);
   U2217 : NOR2_X1 port map( A1 => n1635, A2 => n2400, ZN => n2052);
   U2218 : OR2_X1 port map( A1 => n2236, A2 => n2054, ZN => n2053);
   U2219 : INV_X1 port map( A => n2400, ZN => n2054);
   U2220 : NAND2_X1 port map( A1 => n2055, A2 => n2562, ZN => DataP_PC_reg_N30)
                           ;
   U2221 : NAND4_X1 port map( A1 => n2060, A2 => n2058, A3 => n2057, A4 => 
                           n2056, ZN => DataP_PC_reg_N25);
   U2222 : NAND2_X1 port map( A1 => n1613, A2 => n1971, ZN => n2056);
   U2223 : NAND2_X1 port map( A1 => n3679, A2 => n2061, ZN => n2057);
   U2224 : INV_X1 port map( A => n2059, ZN => n2058);
   U2225 : OAI21_X1 port map( B1 => n2064, B2 => n2708, A => n1966, ZN => n2059
                           );
   U2226 : OR2_X1 port map( A1 => n3777, A2 => n1972, ZN => n2060);
   U2227 : INV_X1 port map( A => n4111, ZN => n2061);
   U2228 : NOR2_X1 port map( A1 => n3880, A2 => n4111, ZN => n2062);
   U2229 : NOR2_X1 port map( A1 => n2133, A2 => n1931, ZN => n2066);
   U2230 : NAND2_X1 port map( A1 => n2133, A2 => n1717, ZN => n2067);
   U2231 : NAND4_X1 port map( A1 => n3478, A2 => n3477, A3 => n3475, A4 => 
                           n3476, ZN => DataP_alu_b_in_12_port);
   U2232 : BUF_X1 port map( A => n3641, Z => n2068);
   U2233 : BUF_X1 port map( A => n538, Z => n2069);
   U2234 : OR2_X1 port map( A1 => n2071, A2 => n2746, ZN => n2070);
   U2235 : AOI21_X1 port map( B1 => n2766, B2 => n2432, A => n2765, ZN => n2071
                           );
   U2236 : AND2_X2 port map( A1 => n2634, A2 => n3292, ZN => n2072);
   U2237 : OR4_X2 port map( A1 => n2259, A2 => n2261, A3 => n2309, A4 => n1602,
                           ZN => n2268);
   U2238 : AND2_X2 port map( A1 => n2384, A2 => n2538, ZN => n2073);
   U2239 : AND4_X1 port map( A1 => n3322, A2 => n3321, A3 => n3319, A4 => n3320
                           , ZN => n2074);
   U2240 : AND2_X1 port map( A1 => n1755, A2 => n2093, ZN => n2076);
   U2241 : AND2_X1 port map( A1 => n1755, A2 => n2093, ZN => n3642);
   U2242 : OR2_X2 port map( A1 => n3399, A2 => n2690, ZN => 
                           DataP_alu_a_in_11_port);
   U2243 : AOI22_X1 port map( A1 => n3221, A2 => DataP_B_s_0_port, B1 => n3222,
                           B2 => DataP_IMM_s_0_port, ZN => n2077);
   U2244 : BUF_X1 port map( A => n2783, Z => n2078);
   U2245 : BUF_X1 port map( A => DataP_opcode_M_1_port, Z => n2079);
   U2246 : OR2_X1 port map( A1 => n2100, A2 => n2296, ZN => n2080);
   U2247 : OR2_X1 port map( A1 => DataP_alu_b_in_2_port, A2 => n1719, ZN => 
                           n2081);
   U2248 : INV_X1 port map( A => n3697, ZN => DataP_alu_a_in_27_port);
   U2249 : BUF_X1 port map( A => n3487, Z => n2084);
   U2250 : AND4_X1 port map( A1 => n2176, A2 => n2178, A3 => n2621, A4 => n2175
                           , ZN => n2085);
   U2251 : NOR2_X1 port map( A1 => n3271, A2 => n1970, ZN => n3272);
   U2252 : CLKBUF_X3 port map( A => n3402, Z => n3217);
   U2253 : BUF_X1 port map( A => n2282, Z => n2086);
   U2254 : NAND4_X1 port map( A1 => n2143, A2 => n1962, A3 => n2144, A4 => 
                           n3240, ZN => n2087);
   U2255 : AND2_X1 port map( A1 => n2620, A2 => n2398, ZN => n2088);
   U2256 : NOR2_X1 port map( A1 => n2637, A2 => n2087, ZN => n2089);
   U2257 : NAND4_X1 port map( A1 => n3307, A2 => n3306, A3 => n3305, A4 => 
                           n3304, ZN => n2090);
   U2258 : AND3_X1 port map( A1 => n3239, A2 => DataP_opcode_W_3_port, A3 => 
                           n2625, ZN => n2091);
   U2259 : OAI221_X1 port map( B1 => n2100, B2 => n2296, C1 => 
                           DataP_alu_b_in_2_port, C2 => n1719, A => n2313, ZN 
                           => n2314);
   U2260 : NOR2_X1 port map( A1 => DataP_alu_b_in_13_port, A2 => 
                           DataP_alu_b_in_12_port, ZN => n3639);
   U2261 : NOR2_X1 port map( A1 => n2098, A2 => n2659, ZN => n2094);
   U2262 : BUF_X1 port map( A => n3860, Z => n2095);
   U2263 : AND4_X2 port map( A1 => n3515, A2 => n3514, A3 => n3513, A4 => n3512
                           , ZN => n2230);
   U2264 : INV_X1 port map( A => DataP_alu_b_in_1_port, ZN => n3200);
   U2265 : BUF_X4 port map( A => n3200, Z => n3047);
   U2266 : INV_X1 port map( A => n2781, ZN => n2782);
   U2267 : BUF_X2 port map( A => DataP_alu_b_in_2_port, Z => n3203);
   U2268 : AND2_X1 port map( A1 => n2190, A2 => DataP_alu_a_in_26_port, ZN => 
                           n2096);
   U2269 : NAND4_X1 port map( A1 => n3307, A2 => n3306, A3 => n3305, A4 => 
                           n3304, ZN => n2098);
   U2270 : NAND2_X1 port map( A1 => n3717, A2 => n3797, ZN => n2484);
   U2271 : BUF_X1 port map( A => n2219, Z => n2155);
   U2272 : INV_X1 port map( A => DataP_alu_a_in_9_port, ZN => n2099);
   U2273 : INV_X1 port map( A => n2101, ZN => n2112);
   U2274 : INV_X1 port map( A => n3054, ZN => n2115);
   U2275 : INV_X1 port map( A => n3203, ZN => n3053);
   U2276 : OR2_X1 port map( A1 => n3380, A2 => n3379, ZN => 
                           DataP_alu_a_in_20_port);
   U2277 : INV_X1 port map( A => n2226, ZN => n2118);
   U2278 : INV_X1 port map( A => n2119, ZN => n2100);
   U2279 : BUF_X4 port map( A => n3054, Z => n2101);
   U2280 : INV_X2 port map( A => n2226, ZN => n3199);
   U2281 : BUF_X2 port map( A => n4190, Z => n2104);
   U2282 : BUF_X2 port map( A => n2126, Z => n2105);
   U2283 : INV_X1 port map( A => n2372, ZN => DataP_alu_b_in_7_port);
   U2284 : INV_X1 port map( A => n2141, ZN => n2106);
   U2285 : INV_X1 port map( A => DataP_alu_b_in_24_port, ZN => n2107);
   U2286 : AND2_X1 port map( A1 => n2389, A2 => n2133, ZN => n2193);
   U2287 : INV_X1 port map( A => DataP_alu_a_in_13_port, ZN => n2109);
   U2288 : INV_X1 port map( A => DataP_alu_a_in_8_port, ZN => n2110);
   U2289 : INV_X1 port map( A => DataP_alu_a_in_21_port, ZN => n2111);
   U2290 : INV_X1 port map( A => DataP_alu_a_in_5_port, ZN => n2113);
   U2291 : INV_X1 port map( A => DataP_alu_a_in_20_port, ZN => n2114);
   U2292 : NAND2_X1 port map( A1 => n2139, A2 => n1969, ZN => n2150);
   U2293 : INV_X1 port map( A => DataP_alu_a_in_11_port, ZN => n2116);
   U2294 : OR2_X1 port map( A1 => n3908, A2 => DataP_wrong_br, ZN => n4190);
   U2295 : BUF_X2 port map( A => n3046, Z => n2117);
   U2296 : INV_X1 port map( A => DataP_alu_b_in_3_port, ZN => n2119);
   U2297 : INV_X1 port map( A => DataP_alu_b_in_28_port, ZN => n2120);
   U2298 : NAND2_X1 port map( A1 => DataP_alu_b_in_22_port, A2 => n3886, ZN => 
                           n2402);
   U2299 : BUF_X1 port map( A => DataP_alu_b_in_21_port, Z => n2152);
   U2300 : NAND4_X1 port map( A1 => n3263, A2 => n3262, A3 => n3261, A4 => 
                           n3260, ZN => DataP_alu_b_in_9_port);
   U2301 : NAND4_X1 port map( A1 => n3442, A2 => n3441, A3 => n3439, A4 => 
                           n3440, ZN => DataP_alu_b_in_10_port);
   U2302 : INV_X1 port map( A => DataP_alu_b_in_31_port, ZN => n2121);
   U2303 : INV_X1 port map( A => DataP_alu_b_in_22_port, ZN => n2122);
   U2304 : INV_X1 port map( A => DataP_alu_b_in_18_port, ZN => n2123);
   U2305 : INV_X1 port map( A => DataP_alu_b_in_23_port, ZN => n2124);
   U2306 : INV_X1 port map( A => n3212, ZN => n3211);
   U2307 : INV_X1 port map( A => DataP_alu_b_in_29_port, ZN => n2125);
   U2308 : INV_X1 port map( A => n1601, ZN => n2126);
   U2309 : INV_X1 port map( A => DataP_alu_b_in_26_port, ZN => n2127);
   U2310 : INV_X1 port map( A => n3897, ZN => n2130);
   U2311 : INV_X1 port map( A => n4111, ZN => n2131);
   U2312 : NOR2_X1 port map( A1 => n3246, A2 => n2628, ZN => n2627);
   U2313 : AND4_X1 port map( A1 => n3474, A2 => n3473, A3 => n3472, A4 => n3471
                           , ZN => n2386);
   U2314 : INV_X2 port map( A => n3233, ZN => n2132);
   U2315 : AND2_X1 port map( A1 => n3884, A2 => n2489, ZN => n2755);
   U2316 : AND2_X1 port map( A1 => n2764, A2 => n2760, ZN => n2759);
   U2317 : INV_X1 port map( A => n2758, ZN => n3635);
   U2318 : AND3_X1 port map( A1 => n2168, A2 => n2155, A3 => n2167, ZN => n2763
                           );
   U2319 : AND2_X1 port map( A1 => n3728, A2 => n2365, ZN => n3826);
   U2320 : NAND2_X1 port map( A1 => n2586, A2 => n2186, ZN => n3797);
   U2321 : INV_X1 port map( A => n3713, ZN => n2133);
   U2322 : NOR2_X1 port map( A1 => DataP_alu_a_in_25_port, A2 => n2187, ZN => 
                           n2186);
   U2323 : INV_X1 port map( A => n4190, ZN => n3231);
   U2324 : INV_X1 port map( A => n4190, ZN => n3230);
   U2325 : AND2_X1 port map( A1 => DataP_alu_a_in_9_port, A2 => n3429, ZN => 
                           n2259);
   U2326 : BUF_X1 port map( A => DataP_alu_a_in_9_port, Z => n2207);
   U2327 : AND2_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => n2198, ZN => 
                           n2197);
   U2328 : INV_X1 port map( A => n2182, ZN => n2181);
   U2329 : INV_X1 port map( A => DataP_alu_a_in_12_port, ZN => n2134);
   U2330 : OAI21_X1 port map( B1 => n2703, B2 => n2185, A => n2108, ZN => n2182
                           );
   U2331 : INV_X1 port map( A => n2101, ZN => n3205);
   U2332 : AND2_X1 port map( A1 => n2703, A2 => n2185, ZN => n2184);
   U2333 : BUF_X1 port map( A => DataP_alu_a_in_11_port, Z => n2200);
   U2334 : OR2_X1 port map( A1 => n3368, A2 => n3367, ZN => 
                           DataP_alu_a_in_24_port);
   U2335 : OR2_X1 port map( A1 => n3362, A2 => n3361, ZN => 
                           DataP_alu_a_in_26_port);
   U2336 : INV_X1 port map( A => DataP_alu_a_in_18_port, ZN => n2135);
   U2337 : OR2_X1 port map( A1 => n3359, A2 => n3358, ZN => 
                           DataP_alu_a_in_28_port);
   U2338 : INV_X1 port map( A => DataP_alu_a_in_23_port, ZN => n2136);
   U2339 : OR2_X2 port map( A1 => n3382, A2 => n3381, ZN => 
                           DataP_alu_a_in_19_port);
   U2340 : INV_X1 port map( A => DataP_alu_a_in_25_port, ZN => n2137);
   U2341 : INV_X1 port map( A => DataP_alu_b_in_3_port, ZN => n3054);
   U2342 : INV_X1 port map( A => n2226, ZN => n2916);
   U2343 : INV_X1 port map( A => n2585, ZN => n2187);
   U2344 : INV_X1 port map( A => n3212, ZN => n2209);
   U2345 : INV_X1 port map( A => n2230, ZN => DataP_alu_b_in_15_port);
   U2346 : BUF_X1 port map( A => n1591, Z => n2166);
   U2347 : INV_X1 port map( A => n3214, ZN => n2139);
   U2348 : INV_X1 port map( A => DataP_alu_b_in_6_port, ZN => n2140);
   U2349 : BUF_X2 port map( A => n1550, Z => n2141);
   U2350 : INV_X1 port map( A => n2782, ZN => n2772);
   U2351 : AND3_X1 port map( A1 => n3549, A2 => n3259, A3 => n399, ZN => n3547)
                           ;
   U2352 : OAI21_X1 port map( B1 => n4148, B2 => n4147, A => Rst, ZN => n4149);
   U2353 : OR2_X1 port map( A1 => n4153, A2 => CU_I_cw_7_port, ZN => n4147);
   U2354 : NOR2_X1 port map( A1 => n4052, A2 => n4051, ZN => CU_I_cw_7_port);
   U2355 : AND2_X1 port map( A1 => n2237, A2 => n2639, ZN => n2398);
   U2356 : NAND2_X2 port map( A1 => n3438, A2 => Rst, ZN => n4110);
   U2357 : OR2_X2 port map( A1 => n3229, A2 => n4143, ZN => n4146);
   U2358 : NAND2_X1 port map( A1 => n2626, A2 => n2627, ZN => n3291);
   U2359 : INV_X1 port map( A => n3883, ZN => n2626);
   U2360 : AND2_X2 port map( A1 => WB_MUX_SEL_i_1_port, A2 => n294, ZN => n4143
                           );
   U2361 : CLKBUF_X1 port map( A => DataP_add_D_3_port, Z => n2146);
   U2362 : INV_X4 port map( A => n2380, ZN => n3055);
   U2363 : NAND2_X2 port map( A1 => n3432, A2 => n3435, ZN => n3897);
   U2364 : NOR2_X1 port map( A1 => n2637, A2 => n2142, ZN => n2636);
   U2365 : NAND4_X1 port map( A1 => n2143, A2 => n1962, A3 => n2144, A4 => 
                           n3240, ZN => n2142);
   U2366 : AND2_X1 port map( A1 => n2174, A2 => n2636, ZN => n2620);
   U2367 : OAI211_X1 port map( C1 => n3213, C2 => n41, A => n2149, B => n2148, 
                           ZN => n3334);
   U2368 : NAND2_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_1_port, ZN => 
                           n2148);
   U2369 : NAND2_X1 port map( A1 => n3209, A2 => DataP_alu_out_W_1_port, ZN => 
                           n2149);
   U2370 : NOR2_X1 port map( A1 => n2090, A2 => n2659, ZN => n2658);
   U2371 : AND4_X2 port map( A1 => n3326, A2 => n3325, A3 => n3324, A4 => n3323
                           , ZN => n2242);
   U2372 : NAND2_X1 port map( A1 => n3396, A2 => n2150, ZN => n3398);
   U2373 : NAND4_X4 port map( A1 => n3535, A2 => n3534, A3 => n3533, A4 => 
                           n3532, ZN => DataP_alu_b_in_16_port);
   U2374 : AOI21_X1 port map( B1 => n3843, B2 => n3420, A => n3419, ZN => n3426
                           );
   U2375 : NAND2_X1 port map( A1 => n3845, A2 => n3844, ZN => n3843);
   U2376 : NAND2_X1 port map( A1 => n2154, A2 => n2153, ZN => n3412);
   U2377 : NAND2_X1 port map( A1 => n3054, A2 => n3886, ZN => n2153);
   U2378 : NAND2_X1 port map( A1 => n3411, A2 => n2108, ZN => n2154);
   U2379 : NAND2_X1 port map( A1 => n3869, A2 => n3630, ZN => n2666);
   U2380 : NAND2_X1 port map( A1 => n2642, A2 => n3629, ZN => n3869);
   U2381 : NAND2_X1 port map( A1 => n2158, A2 => n2157, ZN => n3646);
   U2382 : NAND2_X1 port map( A1 => n2370, A2 => n3886, ZN => n2157);
   U2383 : NAND2_X1 port map( A1 => n3644, A2 => n2108, ZN => n2158);
   U2384 : NOR2_X1 port map( A1 => n2159, A2 => n2488, ZN => n2557);
   U2385 : NAND2_X1 port map( A1 => n2161, A2 => n2160, ZN => n2159);
   U2386 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N49, A2 => n3228, ZN =>
                           n2160);
   U2387 : INV_X1 port map( A => n3903, ZN => n2161);
   U2388 : OAI21_X1 port map( B1 => n2533, B2 => n2531, A => n2162, ZN => n2602
                           );
   U2389 : NAND2_X1 port map( A1 => n3763, A2 => n1746, ZN => n2162);
   U2390 : NAND2_X1 port map( A1 => n1738, A2 => n3691, ZN => n2213);
   U2391 : NAND2_X1 port map( A1 => n2074, A2 => n3886, ZN => n2163);
   U2392 : BUF_X1 port map( A => n1752, Z => n2164);
   U2393 : CLKBUF_X1 port map( A => n1566, Z => n2168);
   U2394 : OAI211_X1 port map( C1 => n3662, C2 => n3682, A => n1566, B => n2169
                           , ZN => n3687);
   U2395 : NAND2_X1 port map( A1 => n2549, A2 => n2547, ZN => n2169);
   U2396 : NAND2_X1 port map( A1 => n2546, A2 => n2108, ZN => n2549);
   U2397 : XNOR2_X1 port map( A => n3647, B => n1736, ZN => n2546);
   U2398 : NOR2_X1 port map( A1 => n3694, A2 => n3659, ZN => n3647);
   U2399 : NAND2_X1 port map( A1 => n3643, A2 => n2721, ZN => n2173);
   U2400 : OAI211_X1 port map( C1 => DataP_alu_b_in_17_port, C2 => n1738, A => 
                           n2170, B => n2172, ZN => n3643);
   U2401 : NAND2_X1 port map( A1 => n2245, A2 => n2171, ZN => n2170);
   U2402 : AND2_X1 port map( A1 => DataP_alu_b_in_17_port, A2 => n2370, ZN => 
                           n2171);
   U2403 : NAND2_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n1753, ZN => 
                           n2172);
   U2404 : NAND2_X1 port map( A1 => n2173, A2 => n2528, ZN => n3661);
   U2405 : AND2_X1 port map( A1 => n3289, A2 => n2638, ZN => n2174);
   U2406 : NAND3_X1 port map( A1 => n2174, A2 => n2089, A3 => n2639, ZN => 
                           n3258);
   U2407 : NOR2_X1 port map( A1 => n2097, A2 => n2406, ZN => n2175);
   U2408 : NAND2_X1 port map( A1 => n3250, A2 => n3251, ZN => n2176);
   U2409 : NAND2_X1 port map( A1 => n2177, A2 => n3248, ZN => n3251);
   U2410 : INV_X1 port map( A => n2179, ZN => n2177);
   U2411 : NOR2_X1 port map( A1 => n3883, A2 => n3246, ZN => n2178);
   U2412 : NAND4_X1 port map( A1 => n520, A2 => n17, A3 => n19, A4 => n21, ZN 
                           => n3883);
   U2413 : NAND2_X1 port map( A1 => n521, A2 => n23, ZN => n3246);
   U2414 : OAI211_X1 port map( C1 => n22, C2 => n2079, A => n2180, B => n2387, 
                           ZN => n2179);
   U2415 : NAND2_X1 port map( A1 => DataP_opcode_M_1_port, A2 => 
                           DataP_opcode_M_3_port, ZN => n2180);
   U2416 : NAND2_X1 port map( A1 => n3709, A2 => n2184, ZN => n2183);
   U2417 : OAI211_X1 port map( C1 => n2185, C2 => n1574, A => n2183, B => n2181
                           , ZN => n2189);
   U2418 : INV_X1 port map( A => DataP_alu_b_in_27_port, ZN => n2185);
   U2419 : XNOR2_X1 port map( A => n3720, B => n3697, ZN => n2188);
   U2420 : NAND2_X1 port map( A1 => n2189, A2 => n2540, ZN => n3720);
   U2421 : NAND3_X1 port map( A1 => n2192, A2 => n3690, A3 => n2193, ZN => 
                           n2191);
   U2422 : NAND2_X1 port map( A1 => n1633, A2 => n1717, ZN => n2192);
   U2423 : AND4_X2 port map( A1 => n3303, A2 => n3302, A3 => n3301, A4 => n3300
                           , ZN => n2372);
   U2424 : NAND4_X1 port map( A1 => n3307, A2 => n1583, A3 => n3305, A4 => 
                           n3304, ZN => DataP_alu_b_in_1_port);
   U2425 : OAI211_X1 port map( C1 => DataP_opcode_M_4_port, C2 => 
                           DataP_opcode_M_0_port, A => DataP_opcode_M_1_port, B
                           => DataP_opcode_M_2_port, ZN => n2195);
   U2426 : NAND2_X1 port map( A1 => n2196, A2 => n2197, ZN => n3738);
   U2427 : NAND2_X1 port map( A1 => n3644, A2 => n2534, ZN => n2196);
   U2428 : XNOR2_X1 port map( A => n1760, B => DataP_alu_b_in_16_port, ZN => 
                           n3644);
   U2429 : NAND2_X1 port map( A1 => n2534, A2 => n2535, ZN => n2198);
   U2430 : NAND2_X1 port map( A1 => n3738, A2 => n3660, ZN => n2527);
   U2431 : OAI21_X1 port map( B1 => n3643, B2 => n2128, A => n2397, ZN => n3660
                           );
   U2432 : OAI21_X1 port map( B1 => n2673, B2 => n2234, A => n2674, ZN => n2199
                           );
   U2433 : INV_X1 port map( A => n3537, ZN => n2201);
   U2434 : NOR2_X1 port map( A1 => n3382, A2 => n3381, ZN => n2202);
   U2435 : BUF_X1 port map( A => n3855, Z => n2203);
   U2436 : BUF_X1 port map( A => n3836, Z => n2204);
   U2437 : AND2_X1 port map( A1 => n3443, A2 => n1749, ZN => n2205);
   U2438 : BUF_X2 port map( A => n3401, Z => n3215);
   U2439 : INV_X1 port map( A => n3617, ZN => n2208);
   U2440 : NOR2_X1 port map( A1 => n3389, A2 => n2693, ZN => n2210);
   U2441 : BUF_X1 port map( A => n3611, Z => n2211);
   U2442 : XNOR2_X1 port map( A => n3799, B => n2212, ZN => n3806);
   U2443 : OR2_X1 port map( A1 => n2744, A2 => n3798, ZN => n2212);
   U2444 : BUF_X1 port map( A => n3869, Z => n2214);
   U2445 : BUF_X1 port map( A => n3604, Z => n2215);
   U2446 : AND2_X1 port map( A1 => n2594, A2 => n2593, ZN => n2216);
   U2447 : AOI21_X1 port map( B1 => n2560, B2 => n2129, A => n3679, ZN => n2217
                           );
   U2448 : BUF_X1 port map( A => n1584, Z => n2218);
   U2449 : AND2_X1 port map( A1 => n2525, A2 => n2524, ZN => n2220);
   U2450 : OR2_X2 port map( A1 => n3330, A2 => n3329, ZN => 
                           DataP_alu_a_in_2_port);
   U2451 : BUF_X1 port map( A => n1749, Z => n2221);
   U2452 : AND2_X1 port map( A1 => n3485, A2 => n3484, ZN => n2222);
   U2453 : INV_X1 port map( A => n2234, ZN => n2223);
   U2454 : INV_X1 port map( A => n1746, ZN => n2224);
   U2455 : AND2_X1 port map( A1 => n2687, A2 => n2686, ZN => n2225);
   U2456 : BUF_X1 port map( A => n3221, Z => n2227);
   U2457 : BUF_X2 port map( A => DataP_alu_a_in_0_port, Z => n2231);
   U2458 : OR2_X2 port map( A1 => n3334, A2 => n3333, ZN => n2232);
   U2459 : NAND2_X1 port map( A1 => n2077, A2 => n1593, ZN => n2233);
   U2460 : NAND2_X1 port map( A1 => n2656, A2 => n2657, ZN => 
                           DataP_alu_b_in_0_port);
   U2461 : AND2_X1 port map( A1 => n3308, A2 => n3309, ZN => n2657);
   U2462 : AND3_X1 port map( A1 => n1634, A2 => n2611, A3 => n2609, ZN => n2234
                           );
   U2463 : NAND2_X1 port map( A1 => n3464, A2 => n3491, ZN => n2235);
   U2464 : AND2_X1 port map( A1 => n2583, A2 => n2582, ZN => n2236);
   U2465 : AND2_X1 port map( A1 => n2627, A2 => n2626, ZN => n2237);
   U2466 : AND3_X2 port map( A1 => n3549, A2 => n3259, A3 => n2481, ZN => n3548
                           );
   U2467 : INV_X1 port map( A => n2762, ZN => n2238);
   U2468 : BUF_X1 port map( A => n3738, Z => n2239);
   U2469 : BUF_X2 port map( A => n3402, Z => n3218);
   U2470 : OAI21_X1 port map( B1 => n2096, B2 => n3719, A => n2188, ZN => n2241
                           );
   U2471 : AOI21_X1 port map( B1 => n1733, B2 => n2491, A => n2668, ZN => n2243
                           );
   U2472 : OAI221_X1 port map( B1 => n2293, B2 => n2292, C1 => n2291, C2 => 
                           n2293, A => n2290, ZN => DataP_ALU_C_comp_N24);
   U2473 : NOR2_X1 port map( A1 => n1760, A2 => n3659, ZN => n2244);
   U2474 : BUF_X2 port map( A => n3548, Z => n2246);
   U2475 : BUF_X2 port map( A => n3548, Z => n2247);
   U2476 : AOI21_X1 port map( B1 => n3251, B2 => n3250, A => n2406, ZN => n2248
                           );
   U2477 : NAND4_X1 port map( A1 => n3307, A2 => n1583, A3 => n3305, A4 => 
                           n3304, ZN => n2250);
   U2478 : NOR2_X1 port map( A1 => DataP_alu_b_in_29_port, A2 => n2295, ZN => 
                           n2252);
   U2479 : NAND2_X1 port map( A1 => DataP_alu_b_in_31_port, A2 => n2073, ZN => 
                           n2251);
   U2480 : OAI21_X1 port map( B1 => DataP_alu_b_in_30_port, B2 => n2294, A => 
                           n2251, ZN => n2280);
   U2481 : AOI211_X1 port map( C1 => DataP_alu_a_in_28_port, C2 => n2120, A => 
                           n2252, B => n2280, ZN => n2284);
   U2482 : AOI211_X1 port map( C1 => DataP_alu_a_in_24_port, C2 => n2107, A => 
                           n2086, B => n2297, ZN => n2253);
   U2483 : NAND2_X1 port map( A1 => n2284, A2 => n2253, ZN => n2293);
   U2484 : AOI21_X1 port map( B1 => DataP_alu_a_in_14_port, B2 => n2371, A => 
                           n2307, ZN => n2267);
   U2485 : OAI211_X1 port map( C1 => lt_x_135_B_12_port, C2 => n2134, A => 
                           n2308, B => n2267, ZN => n2261);
   U2486 : AOI21_X1 port map( B1 => DataP_alu_a_in_6_port, B2 => n2140, A => 
                           n2311, ZN => n2257);
   U2487 : OAI22_X1 port map( A1 => n2231, A2 => n2312, B1 => n2232, B2 => 
                           n2126, ZN => n2254);
   U2488 : OAI22_X1 port map( A1 => DataP_alu_a_in_6_port, A2 => n2318, B1 => 
                           DataP_alu_a_in_7_port, B2 => n2030, ZN => n2255);
   U2489 : OAI22_X1 port map( A1 => DataP_alu_a_in_12_port, A2 => n2321, B1 => 
                           DataP_alu_a_in_13_port, B2 => n2106, ZN => n2266);
   U2490 : NOR2_X1 port map( A1 => n2322, A2 => DataP_alu_a_in_10_port, ZN => 
                           n2258);
   U2491 : AOI22_X1 port map( A1 => n2165, A2 => n2258, B1 => n2151, B2 => 
                           n2116, ZN => n2263);
   U2492 : NOR2_X1 port map( A1 => DataP_alu_a_in_8_port, A2 => n2259, ZN => 
                           n2260);
   U2493 : AOI22_X1 port map( A1 => n2164, A2 => n2260, B1 => n2166, B2 => 
                           n2099, ZN => n2262);
   U2494 : AOI221_X1 port map( B1 => n1602, B2 => n2263, C1 => n2263, C2 => 
                           n2262, A => n2261, ZN => n2265);
   U2495 : NOR2_X1 port map( A1 => DataP_alu_b_in_17_port, A2 => n1750, ZN => 
                           n2272);
   U2496 : OAI211_X1 port map( C1 => DataP_alu_b_in_20_port, C2 => n2114, A => 
                           n2279, B => n2338, ZN => n2274);
   U2497 : AOI21_X1 port map( B1 => n2123, B2 => DataP_alu_a_in_18_port, A => 
                           n2341, ZN => n2269);
   U2498 : OAI21_X1 port map( B1 => n2152, B2 => n2111, A => 
                           DataP_alu_b_in_20_port, ZN => n2270);
   U2499 : OAI22_X1 port map( A1 => DataP_alu_a_in_20_port, A2 => n2270, B1 => 
                           DataP_alu_a_in_21_port, B2 => n3663, ZN => n2278);
   U2500 : NOR2_X1 port map( A1 => n2341, A2 => DataP_alu_a_in_18_port, ZN => 
                           n2271);
   U2501 : AOI22_X1 port map( A1 => n2271, A2 => n1736, B1 => n1722, B2 => 
                           n2202, ZN => n2276);
   U2502 : NOR2_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => n2272, ZN => 
                           n2273);
   U2503 : AOI22_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n2273, B1 => 
                           DataP_alu_b_in_17_port, B2 => n1750, ZN => n2275);
   U2504 : AOI221_X1 port map( B1 => n2298, B2 => n2276, C1 => n2275, C2 => 
                           n2276, A => n2274, ZN => n2277);
   U2505 : OAI21_X1 port map( B1 => DataP_alu_b_in_29_port, B2 => n2295, A => 
                           DataP_alu_b_in_28_port, ZN => n2281);
   U2506 : OAI22_X1 port map( A1 => DataP_alu_a_in_28_port, A2 => n2281, B1 => 
                           DataP_alu_a_in_29_port, B2 => n2125, ZN => n2289);
   U2507 : AOI22_X1 port map( A1 => DataP_alu_b_in_26_port, A2 => n2354, B1 => 
                           DataP_alu_b_in_27_port, B2 => n3697, ZN => n2285);
   U2508 : NOR2_X1 port map( A1 => DataP_alu_a_in_24_port, A2 => n2282, ZN => 
                           n2283);
   U2509 : AOI221_X1 port map( B1 => n2297, B2 => n2285, C1 => n2356, C2 => 
                           n2285, A => n2300, ZN => n2288);
   U2510 : OAI21_X1 port map( B1 => DataP_alu_a_in_31_port, B2 => n2121, A => 
                           DataP_alu_b_in_30_port, ZN => n2286);
   U2511 : OAI22_X1 port map( A1 => DataP_alu_a_in_30_port, A2 => n2286, B1 => 
                           DataP_alu_b_in_31_port, B2 => n2073, ZN => n2287);
   U2512 : AND2_X1 port map( A1 => DataP_alu_a_in_22_port, A2 => n2122, ZN => 
                           n2302);
   U2513 : INV_X1 port map( A => DataP_alu_a_in_29_port, ZN => n2295);
   U2514 : INV_X1 port map( A => DataP_alu_a_in_30_port, ZN => n2294);
   U2515 : INV_X1 port map( A => DataP_alu_a_in_3_port, ZN => n2296);
   U2516 : INV_X1 port map( A => DataP_alu_b_in_16_port, ZN => n2301);
   U2517 : AOI21_X1 port map( B1 => DataP_alu_a_in_23_port, B2 => n2124, A => 
                           n2302, ZN => n2279);
   U2518 : INV_X1 port map( A => n2269, ZN => n2298);
   U2519 : INV_X1 port map( A => n2280, ZN => n2299);
   U2520 : INV_X1 port map( A => n2284, ZN => n2300);
   U2521 : NOR2_X1 port map( A1 => DataP_alu_b_in_29_port, A2 => n2365, ZN => 
                           n2304);
   U2522 : NAND2_X1 port map( A1 => DataP_alu_a_in_31_port, A2 => n2121, ZN => 
                           n2303);
   U2523 : OAI21_X1 port map( B1 => DataP_alu_b_in_30_port, B2 => n2364, A => 
                           n2303, ZN => n2351);
   U2524 : AOI211_X1 port map( C1 => DataP_alu_a_in_28_port, C2 => n2120, A => 
                           n2304, B => n2351, ZN => n2355);
   U2525 : NOR2_X1 port map( A1 => n3697, A2 => DataP_alu_b_in_27_port, ZN => 
                           n2353);
   U2526 : AOI21_X1 port map( B1 => n2127, B2 => DataP_alu_a_in_26_port, A => 
                           n2353, ZN => n2305);
   U2527 : AOI211_X1 port map( C1 => DataP_alu_a_in_24_port, C2 => n2107, A => 
                           n2086, B => n2367, ZN => n2306);
   U2528 : NOR2_X1 port map( A1 => n2166, A2 => n2099, ZN => n2324);
   U2529 : NOR2_X1 port map( A1 => DataP_alu_b_in_15_port, A2 => n2210, ZN => 
                           n2307);
   U2530 : AOI21_X1 port map( B1 => DataP_alu_a_in_14_port, B2 => n2371, A => 
                           n2307, ZN => n2333);
   U2531 : NAND2_X1 port map( A1 => DataP_alu_a_in_13_port, A2 => n2106, ZN => 
                           n2308);
   U2532 : OAI211_X1 port map( C1 => lt_x_135_B_12_port, C2 => n2134, A => 
                           n2333, B => n2308, ZN => n2326);
   U2533 : NOR2_X1 port map( A1 => n2164, A2 => n2110, ZN => n2309);
   U2534 : NOR2_X1 port map( A1 => n2151, A2 => n2116, ZN => n2322);
   U2535 : OR4_X1 port map( A1 => n2324, A2 => n2326, A3 => n2309, A4 => n1602,
                           ZN => n2336);
   U2536 : OAI21_X1 port map( B1 => lt_x_135_B_5_port, B2 => n2113, A => n2138,
                           ZN => n2310);
   U2537 : OAI22_X1 port map( A1 => DataP_alu_a_in_4_port, A2 => n2310, B1 => 
                           DataP_alu_a_in_5_port, B2 => n2074, ZN => n2320);
   U2538 : NOR2_X1 port map( A1 => n2366, A2 => DataP_alu_b_in_7_port, ZN => 
                           n2311);
   U2539 : OAI21_X1 port map( B1 => n2100, B2 => n2296, A => 
                           DataP_alu_b_in_2_port, ZN => n2315);
   U2540 : OAI21_X1 port map( B1 => n2373, B2 => n2206, A => n2226, ZN => n2312
                           );
   U2541 : OAI22_X1 port map( A1 => n2231, A2 => n2312, B1 => n2232, B2 => 
                           n2126, ZN => n2313);
   U2542 : OAI221_X1 port map( B1 => n1973, B2 => n2119, C1 => 
                           DataP_alu_a_in_2_port, C2 => n2315, A => n2314, ZN 
                           => n2316);
   U2543 : OAI21_X1 port map( B1 => lt_x_135_B_5_port, B2 => n2113, A => n2316,
                           ZN => n2317);
   U2544 : AOI21_X1 port map( B1 => DataP_alu_a_in_4_port, B2 => n3206, A => 
                           n2317, ZN => n2319);
   U2545 : OAI21_X1 port map( B1 => n2366, B2 => DataP_alu_b_in_7_port, A => 
                           DataP_alu_b_in_6_port, ZN => n2318);
   U2546 : AOI221_X1 port map( B1 => n2320, B2 => n2257, C1 => n2319, C2 => 
                           n2257, A => n2255, ZN => n2335);
   U2547 : OAI21_X1 port map( B1 => n2141, B2 => n2109, A => lt_x_135_B_12_port
                           , ZN => n2321);
   U2548 : OAI22_X1 port map( A1 => DataP_alu_a_in_12_port, A2 => n2321, B1 => 
                           DataP_alu_a_in_13_port, B2 => n2106, ZN => n2332);
   U2549 : NOR2_X1 port map( A1 => DataP_alu_a_in_10_port, A2 => n2322, ZN => 
                           n2323);
   U2550 : AOI22_X1 port map( A1 => n2165, A2 => n2323, B1 => n2151, B2 => 
                           n2116, ZN => n2328);
   U2551 : NOR2_X1 port map( A1 => DataP_alu_a_in_8_port, A2 => n2324, ZN => 
                           n2325);
   U2552 : AOI22_X1 port map( A1 => n2164, A2 => n2325, B1 => n2166, B2 => 
                           n2099, ZN => n2327);
   U2553 : AOI221_X1 port map( B1 => n1602, B2 => n2328, C1 => n2327, C2 => 
                           n2328, A => n2326, ZN => n2331);
   U2554 : OAI22_X1 port map( A1 => DataP_alu_a_in_14_port, A2 => n2329, B1 => 
                           DataP_alu_a_in_15_port, B2 => n2230, ZN => n2330);
   U2555 : AOI211_X1 port map( C1 => n2333, C2 => n2332, A => n2331, B => n2330
                           , ZN => n2334);
   U2556 : OAI21_X1 port map( B1 => n2336, B2 => n2335, A => n2334, ZN => n2340
                           );
   U2557 : NOR2_X1 port map( A1 => DataP_alu_b_in_17_port, A2 => n1750, ZN => 
                           n2342);
   U2558 : NOR2_X1 port map( A1 => DataP_alu_b_in_23_port, A2 => n2136, ZN => 
                           n2337);
   U2559 : AOI21_X1 port map( B1 => DataP_alu_a_in_22_port, B2 => n2122, A => 
                           n2337, ZN => n2350);
   U2560 : NAND2_X1 port map( A1 => DataP_alu_a_in_21_port, A2 => n3663, ZN => 
                           n2338);
   U2561 : OAI211_X1 port map( C1 => DataP_alu_b_in_20_port, C2 => n2114, A => 
                           n2350, B => n2338, ZN => n2344);
   U2562 : NOR2_X1 port map( A1 => n1722, A2 => n2202, ZN => n2341);
   U2563 : AOI211_X1 port map( C1 => DataP_alu_a_in_16_port, C2 => n2370, A => 
                           n2344, B => n2298, ZN => n2339);
   U2564 : NAND3_X1 port map( A1 => n2340, A2 => n2369, A3 => n2339, ZN => 
                           n2363);
   U2565 : NOR2_X1 port map( A1 => DataP_alu_a_in_16_port, A2 => n2342, ZN => 
                           n2343);
   U2566 : AOI22_X1 port map( A1 => DataP_alu_b_in_16_port, A2 => n2343, B1 => 
                           DataP_alu_b_in_17_port, B2 => n1750, ZN => n2345);
   U2567 : AOI221_X1 port map( B1 => n2298, B2 => n2346, C1 => n2345, C2 => 
                           n2346, A => n2344, ZN => n2349);
   U2568 : OAI21_X1 port map( B1 => DataP_alu_b_in_23_port, B2 => n2136, A => 
                           DataP_alu_b_in_22_port, ZN => n2347);
   U2569 : OAI22_X1 port map( A1 => DataP_alu_a_in_22_port, A2 => n2347, B1 => 
                           DataP_alu_a_in_23_port, B2 => n2124, ZN => n2348);
   U2570 : AOI211_X1 port map( C1 => n2350, C2 => n2278, A => n2349, B => n2348
                           , ZN => n2362);
   U2571 : OAI21_X1 port map( B1 => DataP_alu_b_in_29_port, B2 => n2365, A => 
                           DataP_alu_b_in_28_port, ZN => n2352);
   U2572 : OAI22_X1 port map( A1 => DataP_alu_a_in_28_port, A2 => n2352, B1 => 
                           DataP_alu_a_in_29_port, B2 => n2125, ZN => n2360);
   U2573 : NOR2_X1 port map( A1 => DataP_alu_a_in_26_port, A2 => n2353, ZN => 
                           n2354);
   U2574 : OAI21_X1 port map( B1 => DataP_alu_b_in_31_port, B2 => n2073, A => 
                           DataP_alu_b_in_30_port, ZN => n2357);
   U2575 : OAI22_X1 port map( A1 => DataP_alu_a_in_30_port, A2 => n2357, B1 => 
                           DataP_alu_a_in_31_port, B2 => n2121, ZN => n2358);
   U2576 : AOI211_X1 port map( C1 => n2368, C2 => n2360, A => n2359, B => n2358
                           , ZN => n2361);
   U2577 : INV_X1 port map( A => n2126, ZN => n2373);
   U2578 : INV_X1 port map( A => DataP_alu_a_in_29_port, ZN => n2365);
   U2579 : INV_X1 port map( A => DataP_alu_a_in_30_port, ZN => n2364);
   U2580 : INV_X1 port map( A => n2305, ZN => n2367);
   U2581 : INV_X1 port map( A => DataP_alu_a_in_7_port, ZN => n2366);
   U2582 : INV_X1 port map( A => n2342, ZN => n2369);
   U2583 : INV_X1 port map( A => DataP_alu_b_in_16_port, ZN => n2370);
   U2584 : INV_X1 port map( A => n2351, ZN => n2368);
   U2585 : NAND2_X1 port map( A1 => n2620, A2 => n2398, ZN => n3259);
   U2586 : INV_X1 port map( A => DataP_alu_b_in_20_port, ZN => n3664);
   U2587 : INV_X1 port map( A => DataP_alu_b_in_21_port, ZN => n3663);
   U2588 : BUF_X2 port map( A => n3547, Z => n3219);
   U2589 : NOR2_X1 port map( A1 => n516, A2 => n4044, ZN => n4049);
   U2590 : AND2_X1 port map( A1 => n2776, A2 => n2403, ZN => n2480);
   U2591 : INV_X1 port map( A => n4055, ZN => n4036);
   U2592 : NOR2_X1 port map( A1 => IR_CU_27, A2 => IR_CU_26, ZN => n4055);
   U2593 : INV_X1 port map( A => n3131, ZN => n3195);
   U2594 : AND3_X1 port map( A1 => DataP_opcode_W_2_port, A2 => 
                           DataP_opcode_W_4_port, A3 => n2401, ZN => n2483);
   U2595 : INV_X1 port map( A => n4188, ZN => n491);
   U2596 : INV_X1 port map( A => n4187, ZN => n492);
   U2597 : INV_X1 port map( A => n4156, ZN => n4148);
   U2598 : NAND2_X1 port map( A1 => n516, A2 => n1960, ZN => n3994);
   U2599 : BUF_X1 port map( A => n3900, Z => n3227);
   U2600 : AND3_X1 port map( A1 => n3409, A2 => n3886, A3 => n3408, ZN => n3880
                           );
   U2601 : INV_X1 port map( A => n3892, ZN => n3877);
   U2602 : INV_X1 port map( A => n4186, ZN => n493);
   U2603 : INV_X1 port map( A => n4185, ZN => n494);
   U2604 : INV_X1 port map( A => n4189, ZN => n490);
   U2605 : NOR2_X1 port map( A1 => n486, A2 => n4149, ZN => DataP_add_S2_1_port
                           );
   U2606 : NOR2_X1 port map( A1 => n487, A2 => n4149, ZN => DataP_add_S2_2_port
                           );
   U2607 : NOR2_X1 port map( A1 => n488, A2 => n4149, ZN => DataP_add_S2_3_port
                           );
   U2608 : NOR2_X1 port map( A1 => n489, A2 => n4149, ZN => DataP_add_S2_4_port
                           );
   U2609 : NOR2_X1 port map( A1 => n485, A2 => n4149, ZN => DataP_add_S2_0_port
                           );
   U2610 : INV_X1 port map( A => n4151, ZN => n4052);
   U2611 : NOR3_X1 port map( A1 => n3994, A2 => n4155, A3 => n4036, ZN => n4153
                           );
   U2612 : NOR2_X1 port map( A1 => n3994, A2 => n2374, ZN => n16);
   U2613 : BUF_X1 port map( A => n3904, Z => n3228);
   U2614 : OR2_X1 port map( A1 => n2773, A2 => n2471, ZN => n3312);
   U2615 : AND4_X1 port map( A1 => n3249, A2 => n1638, A3 => n528, A4 => n1637,
                           ZN => n2406);
   U2616 : NOR2_X1 port map( A1 => n504, A2 => n497, ZN => n4166);
   U2617 : OR2_X1 port map( A1 => n4101, A2 => ALU_OPCODE_i_0_port, ZN => n4184
                           );
   U2618 : AND2_X2 port map( A1 => n3638, A2 => n3637, ZN => n3680);
   U2619 : AND2_X1 port map( A1 => BR_EN_i, A2 => n4102, ZN => n3908);
   U2620 : NOR2_X1 port map( A1 => ALU_OPCODE_i_3_port, A2 => 
                           ALU_OPCODE_i_0_port, ZN => n3561);
   U2621 : BUF_X1 port map( A => n4222, Z => n3232);
   U2622 : NOR2_X1 port map( A1 => n3231, A2 => n3235, ZN => n4222);
   U2623 : INV_X1 port map( A => Rst, ZN => n3236);
   U2624 : INV_X1 port map( A => Rst, ZN => n3235);
   U2625 : INV_X1 port map( A => DataP_npc_mux_sel, ZN => n3233);
   U2626 : BUF_X1 port map( A => n4144, Z => n3229);
   U2627 : NOR2_X1 port map( A1 => WB_MUX_SEL_i_1_port, A2 => n294, ZN => n4144
                           );
   U2628 : INV_X1 port map( A => n4165, ZN => n4181);
   U2629 : NAND2_X2 port map( A1 => n1586, A2 => n3310, ZN => 
                           DataP_alu_b_in_3_port);
   U2630 : OR2_X2 port map( A1 => n3392, A2 => n3391, ZN => 
                           DataP_alu_a_in_14_port);
   U2631 : INV_X2 port map( A => n3212, ZN => n3210);
   U2632 : BUF_X2 port map( A => n3547, Z => n3221);
   U2633 : NOR4_X1 port map( A1 => n443, A2 => ALU_OPCODE_i_3_port, A3 => 
                           ALU_OPCODE_i_2_port, A4 => ALU_OPCODE_i_1_port, ZN 
                           => n4102);
   U2634 : INV_X2 port map( A => n3891, ZN => n3894);
   U2635 : INV_X2 port map( A => DataP_alu_b_in_2_port, ZN => n3052);
   U2636 : OR2_X2 port map( A1 => n3371, A2 => n3370, ZN => 
                           DataP_alu_a_in_23_port);
   U2637 : OR2_X2 port map( A1 => n3374, A2 => n3373, ZN => 
                           DataP_alu_a_in_22_port);
   U2638 : OR2_X2 port map( A1 => n3388, A2 => n3387, ZN => 
                           DataP_alu_a_in_16_port);
   U2639 : OR2_X2 port map( A1 => n3299, A2 => n3298, ZN => 
                           DataP_alu_a_in_7_port);
   U2640 : OR2_X2 port map( A1 => n3337, A2 => n3336, ZN => 
                           DataP_alu_a_in_4_port);
   U2641 : OR2_X2 port map( A1 => n3346, A2 => n3345, ZN => 
                           DataP_alu_a_in_8_port);
   U2642 : OR2_X2 port map( A1 => n3395, A2 => n3394, ZN => 
                           DataP_alu_a_in_13_port);
   U2643 : OR2_X2 port map( A1 => n3389, A2 => n2693, ZN => 
                           DataP_alu_a_in_15_port);
   U2644 : BUF_X2 port map( A => n2088, Z => n3226);
   U2645 : OR2_X2 port map( A1 => n3353, A2 => n3352, ZN => 
                           DataP_alu_a_in_30_port);
   U2646 : BUF_X2 port map( A => n2088, Z => n3224);
   U2647 : BUF_X2 port map( A => n2088, Z => n3225);
   U2648 : BUF_X2 port map( A => n3547, Z => n3220);
   U2649 : INV_X2 port map( A => n2072, ZN => n3208);
   U2650 : AOI211_X1 port map( C1 => n4183, C2 => n3907, A => n4182, B => n3906
                           , ZN => DataP_right_br);
   U2651 : AND2_X1 port map( A1 => n4184, A2 => n1905, ZN => n3906);
   U2652 : NAND2_X1 port map( A1 => n3435, A2 => ALU_OPCODE_i_0_port, ZN => 
                           n3907);
   U2653 : INV_X1 port map( A => DataP_add_S2_3_port, ZN => n2767);
   U2654 : INV_X1 port map( A => DataP_add_S2_1_port, ZN => n2770);
   U2655 : AOI211_X1 port map( C1 => n3877, C2 => DataP_ALU_C_shifter_N83, A =>
                           n3584, B => n3583, ZN => n358);
   U2656 : AND2_X1 port map( A1 => DataP_ALU_C_shifter_N51, A2 => n3227, ZN => 
                           n3583);
   U2657 : OAI211_X1 port map( C1 => n3880, C2 => n3582, A => n3581, B => n3580
                           , ZN => n3584);
   U2658 : AOI21_X1 port map( B1 => n2130, B2 => n3579, A => n3578, ZN => n3580
                           );
   U2659 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N19, A2 => n3904, ZN =>
                           n3581);
   U2660 : INV_X1 port map( A => n2827, ZN => n2908);
   U2661 : NAND2_X1 port map( A1 => n1622, A2 => n1754, ZN => n3576);
   U2662 : AOI211_X1 port map( C1 => n3877, C2 => DataP_ALU_C_shifter_N84, A =>
                           n3596, B => n3595, ZN => n357);
   U2663 : OAI211_X1 port map( C1 => n3880, C2 => n3594, A => n3593, B => n3592
                           , ZN => n3595);
   U2664 : AOI21_X1 port map( B1 => n2130, B2 => n3591, A => n3590, ZN => n3592
                           );
   U2665 : OAI22_X1 port map( A1 => n1719, A2 => n3589, B1 => n3052, B2 => 
                           n3891, ZN => n3590);
   U2666 : AOI21_X1 port map( B1 => DataP_alu_b_in_2_port, B2 => n3890, A => 
                           n3894, ZN => n3589);
   U2667 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N20, A2 => n3228, ZN =>
                           n3593);
   U2668 : INV_X1 port map( A => n2884, ZN => n2909);
   U2669 : NAND2_X1 port map( A1 => n3586, A2 => n3585, ZN => n3587);
   U2670 : AND2_X1 port map( A1 => DataP_ALU_C_shifter_N52, A2 => n3227, ZN => 
                           n3596);
   U2671 : INV_X1 port map( A => DataP_add_S2_0_port, ZN => n2768);
   U2672 : INV_X1 port map( A => DataP_add_S2_4_port, ZN => n2769);
   U2673 : OAI22_X1 port map( A1 => n356, A2 => n4111, B1 => n4219, B2 => n4110
                           , ZN => DataP_PC_reg_N5);
   U2674 : AOI21_X1 port map( B1 => n2101, B2 => n3891, A => n3856, ZN => n3846
                           );
   U2675 : OAI211_X1 port map( C1 => n1644, C2 => n1662, A => n2218, B => n2129
                           , ZN => n3847);
   U2676 : INV_X1 port map( A => n2895, ZN => n2910);
   U2677 : INV_X1 port map( A => n2897, ZN => n2912);
   U2678 : OAI22_X1 port map( A1 => n355, A2 => n4111, B1 => n4218, B2 => n4110
                           , ZN => DataP_PC_reg_N6);
   U2679 : OAI21_X1 port map( B1 => n3851, B2 => n2102, A => n3891, ZN => n3852
                           );
   U2680 : INV_X1 port map( A => n2896, ZN => n2911);
   U2681 : OAI22_X1 port map( A1 => n353, A2 => n4111, B1 => n4216, B2 => n4110
                           , ZN => DataP_PC_reg_N8);
   U2682 : AOI211_X1 port map( C1 => n3857, C2 => n3891, A => n1748, B => n3856
                           , ZN => n3858);
   U2683 : OAI22_X1 port map( A1 => n345, A2 => n4111, B1 => n4214, B2 => n4110
                           , ZN => DataP_PC_reg_N10);
   U2684 : AOI21_X1 port map( B1 => n3841, B2 => n2130, A => n3894, ZN => n3840
                           );
   U2685 : INV_X1 port map( A => n3838, ZN => n3856);
   U2686 : NOR2_X1 port map( A1 => n2130, A2 => n3894, ZN => n3839);
   U2687 : INV_X1 port map( A => n2900, ZN => n2914);
   U2688 : AOI22_X1 port map( A1 => n3436, A2 => n2166, B1 => n3894, B2 => 
                           n2207, ZN => n3437);
   U2689 : OAI21_X1 port map( B1 => n2099, B2 => n3851, A => n3891, ZN => n3436
                           );
   U2690 : INV_X1 port map( A => n2901, ZN => n2915);
   U2691 : INV_X1 port map( A => n3835, ZN => n3428);
   U2692 : OAI21_X1 port map( B1 => n2366, B2 => n3851, A => n3891, ZN => n3612
                           );
   U2693 : INV_X1 port map( A => n2899, ZN => n2913);
   U2694 : INV_X1 port map( A => n1655, ZN => n3610);
   U2695 : AOI21_X1 port map( B1 => n3607, B2 => n2156, A => n3605, ZN => n3854
                           );
   U2696 : INV_X1 port map( A => n2215, ZN => n3605);
   U2697 : OAI21_X1 port map( B1 => n3850, B2 => n3600, A => n3599, ZN => n3607
                           );
   U2698 : INV_X1 port map( A => n3598, ZN => n3600);
   U2699 : NAND2_X1 port map( A1 => n2218, A2 => n3597, ZN => n3850);
   U2700 : AOI22_X1 port map( A1 => n3452, A2 => n2165, B1 => n3894, B2 => 
                           DataP_alu_a_in_10_port, ZN => n3453);
   U2701 : OAI21_X1 port map( B1 => n3451, B2 => n3851, A => n3891, ZN => n3452
                           );
   U2702 : INV_X1 port map( A => n2863, ZN => n2902);
   U2703 : INV_X1 port map( A => n3484, ZN => n3450);
   U2704 : INV_X1 port map( A => n2875, ZN => n2904);
   U2705 : NAND2_X1 port map( A1 => DataP_alu_a_in_12_port, A2 => n2655, ZN => 
                           n3492);
   U2706 : NOR2_X1 port map( A1 => n1573, A2 => n3851, ZN => n2655);
   U2707 : OAI21_X1 port map( B1 => DataP_alu_a_in_12_port, B2 => 
                           lt_x_135_B_12_port, A => n3894, ZN => n3493);
   U2708 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N29, A2 => n3228, ZN =>
                           n3471);
   U2709 : INV_X1 port map( A => n2868, ZN => n2903);
   U2710 : AOI21_X1 port map( B1 => n3540, B2 => n2130, A => n3470, ZN => n3472
                           );
   U2711 : OAI22_X1 port map( A1 => n3469, A2 => n3468, B1 => n3467, B2 => 
                           n3891, ZN => n3470);
   U2712 : AOI21_X1 port map( B1 => n2200, B2 => n3890, A => n3894, ZN => n3469
                           );
   U2713 : AOI22_X1 port map( A1 => n3227, A2 => DataP_ALU_C_shifter_N61, B1 =>
                           DataP_ALU_C_shifter_N93, B2 => n3877, ZN => n3473);
   U2714 : NAND2_X1 port map( A1 => n3466, A2 => n2129, ZN => n3474);
   U2715 : XNOR2_X1 port map( A => n3465, B => n3488, ZN => n3466);
   U2716 : OAI21_X1 port map( B1 => n3458, B2 => n3489, A => n3484, ZN => n3465
                           );
   U2717 : NAND2_X1 port map( A1 => n3446, A2 => n3445, ZN => n3458);
   U2718 : NAND2_X1 port map( A1 => n3444, A2 => n3443, ZN => n3445);
   U2719 : NAND2_X1 port map( A1 => n3483, A2 => n3835, ZN => n3444);
   U2720 : NAND2_X1 port map( A1 => n3837, A2 => n2205, ZN => n3446);
   U2721 : NAND2_X1 port map( A1 => n2084, A2 => n3482, ZN => n3837);
   U2722 : OAI22_X1 port map( A1 => n333, A2 => n4111, B1 => n4110, B2 => n4209
                           , ZN => DataP_PC_reg_N15);
   U2723 : INV_X1 port map( A => DataP_npc_13_port, ZN => n4209);
   U2724 : OAI21_X1 port map( B1 => DataP_alu_a_in_13_port, B2 => n2141, A => 
                           n3894, ZN => n3871);
   U2725 : INV_X1 port map( A => n2882, ZN => n2905);
   U2726 : NAND2_X1 port map( A1 => n1710, A2 => n3863, ZN => n3866);
   U2727 : OAI22_X1 port map( A1 => n326, A2 => n4111, B1 => n4110, B2 => n4206
                           , ZN => DataP_PC_reg_N18);
   U2728 : INV_X1 port map( A => DataP_npc_16_port, ZN => n4206);
   U2729 : AOI21_X1 port map( B1 => n3737, B2 => n2129, A => n3736, ZN => n326)
                           ;
   U2730 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N34, A2 => n3228, ZN =>
                           n3733);
   U2731 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N66, B2 => n3227, A => 
                           n3732, ZN => n3735);
   U2732 : OAI22_X1 port map( A1 => n319, A2 => n4111, B1 => n4110, B2 => n4203
                           , ZN => DataP_PC_reg_N21);
   U2733 : INV_X1 port map( A => DataP_npc_19_port, ZN => n4203);
   U2734 : AOI21_X1 port map( B1 => n3658, B2 => n2129, A => n3657, ZN => n319)
                           ;
   U2735 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N37, A2 => n3904, ZN =>
                           n3654);
   U2736 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N69, B2 => n3900, A => 
                           n3653, ZN => n3655);
   U2737 : OAI211_X1 port map( C1 => n4106, C2 => n3897, A => n3652, B => n3651
                           , ZN => n3653);
   U2738 : NAND2_X1 port map( A1 => DataP_alu_a_in_19_port, A2 => n3894, ZN => 
                           n3651);
   U2739 : OAI211_X1 port map( C1 => DataP_alu_a_in_19_port, C2 => n3894, A => 
                           n1722, B => n3838, ZN => n3652);
   U2740 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N101, A2 => n3877, ZN 
                           => n3656);
   U2741 : OAI22_X1 port map( A1 => n322, A2 => n4111, B1 => n4110, B2 => n4204
                           , ZN => DataP_PC_reg_N20);
   U2742 : INV_X1 port map( A => DataP_npc_18_port, ZN => n4204);
   U2743 : INV_X1 port map( A => n3752, ZN => n322);
   U2744 : OAI211_X1 port map( C1 => n3751, C2 => n3880, A => n3750, B => n3749
                           , ZN => n3752);
   U2745 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N100, A2 => n3877, ZN 
                           => n3749);
   U2746 : AOI21_X1 port map( B1 => n3904, B2 => DataP_ALU_C_shifter_N36, A => 
                           n3748, ZN => n3750);
   U2747 : NAND3_X1 port map( A1 => n2724, A2 => n3635, A3 => n2378, ZN => 
                           n2673);
   U2748 : OAI22_X1 port map( A1 => n323, A2 => n4111, B1 => n4110, B2 => n4205
                           , ZN => DataP_PC_reg_N19);
   U2749 : INV_X1 port map( A => DataP_npc_17_port, ZN => n4205);
   U2750 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N67, B2 => n3227, A => 
                           n3742, ZN => n3744);
   U2751 : OAI211_X1 port map( C1 => n3741, C2 => n3897, A => n3740, B => n3739
                           , ZN => n3742);
   U2752 : OAI211_X1 port map( C1 => n1751, C2 => n3894, A => 
                           DataP_alu_b_in_17_port, B => n3838, ZN => n3739);
   U2753 : NAND2_X1 port map( A1 => n1751, A2 => n3894, ZN => n3740);
   U2754 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N99, A2 => n3877, ZN =>
                           n3745);
   U2755 : NAND2_X1 port map( A1 => n2078, A2 => n3680, ZN => n3729);
   U2756 : OAI22_X1 port map( A1 => n311, A2 => n4111, B1 => n4110, B2 => n4200
                           , ZN => DataP_PC_reg_N24);
   U2757 : INV_X1 port map( A => DataP_npc_22_port, ZN => n4200);
   U2758 : AOI21_X1 port map( B1 => n3787, B2 => n2129, A => n3786, ZN => n311)
                           ;
   U2759 : OAI21_X1 port map( B1 => n3892, B2 => n3785, A => n3784, ZN => n3786
                           );
   U2760 : AOI21_X1 port map( B1 => n3904, B2 => DataP_ALU_C_shifter_N40, A => 
                           n3783, ZN => n3784);
   U2761 : OAI211_X1 port map( C1 => n3897, C2 => n3782, A => n3781, B => n3780
                           , ZN => n3783);
   U2762 : AOI22_X1 port map( A1 => n3779, A2 => DataP_alu_b_in_22_port, B1 => 
                           n3894, B2 => DataP_alu_a_in_22_port, ZN => n3780);
   U2763 : OAI21_X1 port map( B1 => n3778, B2 => n3851, A => n3891, ZN => n3779
                           );
   U2764 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N72, A2 => n3227, ZN =>
                           n3781);
   U2765 : INV_X1 port map( A => DataP_ALU_C_shifter_N104, ZN => n3785);
   U2766 : XNOR2_X1 port map( A => n3777, B => n3776, ZN => n3787);
   U2767 : INV_X1 port map( A => DataP_npc_21_port, ZN => n4201);
   U2768 : OAI21_X1 port map( B1 => n3892, B2 => n3774, A => n3773, ZN => n3775
                           );
   U2769 : AOI21_X1 port map( B1 => n3904, B2 => DataP_ALU_C_shifter_N39, A => 
                           n3772, ZN => n3773);
   U2770 : OAI211_X1 port map( C1 => n3897, C2 => n3771, A => n3770, B => n3769
                           , ZN => n3772);
   U2771 : AOI22_X1 port map( A1 => n3768, A2 => n2152, B1 => n3894, B2 => 
                           DataP_alu_a_in_21_port, ZN => n3769);
   U2772 : OAI21_X1 port map( B1 => n2111, B2 => n3851, A => n3891, ZN => n3768
                           );
   U2773 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N71, A2 => n3227, ZN =>
                           n3770);
   U2774 : INV_X1 port map( A => DataP_ALU_C_shifter_N103, ZN => n3774);
   U2775 : INV_X1 port map( A => n1588, ZN => n3765);
   U2776 : OAI22_X1 port map( A1 => n317, A2 => n4111, B1 => n4110, B2 => n4202
                           , ZN => DataP_PC_reg_N22);
   U2777 : INV_X1 port map( A => DataP_npc_20_port, ZN => n4202);
   U2778 : AOI21_X1 port map( B1 => n3761, B2 => n2129, A => n3760, ZN => n317)
                           ;
   U2779 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N38, A2 => n3228, ZN =>
                           n3757);
   U2780 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N70, B2 => n3227, A => 
                           n3756, ZN => n3758);
   U2781 : OAI211_X1 port map( C1 => n4107, C2 => n3897, A => n3755, B => n3754
                           , ZN => n3756);
   U2782 : NAND2_X1 port map( A1 => DataP_alu_a_in_20_port, A2 => n3894, ZN => 
                           n3754);
   U2783 : OAI211_X1 port map( C1 => DataP_alu_a_in_20_port, C2 => n3894, A => 
                           DataP_alu_b_in_20_port, B => n3838, ZN => n3755);
   U2784 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N102, A2 => n3877, ZN 
                           => n3759);
   U2785 : OAI22_X1 port map( A1 => n308, A2 => n4111, B1 => n4110, B2 => n4198
                           , ZN => DataP_PC_reg_N26);
   U2786 : INV_X1 port map( A => DataP_npc_24_port, ZN => n4198);
   U2787 : AOI21_X1 port map( B1 => n3796, B2 => n2129, A => n3795, ZN => n308)
                           ;
   U2788 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N42, A2 => n3228, ZN =>
                           n3792);
   U2789 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N74, B2 => n3227, A => 
                           n3791, ZN => n3793);
   U2790 : OAI211_X1 port map( C1 => n4109, C2 => n3897, A => n3790, B => n3789
                           , ZN => n3791);
   U2791 : NAND2_X1 port map( A1 => DataP_alu_a_in_24_port, A2 => n3894, ZN => 
                           n3789);
   U2792 : OAI211_X1 port map( C1 => DataP_alu_a_in_24_port, C2 => n3894, A => 
                           DataP_alu_b_in_24_port, B => n3838, ZN => n3790);
   U2793 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N106, A2 => n3877, ZN 
                           => n3794);
   U2794 : INV_X1 port map( A => n3127, ZN => n3197);
   U2795 : AND3_X1 port map( A1 => n2555, A2 => n2556, A3 => n2558, ZN => n297)
                           ;
   U2796 : OR2_X1 port map( A1 => n2752, A2 => n2083, ZN => n2555);
   U2797 : AOI21_X1 port map( B1 => n2654, B2 => n2129, A => n3824, ZN => n300)
                           ;
   U2798 : INV_X1 port map( A => DataP_npc_26_port, ZN => n4196);
   U2799 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N108, A2 => n3877, ZN 
                           => n3812);
   U2800 : INV_X1 port map( A => n3133, ZN => DataP_ALU_C_shifter_N108);
   U2801 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N76, B2 => n3227, A => 
                           n3811, ZN => n3813);
   U2802 : OAI211_X1 port map( C1 => n3810, C2 => n3897, A => n3809, B => n3808
                           , ZN => n3811);
   U2803 : NAND2_X1 port map( A1 => DataP_alu_a_in_26_port, A2 => n3894, ZN => 
                           n3808);
   U2804 : OAI211_X1 port map( C1 => DataP_alu_a_in_26_port, C2 => n3894, A => 
                           DataP_alu_b_in_26_port, B => n3838, ZN => n3809);
   U2805 : NAND2_X1 port map( A1 => n3719, A2 => n2584, ZN => n3807);
   U2806 : OAI211_X1 port map( C1 => n2216, C2 => n2756, A => n2574, B => n2482
                           , ZN => n2774);
   U2807 : INV_X1 port map( A => n2756, ZN => n2575);
   U2808 : INV_X1 port map( A => DataP_npc_31_port, ZN => n4191);
   U2809 : NAND2_X1 port map( A1 => n1721, A2 => n2754, ZN => n2753);
   U2810 : OAI21_X1 port map( B1 => n3905, B2 => n3902, A => n3901, ZN => n3903
                           );
   U2811 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N81, B2 => n3227, A => 
                           n3899, ZN => n3901);
   U2812 : OAI21_X1 port map( B1 => n3898, B2 => n3897, A => n3896, ZN => n3899
                           );
   U2813 : AOI22_X1 port map( A1 => DataP_alu_a_in_31_port, A2 => n3895, B1 => 
                           n3894, B2 => DataP_alu_b_in_31_port, ZN => n3896);
   U2814 : NAND2_X1 port map( A1 => DataP_alu_b_in_31_port, A2 => n3890, ZN => 
                           n3893);
   U2815 : NOR2_X1 port map( A1 => n3905, A2 => n2750, ZN => n2749);
   U2816 : NOR2_X1 port map( A1 => n2754, A2 => n3905, ZN => n2751);
   U2817 : NAND2_X1 port map( A1 => n3888, A2 => n2129, ZN => n3905);
   U2818 : INV_X1 port map( A => n3889, ZN => n3888);
   U2819 : AOI21_X1 port map( B1 => n2663, B2 => n2129, A => n3704, ZN => n301)
                           ;
   U2820 : INV_X1 port map( A => DataP_npc_23_port, ZN => n4199);
   U2821 : OAI211_X1 port map( C1 => n3678, C2 => n3892, A => n3677, B => n3676
                           , ZN => n3679);
   U2822 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N41, A2 => n3228, ZN =>
                           n3676);
   U2823 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N73, B2 => n3227, A => 
                           n3675, ZN => n3677);
   U2824 : OAI211_X1 port map( C1 => n4108, C2 => n3897, A => n3674, B => n3673
                           , ZN => n3675);
   U2825 : NAND2_X1 port map( A1 => DataP_alu_a_in_23_port, A2 => n3894, ZN => 
                           n3673);
   U2826 : OAI211_X1 port map( C1 => DataP_alu_a_in_23_port, C2 => n3894, A => 
                           DataP_alu_b_in_23_port, B => n3838, ZN => n3674);
   U2827 : INV_X1 port map( A => DataP_ALU_C_shifter_N105, ZN => n3678);
   U2828 : INV_X1 port map( A => n3125, ZN => n3196);
   U2829 : INV_X1 port map( A => n1717, ZN => n3672);
   U2830 : NAND2_X1 port map( A1 => n2763, A2 => n2761, ZN => n2760);
   U2831 : NOR2_X1 port map( A1 => n3680, A2 => n2762, ZN => n2761);
   U2832 : INV_X1 port map( A => n3683, ZN => n2762);
   U2833 : INV_X1 port map( A => DataP_npc_28_port, ZN => n4194);
   U2834 : OAI211_X1 port map( C1 => n3892, C2 => n3137, A => n3823, B => n3822
                           , ZN => n3824);
   U2835 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N78, B2 => n3227, A => 
                           n3821, ZN => n3822);
   U2836 : OAI21_X1 port map( B1 => n3897, B2 => n3820, A => n3819, ZN => n3821
                           );
   U2837 : AOI22_X1 port map( A1 => n3818, A2 => DataP_alu_b_in_28_port, B1 => 
                           n3894, B2 => DataP_alu_a_in_28_port, ZN => n3819);
   U2838 : OAI21_X1 port map( B1 => n3817, B2 => n3851, A => n3891, ZN => n3818
                           );
   U2839 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N46, A2 => n3228, ZN =>
                           n3823);
   U2840 : INV_X1 port map( A => n3798, ZN => n2747);
   U2841 : OAI22_X1 port map( A1 => n304, A2 => n4111, B1 => n4110, B2 => n4197
                           , ZN => DataP_PC_reg_N27);
   U2842 : INV_X1 port map( A => DataP_npc_25_port, ZN => n4197);
   U2843 : AOI21_X1 port map( B1 => n3806, B2 => n2129, A => n3805, ZN => n304)
                           ;
   U2844 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N75, B2 => n3227, A => 
                           n3801, ZN => n3802);
   U2845 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N43, A2 => n3228, ZN =>
                           n3803);
   U2846 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N107, A2 => n3877, ZN 
                           => n3804);
   U2847 : INV_X1 port map( A => n3130, ZN => n3198);
   U2848 : OAI22_X1 port map( A1 => n330, A2 => n4111, B1 => n4110, B2 => n4207
                           , ZN => DataP_PC_reg_N17);
   U2849 : INV_X1 port map( A => DataP_npc_15_port, ZN => n4207);
   U2850 : AOI21_X1 port map( B1 => n2689, B2 => n2129, A => n2688, ZN => n330)
                           ;
   U2851 : NAND2_X1 port map( A1 => n3626, A2 => n3627, ZN => n2688);
   U2852 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N65, B2 => n3900, A => 
                           n3625, ZN => n3627);
   U2853 : OAI211_X1 port map( C1 => n3624, C2 => n3891, A => n3623, B => n3622
                           , ZN => n3625);
   U2854 : OAI211_X1 port map( C1 => DataP_alu_a_in_15_port, C2 => n3894, A => 
                           DataP_alu_b_in_15_port, B => n3838, ZN => n3622);
   U2855 : NAND2_X1 port map( A1 => n3621, A2 => n2130, ZN => n3623);
   U2856 : AOI22_X1 port map( A1 => DataP_ALU_C_shifter_N33, A2 => n3228, B1 =>
                           n3877, B2 => DataP_ALU_C_shifter_N97, ZN => n3626);
   U2857 : INV_X1 port map( A => n2894, ZN => n2907);
   U2858 : INV_X1 port map( A => DataP_npc_29_port, ZN => n4193);
   U2859 : OAI211_X1 port map( C1 => n3892, C2 => n3139, A => n3832, B => n3831
                           , ZN => n3833);
   U2860 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N79, B2 => n3227, A => 
                           n3830, ZN => n3831);
   U2861 : OAI21_X1 port map( B1 => n3897, B2 => n3829, A => n3828, ZN => n3830
                           );
   U2862 : AOI22_X1 port map( A1 => n3827, A2 => DataP_alu_b_in_29_port, B1 => 
                           n3894, B2 => DataP_alu_a_in_29_port, ZN => n3828);
   U2863 : OAI21_X1 port map( B1 => n2365, B2 => n3851, A => n3891, ZN => n3827
                           );
   U2864 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N47, A2 => n3904, ZN =>
                           n3832);
   U2865 : AND2_X1 port map( A1 => n2766, A2 => n2748, ZN => n2717);
   U2866 : AOI21_X1 port map( B1 => n2756, B2 => n2131, A => n2474, ZN => n2707
                           );
   U2867 : INV_X1 port map( A => DataP_npc_30_port, ZN => n4192);
   U2868 : NAND2_X1 port map( A1 => DataP_alu_a_in_30_port, A2 => n3894, ZN => 
                           n3705);
   U2869 : OAI211_X1 port map( C1 => DataP_alu_a_in_30_port, C2 => n3894, A => 
                           DataP_alu_b_in_30_port, B => n3838, ZN => n3706);
   U2870 : NAND2_X1 port map( A1 => n3891, A2 => n3851, ZN => n3838);
   U2871 : OR2_X1 port map( A1 => n3880, A2 => n4111, ZN => n2708);
   U2872 : AOI21_X1 port map( B1 => n3713, B2 => n1548, A => n3788, ZN => n3717
                           );
   U2873 : AND2_X1 port map( A1 => n3715, A2 => n1717, ZN => n2726);
   U2874 : NOR2_X1 port map( A1 => n3725, A2 => n3798, ZN => n2748);
   U2875 : NAND2_X1 port map( A1 => n3711, A2 => DataP_alu_a_in_30_port, ZN => 
                           n3884);
   U2876 : INV_X1 port map( A => n3710, ZN => n3711);
   U2877 : NAND2_X1 port map( A1 => n3710, A2 => n2364, ZN => n3902);
   U2878 : OAI21_X1 port map( B1 => n2566, B2 => n2535, A => n2565, ZN => n3710
                           );
   U2879 : NAND2_X1 port map( A1 => n2614, A2 => n2535, ZN => n2565);
   U2880 : XNOR2_X1 port map( A => n2567, B => DataP_alu_b_in_30_port, ZN => 
                           n2566);
   U2881 : NOR2_X1 port map( A1 => n3722, A2 => n2381, ZN => n2567);
   U2882 : INV_X1 port map( A => n3728, ZN => n3727);
   U2883 : NOR2_X1 port map( A1 => n3724, A2 => DataP_alu_a_in_28_port, ZN => 
                           n2765);
   U2884 : INV_X1 port map( A => n3816, ZN => n3724);
   U2885 : NOR2_X1 port map( A1 => n3816, A2 => n3817, ZN => n3725);
   U2886 : INV_X1 port map( A => DataP_alu_a_in_28_port, ZN => n3817);
   U2887 : XNOR2_X1 port map( A => n3722, B => DataP_alu_b_in_28_port, ZN => 
                           n3723);
   U2888 : NAND2_X1 port map( A1 => n3709, A2 => n3726, ZN => n3722);
   U2889 : NOR2_X1 port map( A1 => n3708, A2 => DataP_alu_b_in_27_port, ZN => 
                           n3726);
   U2890 : AOI21_X1 port map( B1 => n3704, B2 => n2131, A => n2592, ZN => n2591
                           );
   U2891 : NOR2_X1 port map( A1 => n4110, A2 => n4195, ZN => n2592);
   U2892 : INV_X1 port map( A => DataP_npc_27_port, ZN => n4195);
   U2893 : OAI211_X1 port map( C1 => n3892, C2 => n3135, A => n3703, B => n3702
                           , ZN => n3704);
   U2894 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N77, B2 => n3227, A => 
                           n3701, ZN => n3702);
   U2895 : OAI21_X1 port map( B1 => n3897, B2 => n3700, A => n3699, ZN => n3701
                           );
   U2896 : AOI22_X1 port map( A1 => n3698, A2 => DataP_alu_b_in_27_port, B1 => 
                           n3894, B2 => DataP_alu_a_in_27_port, ZN => n3699);
   U2897 : OAI21_X1 port map( B1 => n3697, B2 => n3851, A => n3891, ZN => n3698
                           );
   U2898 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N45, A2 => n3228, ZN =>
                           n3703);
   U2899 : INV_X1 port map( A => n3708, ZN => n2703);
   U2900 : NAND2_X1 port map( A1 => n2485, A2 => n2127, ZN => n3708);
   U2901 : AND2_X1 port map( A1 => n2588, A2 => n2107, ZN => n2485);
   U2902 : AOI21_X1 port map( B1 => n2389, B2 => n2715, A => n2706, ZN => n2705
                           );
   U2903 : INV_X1 port map( A => n3696, ZN => n2706);
   U2904 : OAI21_X1 port map( B1 => n3798, B2 => n2727, A => n3797, ZN => n3696
                           );
   U2905 : NAND2_X1 port map( A1 => DataP_alu_b_in_23_port, A2 => n2535, ZN => 
                           n2701);
   U2906 : NAND2_X1 port map( A1 => n3692, A2 => n2122, ZN => n2702);
   U2907 : INV_X1 port map( A => DataP_alu_a_in_22_port, ZN => n3778);
   U2908 : AND2_X1 port map( A1 => n3683, A2 => n2239, ZN => n3730);
   U2909 : NAND2_X1 port map( A1 => n3646, A2 => n3645, ZN => n3683);
   U2910 : INV_X1 port map( A => DataP_alu_a_in_16_port, ZN => n3645);
   U2911 : NAND2_X1 port map( A1 => n3763, A2 => n1588, ZN => n2606);
   U2912 : XNOR2_X1 port map( A => n1574, B => DataP_alu_b_in_24_port, ZN => 
                           n3695);
   U2913 : INV_X1 port map( A => n3668, ZN => n3692);
   U2914 : NAND2_X1 port map( A1 => n2679, A2 => n3886, ZN => n2676);
   U2915 : INV_X1 port map( A => n2679, ZN => n2598);
   U2916 : AND3_X1 port map( A1 => n2224, A2 => n3714, A3 => n3680, ZN => n3681
                           );
   U2917 : NAND2_X1 port map( A1 => n2402, A2 => n3886, ZN => n2569);
   U2918 : NAND2_X1 port map( A1 => n3663, A2 => n3664, ZN => n3668);
   U2919 : NOR2_X1 port map( A1 => DataP_alu_a_in_18_port, A2 => n2548, ZN => 
                           n2547);
   U2920 : INV_X1 port map( A => n2757, ZN => n2548);
   U2921 : NAND2_X1 port map( A1 => n2732, A2 => n2731, ZN => n2730);
   U2922 : INV_X1 port map( A => DataP_alu_b_in_19_port, ZN => n2732);
   U2923 : OR2_X1 port map( A1 => n2244, A2 => n2486, ZN => n2733);
   U2924 : OR2_X1 port map( A1 => n2135, A2 => n2757, ZN => n2524);
   U2925 : NAND2_X1 port map( A1 => n2546, A2 => n2526, ZN => n2525);
   U2926 : NOR2_X1 port map( A1 => n2135, A2 => n2535, ZN => n2526);
   U2927 : NAND2_X1 port map( A1 => n2301, A2 => n1753, ZN => n3659);
   U2928 : NAND2_X1 port map( A1 => n3616, A2 => n3615, ZN => n3638);
   U2929 : AND2_X1 port map( A1 => DataP_alu_a_in_15_port, A2 => n2108, ZN => 
                           n3615);
   U2930 : NAND2_X1 port map( A1 => n3614, A2 => n2479, ZN => n2577);
   U2931 : INV_X1 port map( A => DataP_alu_a_in_15_port, ZN => n3624);
   U2932 : INV_X1 port map( A => n3616, ZN => n3614);
   U2933 : NAND2_X1 port map( A1 => n3633, A2 => n3632, ZN => n2724);
   U2934 : AND2_X1 port map( A1 => n2647, A2 => n2643, ZN => n2642);
   U2935 : AND2_X1 port map( A1 => n3632, A2 => n1739, ZN => n2611);
   U2936 : INV_X1 port map( A => n3632, ZN => n3636);
   U2937 : INV_X1 port map( A => n3630, ZN => n3868);
   U2938 : NAND2_X1 port map( A1 => n3628, A2 => n3865, ZN => n3861);
   U2939 : OAI22_X1 port map( A1 => n332, A2 => n4111, B1 => n4110, B2 => n4208
                           , ZN => DataP_PC_reg_N16);
   U2940 : INV_X1 port map( A => DataP_npc_14_port, ZN => n4208);
   U2941 : INV_X1 port map( A => n3882, ZN => n332);
   U2942 : OAI211_X1 port map( C1 => n3881, C2 => n3880, A => n3879, B => n3878
                           , ZN => n3882);
   U2943 : AOI22_X1 port map( A1 => DataP_ALU_C_shifter_N32, A2 => n3228, B1 =>
                           n3877, B2 => DataP_ALU_C_shifter_N96, ZN => n3878);
   U2944 : INV_X1 port map( A => n2890, ZN => n2906);
   U2945 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N64, B2 => n3227, A => 
                           n3876, ZN => n3879);
   U2946 : XNOR2_X1 port map( A => n3874, B => n3873, ZN => n3881);
   U2947 : AND2_X1 port map( A1 => n3631, A2 => n3632, ZN => n3873);
   U2948 : NOR2_X1 port map( A1 => n2652, A2 => n2650, ZN => n2649);
   U2949 : NOR2_X1 port map( A1 => n2390, A2 => n2108, ZN => n2650);
   U2950 : INV_X1 port map( A => n2390, ZN => n2651);
   U2951 : INV_X1 port map( A => n3629, ZN => n3867);
   U2952 : OAI21_X1 port map( B1 => n1713, B2 => n2738, A => n2393, ZN => n3630
                           );
   U2953 : NAND2_X1 port map( A1 => n2740, A2 => n2128, ZN => n2737);
   U2954 : XNOR2_X1 port map( A => n3618, B => n2106, ZN => n3619);
   U2955 : OAI21_X1 port map( B1 => n1597, B2 => n2736, A => n1726, ZN => n3863
                           );
   U2956 : INV_X1 port map( A => n2739, ZN => n2736);
   U2957 : INV_X1 port map( A => n3865, ZN => n3617);
   U2958 : NOR2_X1 port map( A1 => DataP_alu_b_in_11_port, A2 => 
                           DataP_alu_b_in_10_port, ZN => n3479);
   U2959 : AND2_X1 port map( A1 => n3491, A2 => n3490, ZN => n3628);
   U2960 : NAND2_X1 port map( A1 => n1714, A2 => n3463, ZN => n3491);
   U2961 : AND2_X1 port map( A1 => n2200, A2 => n2108, ZN => n3463);
   U2962 : INV_X1 port map( A => n2200, ZN => n3467);
   U2963 : XNOR2_X1 port map( A => n3461, B => n2151, ZN => n3462);
   U2964 : NAND2_X1 port map( A1 => n3460, A2 => n3459, ZN => n3461);
   U2965 : NAND2_X1 port map( A1 => n3485, A2 => n3484, ZN => n3486);
   U2966 : NAND2_X1 port map( A1 => n3447, A2 => n3451, ZN => n3484);
   U2967 : INV_X1 port map( A => DataP_alu_a_in_10_port, ZN => n3451);
   U2968 : OAI211_X1 port map( C1 => n3426, C2 => n3425, A => n3424, B => n3611
                           , ZN => n3487);
   U2969 : NAND2_X1 port map( A1 => n3855, A2 => n1655, ZN => n3424);
   U2970 : XNOR2_X1 port map( A => n3427, B => DataP_alu_a_in_7_port, ZN => 
                           n3611);
   U2971 : NAND2_X1 port map( A1 => n3608, A2 => n3606, ZN => n3425);
   U2972 : NAND2_X1 port map( A1 => n3422, A2 => DataP_alu_a_in_5_port, ZN => 
                           n3606);
   U2973 : INV_X1 port map( A => n1747, ZN => n3422);
   U2974 : NAND2_X1 port map( A1 => n3604, A2 => n3599, ZN => n3419);
   U2975 : NAND2_X1 port map( A1 => n3849, A2 => n3418, ZN => n3599);
   U2976 : INV_X1 port map( A => DataP_alu_a_in_4_port, ZN => n3418);
   U2977 : INV_X1 port map( A => n3414, ZN => n3415);
   U2978 : XNOR2_X1 port map( A => n3412, B => n1973, ZN => n3845);
   U2979 : AND2_X1 port map( A1 => n3598, A2 => n3597, ZN => n3420);
   U2980 : NAND2_X1 port map( A1 => n1589, A2 => n1973, ZN => n3597);
   U2981 : XNOR2_X1 port map( A => n3410, B => DataP_alu_b_in_3_port, ZN => 
                           n3411);
   U2982 : NOR2_X1 port map( A1 => DataP_alu_b_in_0_port, A2 => 
                           DataP_alu_b_in_1_port, ZN => n3416);
   U2983 : NAND2_X1 port map( A1 => n1712, A2 => DataP_alu_a_in_4_port, ZN => 
                           n3598);
   U2984 : NAND2_X1 port map( A1 => n2225, A2 => DataP_alu_a_in_8_port, ZN => 
                           n3835);
   U2985 : NAND2_X1 port map( A1 => n1610, A2 => DataP_alu_a_in_7_port, ZN => 
                           n3482);
   U2986 : INV_X1 port map( A => n1577, ZN => n3429);
   U2987 : INV_X1 port map( A => n3310, ZN => n2659);
   U2988 : INV_X1 port map( A => n3908, ZN => n3438);
   U2989 : AOI21_X1 port map( B1 => n3572, B2 => n2491, A => n2668, ZN => n296)
                           ;
   U2990 : OAI21_X1 port map( B1 => n2670, B2 => n2491, A => n2669, ZN => n2668
                           );
   U2991 : AOI21_X1 port map( B1 => DataP_ALU_C_shifter_N82, B2 => n3877, A => 
                           n3573, ZN => n2669);
   U2992 : NAND4_X1 port map( A1 => n3559, A2 => n3558, A3 => n3557, A4 => 
                           n3556, ZN => n3573);
   U2993 : OAI21_X1 port map( B1 => n3555, B2 => n3894, A => n3554, ZN => n3556
                           );
   U2994 : NAND2_X1 port map( A1 => n3435, A2 => n3561, ZN => n3891);
   U2995 : AOI21_X1 port map( B1 => n3880, B2 => n3897, A => n3577, ZN => n3555
                           );
   U2996 : NOR2_X1 port map( A1 => n3237, A2 => ALU_OPCODE_i_1_port, ZN => 
                           n3435);
   U2997 : NAND2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => n443, ZN => 
                           n3237);
   U2998 : INV_X1 port map( A => n3562, ZN => n3432);
   U2999 : XNOR2_X1 port map( A => ALU_OPCODE_i_2_port, B => n4100, ZN => n3407
                           );
   U3000 : NAND2_X1 port map( A1 => n3405, A2 => n3563, ZN => n3409);
   U3001 : OAI21_X1 port map( B1 => n443, B2 => ALU_OPCODE_i_3_port, A => n3562
                           , ZN => n3405);
   U3002 : NAND2_X1 port map( A1 => n1741, A2 => n3890, ZN => n3557);
   U3003 : OR2_X1 port map( A1 => n3434, A2 => n3562, ZN => n3851);
   U3004 : INV_X1 port map( A => n3433, ZN => n3434);
   U3005 : AND2_X1 port map( A1 => n3406, A2 => ALU_OPCODE_i_1_port, ZN => 
                           n3433);
   U3006 : NOR2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => n2491, ZN => 
                           n3406);
   U3007 : INV_X1 port map( A => n3561, ZN => n3430);
   U3008 : NAND2_X1 port map( A1 => DataP_ALU_C_shifter_N50, A2 => n3900, ZN =>
                           n3559);
   U3009 : NOR2_X1 port map( A1 => n3562, A2 => n4101, ZN => n3900);
   U3010 : INV_X1 port map( A => n4101, ZN => n3431);
   U3011 : NOR2_X1 port map( A1 => n3571, A2 => n3570, ZN => n2671);
   U3012 : OAI211_X1 port map( C1 => n3568, C2 => n2391, A => n3567, B => n3566
                           , ZN => n3572);
   U3013 : OAI21_X1 port map( B1 => n3565, B2 => n3571, A => n3564, ZN => n3566
                           );
   U3014 : INV_X1 port map( A => n3570, ZN => n3564);
   U3015 : NOR2_X1 port map( A1 => ALU_OPCODE_i_2_port, A2 => 
                           ALU_OPCODE_i_1_port, ZN => n3563);
   U3016 : INV_X1 port map( A => DataP_ALU_C_comp_N50, ZN => n3565);
   U3017 : AOI22_X1 port map( A1 => DataP_ALU_C_comp_N50, A2 => n3560, B1 => 
                           n3561, B2 => n3571, ZN => n3568);
   U3018 : INV_X1 port map( A => n3569, ZN => n3571);
   U3019 : NAND2_X1 port map( A1 => n2683, A2 => n2682, ZN => n3560);
   U3020 : NAND2_X1 port map( A1 => n3561, A2 => ALU_OPCODE_i_1_port, ZN => 
                           n2682);
   U3021 : NAND2_X1 port map( A1 => n3569, A2 => n2684, ZN => n2683);
   U3022 : NOR2_X1 port map( A1 => n3562, A2 => ALU_OPCODE_i_1_port, ZN => 
                           n2684);
   U3023 : NAND2_X1 port map( A1 => n2672, A2 => ALU_OPCODE_i_0_port, ZN => 
                           n3562);
   U3024 : NAND2_X1 port map( A1 => n4103, A2 => n2741, ZN => n3569);
   U3025 : AND2_X1 port map( A1 => n2742, A2 => n4104, ZN => n2741);
   U3026 : NOR3_X1 port map( A1 => n3511, A2 => n3579, A3 => n3510, ZN => n4104
                           );
   U3027 : NAND4_X1 port map( A1 => n3829, A2 => n3820, A3 => n3700, A4 => 
                           n3810, ZN => n3510);
   U3028 : XNOR2_X1 port map( A => DataP_alu_a_in_26_port, B => 
                           DataP_alu_b_in_26_port, ZN => n3810);
   U3029 : XNOR2_X1 port map( A => DataP_alu_a_in_27_port, B => 
                           DataP_alu_b_in_27_port, ZN => n3700);
   U3030 : XNOR2_X1 port map( A => DataP_alu_a_in_28_port, B => 
                           DataP_alu_b_in_28_port, ZN => n3820);
   U3031 : XNOR2_X1 port map( A => DataP_alu_a_in_29_port, B => 
                           DataP_alu_b_in_29_port, ZN => n3829);
   U3032 : BUF_X1 port map( A => n3200, Z => n3201);
   U3033 : INV_X1 port map( A => n3800, ZN => n3511);
   U3034 : NOR2_X1 port map( A1 => n4105, A2 => n2743, ZN => n2742);
   U3035 : XNOR2_X1 port map( A => DataP_alu_a_in_22_port, B => 
                           DataP_alu_b_in_22_port, ZN => n3782);
   U3036 : XNOR2_X1 port map( A => DataP_alu_a_in_21_port, B => n2152, ZN => 
                           n3771);
   U3037 : XNOR2_X1 port map( A => DataP_alu_a_in_24_port, B => 
                           DataP_alu_b_in_24_port, ZN => n4109);
   U3038 : XNOR2_X1 port map( A => DataP_alu_a_in_23_port, B => 
                           DataP_alu_b_in_23_port, ZN => n4108);
   U3039 : XNOR2_X1 port map( A => DataP_alu_a_in_19_port, B => n1722, ZN => 
                           n4106);
   U3040 : XNOR2_X1 port map( A => DataP_alu_a_in_20_port, B => 
                           DataP_alu_b_in_20_port, ZN => n4107);
   U3041 : AND4_X1 port map( A1 => n3747, A2 => n3496, A3 => n3495, A4 => n3494
                           , ZN => n2434);
   U3042 : XNOR2_X1 port map( A => DataP_alu_a_in_9_port, B => n2166, ZN => 
                           n3494);
   U3043 : XNOR2_X1 port map( A => DataP_alu_a_in_10_port, B => n2165, ZN => 
                           n3495);
   U3044 : XNOR2_X1 port map( A => DataP_alu_a_in_12_port, B => 
                           lt_x_135_B_12_port, ZN => n3496);
   U3045 : XNOR2_X1 port map( A => DataP_alu_a_in_18_port, B => n1736, ZN => 
                           n3747);
   U3046 : XNOR2_X1 port map( A => DataP_alu_b_in_3_port, B => n1973, ZN => 
                           n3848);
   U3047 : INV_X1 port map( A => n3540, ZN => n3541);
   U3048 : XNOR2_X1 port map( A => DataP_alu_a_in_11_port, B => n3468, ZN => 
                           n3540);
   U3049 : INV_X1 port map( A => n2151, ZN => n3468);
   U3050 : AOI211_X1 port map( C1 => n3539, C2 => n3554, A => n3538, B => n3621
                           , ZN => n3542);
   U3051 : XNOR2_X1 port map( A => DataP_alu_a_in_15_port, B => n2230, ZN => 
                           n3621);
   U3052 : XNOR2_X1 port map( A => n3841, B => DataP_alu_a_in_8_port, ZN => 
                           n3538);
   U3053 : INV_X1 port map( A => n1575, ZN => n3841);
   U3054 : INV_X1 port map( A => n2231, ZN => n3537);
   U3055 : INV_X1 port map( A => n3577, ZN => n3539);
   U3056 : INV_X1 port map( A => n3591, ZN => n3536);
   U3057 : XNOR2_X1 port map( A => DataP_alu_a_in_2_port, B => n3052, ZN => 
                           n3591);
   U3058 : XNOR2_X1 port map( A => DataP_alu_a_in_4_port, B => n3055, ZN => 
                           n3853);
   U3059 : XNOR2_X1 port map( A => DataP_alu_a_in_6_port, B => 
                           DataP_alu_b_in_6_port, ZN => n3859);
   U3060 : XNOR2_X1 port map( A => DataP_alu_a_in_7_port, B => 
                           DataP_alu_b_in_7_port, ZN => n3613);
   U3061 : XNOR2_X1 port map( A => DataP_alu_a_in_13_port, B => n2141, ZN => 
                           n3872);
   U3062 : XNOR2_X1 port map( A => DataP_alu_a_in_16_port, B => 
                           DataP_alu_b_in_16_port, ZN => n3731);
   U3063 : XNOR2_X1 port map( A => n1751, B => DataP_alu_b_in_17_port, ZN => 
                           n3741);
   U3064 : XNOR2_X1 port map( A => DataP_alu_a_in_14_port, B => n2145, ZN => 
                           n3875);
   U3065 : INV_X1 port map( A => n3885, ZN => n3898);
   U3066 : XNOR2_X1 port map( A => DataP_alu_a_in_31_port, B => n2121, ZN => 
                           n3885);
   U3067 : XNOR2_X1 port map( A => DataP_alu_a_in_30_port, B => 
                           DataP_alu_b_in_30_port, ZN => n3707);
   U3068 : NOR2_X1 port map( A1 => n3216, A2 => n2447, ZN => n3381);
   U3069 : NOR2_X1 port map( A1 => n3216, A2 => n2455, ZN => n3384);
   U3070 : OAI21_X1 port map( B1 => n3214, B2 => n109, A => n3383, ZN => n3385)
                           ;
   U3071 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_18_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_18_port, ZN => n3383);
   U3072 : NAND4_X1 port map( A1 => n3553, A2 => n3552, A3 => n3551, A4 => 
                           n3550, ZN => DataP_alu_b_in_21_port);
   U3073 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_21_port, ZN =>
                           n3550);
   U3074 : OR2_X1 port map( A1 => n2771, A2 => n2419, ZN => n3551);
   U3075 : NAND2_X1 port map( A1 => n3223, A2 => DataP_IMM_s_21_port, ZN => 
                           n3552);
   U3076 : NAND2_X1 port map( A1 => n1572, A2 => DataP_B_s_21_port, ZN => n3553
                           );
   U3077 : NOR2_X1 port map( A1 => n3216, A2 => n2446, ZN => n3376);
   U3078 : OAI21_X1 port map( B1 => n3215, B2 => n121, A => n3375, ZN => n3377)
                           ;
   U3079 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_21_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_21_port, ZN => n3375);
   U3080 : NOR2_X1 port map( A1 => n3217, A2 => n2439, ZN => n3370);
   U3081 : OAI21_X1 port map( B1 => n3215, B2 => n129, A => n3369, ZN => n3371)
                           ;
   U3082 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_23_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_23_port, ZN => n3369);
   U3083 : NAND4_X1 port map( A1 => n3546, A2 => n3545, A3 => n3544, A4 => 
                           n3543, ZN => DataP_alu_b_in_23_port);
   U3084 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_23_port, ZN =>
                           n3543);
   U3085 : OR2_X1 port map( A1 => n1627, A2 => n2413, ZN => n3544);
   U3086 : NAND2_X1 port map( A1 => n1614, A2 => DataP_IMM_s_23_port, ZN => 
                           n3545);
   U3087 : NAND2_X1 port map( A1 => n1620, A2 => DataP_B_s_23_port, ZN => n3546
                           );
   U3088 : NOR2_X1 port map( A1 => n3217, A2 => n2464, ZN => n3373);
   U3089 : OAI21_X1 port map( B1 => n3213, B2 => n125, A => n3372, ZN => n3374)
                           ;
   U3090 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_22_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_22_port, ZN => n3372);
   U3091 : NOR2_X1 port map( A1 => n3216, A2 => n2454, ZN => n3379);
   U3092 : OAI21_X1 port map( B1 => n3215, B2 => n117, A => n3378, ZN => n3380)
                           ;
   U3093 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_20_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_20_port, ZN => n3378);
   U3094 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_20_port, ZN =>
                           n3497);
   U3095 : OR2_X1 port map( A1 => n2772, A2 => n2420, ZN => n3498);
   U3096 : NAND2_X1 port map( A1 => n2247, A2 => DataP_IMM_s_20_port, ZN => 
                           n3499);
   U3097 : NAND2_X1 port map( A1 => n3221, A2 => DataP_B_s_20_port, ZN => n3500
                           );
   U3098 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_16_port, ZN =>
                           n3532);
   U3099 : OR2_X1 port map( A1 => n2773, A2 => n2412, ZN => n3533);
   U3100 : NAND2_X1 port map( A1 => n3223, A2 => DataP_IMM_s_16_port, ZN => 
                           n3534);
   U3101 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_16_port, ZN => n3535
                           );
   U3102 : NOR2_X1 port map( A1 => n3216, A2 => n2465, ZN => n3387);
   U3103 : OAI21_X1 port map( B1 => n3215, B2 => n101, A => n3386, ZN => n3388)
                           ;
   U3104 : AOI22_X1 port map( A1 => n2209, A2 => DataP_alu_out_M_16_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_16_port, ZN => n3386);
   U3105 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_17_port, ZN =>
                           n3519);
   U3106 : OR2_X1 port map( A1 => n1627, A2 => n2416, ZN => n3520);
   U3107 : NAND2_X1 port map( A1 => n1623, A2 => DataP_IMM_s_17_port, ZN => 
                           n3521);
   U3108 : NAND2_X1 port map( A1 => n1645, A2 => DataP_B_s_17_port, ZN => n3522
                           );
   U3109 : AOI22_X1 port map( A1 => n3221, A2 => DataP_B_s_0_port, B1 => n3222,
                           B2 => DataP_IMM_s_0_port, ZN => n2656);
   U3110 : NOR2_X1 port map( A1 => n3218, A2 => n2461, ZN => n3333);
   U3111 : NOR2_X1 port map( A1 => n3218, A2 => n2460, ZN => n3331);
   U3112 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_2_port, ZN => 
                           n3311);
   U3113 : NOR2_X1 port map( A1 => n3218, A2 => n2459, ZN => n3329);
   U3114 : OAI21_X1 port map( B1 => n3215, B2 => n45, A => n3328, ZN => n3330);
   U3115 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_2_port, B1 => 
                           n3208, B2 => DataP_alu_out_W_2_port, ZN => n3328);
   U3116 : NAND2_X1 port map( A1 => n2246, A2 => DataP_IMM_s_3_port, ZN => 
                           n2661);
   U3117 : NAND2_X1 port map( A1 => n3220, A2 => DataP_B_s_3_port, ZN => n2662)
                           ;
   U3118 : NOR2_X1 port map( A1 => n3218, A2 => n2458, ZN => n3327);
   U3119 : NOR2_X1 port map( A1 => n3218, A2 => n2451, ZN => n3298);
   U3120 : OAI21_X1 port map( B1 => n3213, B2 => n65, A => n3297, ZN => n3299);
   U3121 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_7_port, B1 => 
                           n3208, B2 => DataP_alu_out_W_7_port, ZN => n3297);
   U3122 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_7_port, ZN => 
                           n3300);
   U3123 : NAND2_X1 port map( A1 => n3223, A2 => DataP_IMM_s_7_port, ZN => 
                           n3302);
   U3124 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_6_port, ZN => 
                           n3323);
   U3125 : OR2_X1 port map( A1 => n2773, A2 => n2410, ZN => n3324);
   U3126 : NOR2_X1 port map( A1 => n3218, A2 => n2462, ZN => n3342);
   U3127 : OAI21_X1 port map( B1 => n3213, B2 => n61, A => n3341, ZN => n3343);
   U3128 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_6_port, B1 => 
                           n3207, B2 => DataP_alu_out_W_6_port, ZN => n3341);
   U3129 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_4_port, ZN => 
                           n3315);
   U3130 : NOR2_X1 port map( A1 => n3217, A2 => n2443, ZN => n3339);
   U3131 : OAI21_X1 port map( B1 => n3215, B2 => n57, A => n3338, ZN => n3340);
   U3132 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_5_port, B1 => 
                           n3208, B2 => DataP_alu_out_W_5_port, ZN => n3338);
   U3133 : NOR2_X1 port map( A1 => n3214, A2 => n53, ZN => n3336);
   U3134 : OAI21_X1 port map( B1 => n3218, B2 => n2470, A => n3335, ZN => n3337
                           );
   U3135 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_4_port, B1 => 
                           n3208, B2 => DataP_alu_out_W_4_port, ZN => n3335);
   U3136 : OR2_X1 port map( A1 => n2072, A2 => n2518, ZN => n2692);
   U3137 : NOR2_X1 port map( A1 => n3216, A2 => n2449, ZN => n3399);
   U3138 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_11_port, ZN =>
                           n3454);
   U3139 : OR2_X1 port map( A1 => n2773, A2 => n2431, ZN => n3455);
   U3140 : NOR2_X1 port map( A1 => n3217, A2 => n2457, ZN => n3403);
   U3141 : OAI21_X1 port map( B1 => n3215, B2 => n77, A => n3400, ZN => n3404);
   U3142 : AOI22_X1 port map( A1 => n2209, A2 => DRAM_ADDRESS_10_port, B1 => 
                           n3209, B2 => DataP_alu_out_W_10_port, ZN => n3400);
   U3143 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_10_port, ZN =>
                           n3439);
   U3144 : OR2_X1 port map( A1 => n2773, A2 => n2409, ZN => n3440);
   U3145 : NOR2_X1 port map( A1 => n3213, A2 => n69, ZN => n3345);
   U3146 : OAI21_X1 port map( B1 => n3218, B2 => n2467, A => n3344, ZN => n3346
                           );
   U3147 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_8_port, B1 => 
                           n3208, B2 => DataP_alu_out_W_8_port, ZN => n3344);
   U3148 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_8_port, ZN => 
                           n3347);
   U3149 : OR2_X1 port map( A1 => n2773, A2 => n2408, ZN => n3348);
   U3150 : NAND4_X1 port map( A1 => n3527, A2 => n3526, A3 => n3525, A4 => 
                           n3524, ZN => DataP_alu_b_in_13_port);
   U3151 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_13_port, ZN =>
                           n3524);
   U3152 : OR2_X1 port map( A1 => n2772, A2 => n2423, ZN => n3525);
   U3153 : NAND2_X1 port map( A1 => n2247, A2 => DataP_IMM_s_13_port, ZN => 
                           n3526);
   U3154 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_13_port, ZN => n3527
                           );
   U3155 : NOR2_X1 port map( A1 => n3216, A2 => n2456, ZN => n3394);
   U3156 : OAI21_X1 port map( B1 => n3214, B2 => n89, A => n3393, ZN => n3395);
   U3157 : AOI22_X1 port map( A1 => n2209, A2 => DataP_alu_out_M_13_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_13_port, ZN => n3393);
   U3158 : NOR2_X1 port map( A1 => n3216, A2 => n2441, ZN => n3389);
   U3159 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_15_port, ZN =>
                           n3512);
   U3160 : OR2_X1 port map( A1 => n2771, A2 => n2433, ZN => n3513);
   U3161 : NAND2_X1 port map( A1 => n2246, A2 => DataP_IMM_s_15_port, ZN => 
                           n3514);
   U3162 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_15_port, ZN => n3515
                           );
   U3163 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_14_port, ZN =>
                           n3528);
   U3164 : OR2_X1 port map( A1 => n2773, A2 => n2418, ZN => n3529);
   U3165 : NAND2_X1 port map( A1 => n2246, A2 => DataP_IMM_s_14_port, ZN => 
                           n3530);
   U3166 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_14_port, ZN => n3531
                           );
   U3167 : NOR2_X1 port map( A1 => n3216, A2 => n2448, ZN => n3391);
   U3168 : OAI21_X1 port map( B1 => n3214, B2 => n93, A => n3390, ZN => n3392);
   U3169 : AOI22_X1 port map( A1 => n2209, A2 => DataP_alu_out_M_14_port, B1 =>
                           n3209, B2 => DataP_alu_out_W_14_port, ZN => n3390);
   U3170 : NOR2_X1 port map( A1 => n3216, A2 => n2442, ZN => n3397);
   U3171 : AOI22_X1 port map( A1 => n2209, A2 => DataP_alu_out_M_12_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_12_port, ZN => n3396);
   U3172 : BUF_X1 port map( A => n1762, Z => lt_x_135_B_12_port);
   U3173 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_12_port, ZN => n3478
                           );
   U3174 : OR2_X1 port map( A1 => n2773, A2 => n2424, ZN => n3476);
   U3175 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_12_port, ZN =>
                           n3475);
   U3176 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_9_port, ZN => 
                           n3260);
   U3177 : NAND2_X1 port map( A1 => n2247, A2 => DataP_IMM_s_9_port, ZN => 
                           n3262);
   U3178 : NAND4_X1 port map( A1 => n3523, A2 => n3509, A3 => n3508, A4 => 
                           n3507, ZN => DataP_alu_b_in_27_port);
   U3179 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_27_port, ZN =>
                           n3507);
   U3180 : OR2_X1 port map( A1 => n1627, A2 => n2411, ZN => n3508);
   U3181 : NAND2_X1 port map( A1 => n2227, A2 => DataP_B_s_27_port, ZN => n3509
                           );
   U3182 : NOR2_X1 port map( A1 => n3217, A2 => n2445, ZN => n3361);
   U3183 : OAI21_X1 port map( B1 => n3214, B2 => n141, A => n3360, ZN => n3362)
                           ;
   U3184 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_26_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_26_port, ZN => n3360);
   U3185 : NAND4_X1 port map( A1 => n3523, A2 => n3503, A3 => n3502, A4 => 
                           n3501, ZN => DataP_alu_b_in_26_port);
   U3186 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_26_port, ZN =>
                           n3501);
   U3187 : OR2_X1 port map( A1 => n1627, A2 => n2415, ZN => n3502);
   U3188 : NAND2_X1 port map( A1 => n2227, A2 => DataP_B_s_26_port, ZN => n3503
                           );
   U3189 : NOR2_X1 port map( A1 => n3217, A2 => n2453, ZN => n3364);
   U3190 : OAI21_X1 port map( B1 => n3214, B2 => n137, A => n3363, ZN => n3365)
                           ;
   U3191 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_25_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_25_port, ZN => n3363);
   U3192 : OR2_X1 port map( A1 => n2772, A2 => n2422, ZN => n3504);
   U3193 : NAND2_X1 port map( A1 => n3225, A2 => DataP_alu_out_W_25_port, ZN =>
                           n3505);
   U3194 : NAND2_X1 port map( A1 => n1645, A2 => DataP_B_s_25_port, ZN => n3506
                           );
   U3195 : NOR2_X1 port map( A1 => n3217, A2 => n2463, ZN => n3367);
   U3196 : OAI21_X1 port map( B1 => n3213, B2 => n133, A => n3366, ZN => n3368)
                           ;
   U3197 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_24_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_24_port, ZN => n3366);
   U3198 : NAND4_X1 port map( A1 => n3523, A2 => n3518, A3 => n3517, A4 => 
                           n3516, ZN => DataP_alu_b_in_31_port);
   U3199 : NAND2_X1 port map( A1 => n3224, A2 => DataP_alu_out_W_31_port, ZN =>
                           n3516);
   U3200 : OR2_X1 port map( A1 => n1627, A2 => n2414, ZN => n3517);
   U3201 : NAND2_X1 port map( A1 => n2227, A2 => DataP_B_s_31_port, ZN => n3518
                           );
   U3202 : NOR2_X1 port map( A1 => n2539, A2 => n2405, ZN => n2538);
   U3203 : NOR2_X1 port map( A1 => n3217, A2 => n2437, ZN => n3352);
   U3204 : OAI21_X1 port map( B1 => n3215, B2 => n157, A => n3351, ZN => n3353)
                           ;
   U3205 : AOI22_X1 port map( A1 => n3210, A2 => DataP_alu_out_M_30_port, B1 =>
                           n3208, B2 => DataP_alu_out_W_30_port, ZN => n3351);
   U3206 : NOR2_X1 port map( A1 => n3217, A2 => n2444, ZN => n3355);
   U3207 : OAI21_X1 port map( B1 => n3213, B2 => n153, A => n3354, ZN => n3356)
                           ;
   U3208 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_29_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_29_port, ZN => n3354);
   U3209 : NAND2_X1 port map( A1 => n2246, A2 => DataP_IMM_s_30_port, ZN => 
                           n3523);
   U3210 : NOR2_X1 port map( A1 => n3253, A2 => n3252, ZN => n3257);
   U3211 : XNOR2_X1 port map( A => DataP_Rs2_0_port, B => n528, ZN => n3253);
   U3212 : NOR2_X1 port map( A1 => n3255, A2 => n3254, ZN => n3256);
   U3213 : XNOR2_X1 port map( A => DataP_Rs2_2_port, B => n530, ZN => n3254);
   U3214 : XNOR2_X1 port map( A => DataP_Rs2_3_port, B => n2777, ZN => n3255);
   U3215 : NOR2_X1 port map( A1 => n3217, A2 => n2452, ZN => n3358);
   U3216 : OAI21_X1 port map( B1 => n3214, B2 => n149, A => n3357, ZN => n3359)
                           ;
   U3217 : AOI22_X1 port map( A1 => n3211, A2 => DataP_alu_out_M_28_port, B1 =>
                           n3207, B2 => DataP_alu_out_W_28_port, ZN => n3357);
   U3218 : NOR2_X1 port map( A1 => n3246, A2 => n3883, ZN => n2629);
   U3219 : INV_X1 port map( A => Rst, ZN => n2628);
   U3220 : AOI21_X1 port map( B1 => n3287, B2 => n17, A => n3286, ZN => n3296);
   U3221 : NOR2_X1 port map( A1 => n3285, A2 => n3284, ZN => n3286);
   U3222 : NOR2_X1 port map( A1 => n3280, A2 => n521, ZN => n3281);
   U3223 : NOR2_X1 port map( A1 => n3279, A2 => n3288, ZN => n3910);
   U3224 : NOR2_X1 port map( A1 => n3278, A2 => n3277, ZN => n3290);
   U3225 : NAND4_X1 port map( A1 => n3276, A2 => n3275, A3 => n3274, A4 => 
                           n3273, ZN => n3278);
   U3226 : XNOR2_X1 port map( A => n530, B => DataP_Rs1_2_port, ZN => n3270);
   U3227 : XNOR2_X1 port map( A => n528, B => n2392, ZN => n3268);
   U3228 : AOI21_X1 port map( B1 => n3265, B2 => n3264, A => n2091, ZN => n3288
                           );
   U3229 : NAND3_X1 port map( A1 => n3239, A2 => DataP_opcode_W_3_port, A3 => 
                           n2625, ZN => n2635);
   U3230 : NAND2_X1 port map( A1 => n2622, A2 => n2624, ZN => n3265);
   U3231 : AND2_X1 port map( A1 => n3902, A2 => n3884, ZN => n2376);
   U3232 : AND2_X1 port map( A1 => n1570, A2 => n2238, ZN => n2378);
   U3233 : OR2_X1 port map( A1 => DataP_alu_b_in_29_port, A2 => 
                           DataP_alu_b_in_28_port, ZN => n2381);
   U3234 : OAI211_X1 port map( C1 => n3621, C2 => n2108, A => n3638, B => n2577
                           , ZN => n2758);
   U3235 : OR2_X1 port map( A1 => n3217, A2 => n2436, ZN => n2384);
   U3236 : INV_X1 port map( A => n2740, ZN => n2738);
   U3237 : AND2_X1 port map( A1 => DataP_alu_a_in_21_port, A2 => n2679, ZN => 
                           n2388);
   U3238 : INV_X1 port map( A => n1618, ZN => n2754);
   U3239 : NOR2_X1 port map( A1 => n3430, A2 => n4101, ZN => n3904);
   U3240 : INV_X1 port map( A => n2165, ZN => n3459);
   U3241 : INV_X1 port map( A => n2233, ZN => n3046);
   U3242 : AND2_X1 port map( A1 => DataP_alu_a_in_13_port, A2 => n2737, ZN => 
                           n2393);
   U3243 : AND2_X1 port map( A1 => n2763, A2 => n2238, ZN => n2394);
   U3244 : AND2_X1 port map( A1 => n1723, A2 => n3762, ZN => n2396);
   U3245 : INV_X1 port map( A => n3851, ZN => n3890);
   U3246 : AND2_X1 port map( A1 => DataP_alu_a_in_17_port, A2 => n2721, ZN => 
                           n2397);
   U3247 : XOR2_X1 port map( A => n3816, B => n3817, Z => n2400);
   U3248 : INV_X1 port map( A => n3797, ZN => n2744);
   U3249 : INV_X1 port map( A => n3296, ZN => n2619);
   U3250 : NAND2_X1 port map( A1 => n3689, A2 => DataP_alu_a_in_23_port, ZN => 
                           n3715);
   U3251 : OR2_X1 port map( A1 => n2727, A2 => n3788, ZN => n2404);
   U3252 : NAND2_X1 port map( A1 => n3727, A2 => DataP_alu_a_in_29_port, ZN => 
                           n3825);
   U3253 : INV_X1 port map( A => n3825, ZN => n2746);
   U3254 : AND2_X1 port map( A1 => n3210, A2 => DataP_alu_out_M_31_port, ZN => 
                           n2405);
   U3255 : INV_X1 port map( A => n3826, ZN => n2750);
   U3256 : AND3_X1 port map( A1 => n3835, A2 => n3482, A3 => n3483, ZN => n2473
                           );
   U3257 : NOR2_X1 port map( A1 => n4110, A2 => n4192, ZN => n2474);
   U3258 : AND2_X1 port map( A1 => n2725, A2 => n2394, ZN => n2476);
   U3259 : AND2_X1 port map( A1 => n3624, A2 => n2108, ZN => n2479);
   U3260 : OR2_X1 port map( A1 => n2756, A2 => n2129, ZN => n2482);
   U3261 : NAND2_X1 port map( A1 => n2525, A2 => n2524, ZN => n3682);
   U3262 : NAND2_X1 port map( A1 => n3665, A2 => n2114, ZN => n3766);
   U3263 : INV_X1 port map( A => n3766, ZN => n2607);
   U3264 : INV_X1 port map( A => DataP_alu_b_in_30_port, ZN => n2614);
   U3265 : OR2_X1 port map( A1 => n1600, A2 => n2535, ZN => n2486);
   U3266 : AND2_X1 port map( A1 => DataP_alu_a_in_22_port, A2 => n2569, ZN => 
                           n2487);
   U3267 : AND2_X1 port map( A1 => n2755, A2 => n2749, ZN => n2488);
   U3268 : NAND2_X1 port map( A1 => n3720, A2 => DataP_alu_a_in_27_port, ZN => 
                           n3721);
   U3269 : OR2_X1 port map( A1 => n3825, A2 => n3826, ZN => n2489);
   U3270 : AND2_X1 port map( A1 => n2111, A2 => n2676, ZN => n2490);
   U3271 : INV_X1 port map( A => Rst, ZN => n3234);
   U3272 : NAND2_X1 port map( A1 => n3648, A2 => DataP_alu_a_in_19_port, ZN => 
                           n3685);
   U3273 : NAND2_X1 port map( A1 => n2615, A2 => n2733, ZN => n3648);
   U3274 : AND2_X1 port map( A1 => n1750, A2 => n2529, ZN => n2528);
   U3275 : NAND2_X1 port map( A1 => n2721, A2 => n2128, ZN => n2529);
   U3276 : INV_X1 port map( A => n3666, ZN => n3665);
   U3277 : OR2_X1 port map( A1 => n2630, A2 => n2598, ZN => n2530);
   U3278 : INV_X1 port map( A => n2653, ZN => n2532);
   U3279 : NAND4_X1 port map( A1 => n1734, A2 => n2219, A3 => n2220, A4 => 
                           n3684, ZN => n2533);
   U3280 : AOI21_X1 port map( B1 => n2536, B2 => n2129, A => n3775, ZN => n313)
                           ;
   U3281 : XNOR2_X1 port map( A => n2537, B => n2396, ZN => n2536);
   U3282 : AOI21_X1 port map( B1 => n3767, B2 => n3766, A => n3765, ZN => n2537
                           );
   U3283 : OAI22_X1 port map( A1 => n3213, A2 => n161, B1 => n2072, B2 => n2517
                           , ZN => n2539);
   U3284 : NAND2_X1 port map( A1 => DataP_alu_b_in_27_port, A2 => n2535, ZN => 
                           n2540);
   U3285 : XNOR2_X1 port map( A => n2541, B => n3635, ZN => n2689);
   U3286 : OAI21_X1 port map( B1 => n3874, B2 => n3636, A => n3631, ZN => n2541
                           );
   U3287 : AOI21_X1 port map( B1 => n2542, B2 => n3630, A => n3867, ZN => n3874
                           );
   U3288 : OAI21_X1 port map( B1 => n3864, B2 => n3617, A => n3863, ZN => n2542
                           );
   U3289 : AOI21_X1 port map( B1 => n2543, B2 => n2129, A => n3746, ZN => n323)
                           ;
   U3290 : XNOR2_X1 port map( A => n2544, B => n2155, ZN => n2543);
   U3291 : AOI21_X1 port map( B1 => n3729, B2 => n2238, A => n2545, ZN => n2544
                           );
   U3292 : INV_X1 port map( A => n1663, ZN => n2545);
   U3293 : OAI211_X1 port map( C1 => n4111, C2 => n2558, A => n2550, B => n2553
                           , ZN => DataP_PC_reg_N33);
   U3294 : INV_X1 port map( A => n2551, ZN => n2550);
   U3295 : OR2_X1 port map( A1 => n4110, A2 => n4191, ZN => n2552);
   U3296 : NAND2_X1 port map( A1 => n2554, A2 => n2131, ZN => n2553);
   U3297 : INV_X1 port map( A => n2556, ZN => n2554);
   U3298 : AND2_X1 port map( A1 => n2557, A2 => n2753, ZN => n2556);
   U3299 : NAND2_X1 port map( A1 => n2083, A2 => n2751, ZN => n2558);
   U3300 : NAND2_X1 port map( A1 => n2783, A2 => n1646, ZN => n3690);
   U3301 : NAND2_X1 port map( A1 => n2559, A2 => n2759, ZN => n3767);
   U3302 : NAND2_X1 port map( A1 => n2476, A2 => n2700, ZN => n2559);
   U3303 : AND2_X1 port map( A1 => n2724, A2 => n3635, ZN => n2700);
   U3304 : OAI22_X1 port map( A1 => n303, A2 => n4111, B1 => n4110, B2 => n4196
                           , ZN => DataP_PC_reg_N28);
   U3305 : AOI21_X1 port map( B1 => n2561, B2 => n2129, A => n3815, ZN => n303)
                           ;
   U3306 : XNOR2_X1 port map( A => n1711, B => n3807, ZN => n2561);
   U3307 : AOI21_X1 port map( B1 => n3824, B2 => n2131, A => n2563, ZN => n2562
                           );
   U3308 : NOR2_X1 port map( A1 => n4110, A2 => n4194, ZN => n2563);
   U3309 : NOR2_X1 port map( A1 => n3880, A2 => n4111, ZN => n2564);
   U3310 : NAND2_X1 port map( A1 => n3762, A2 => n3764, ZN => n3667);
   U3311 : NAND2_X1 port map( A1 => n3666, A2 => DataP_alu_a_in_20_port, ZN => 
                           n3764);
   U3312 : OAI21_X1 port map( B1 => n3886, B2 => n2678, A => n2388, ZN => n3762
                           );
   U3313 : NAND2_X1 port map( A1 => n2568, A2 => n2487, ZN => n3714);
   U3314 : NAND2_X1 port map( A1 => n3670, A2 => n2402, ZN => n2568);
   U3315 : XNOR2_X1 port map( A => n2570, B => n2122, ZN => n3670);
   U3316 : NOR2_X1 port map( A1 => n3668, A2 => n3669, ZN => n2570);
   U3317 : NAND2_X1 port map( A1 => n2576, A2 => n2571, ZN => n2709);
   U3318 : NAND3_X1 port map( A1 => n2595, A2 => n2376, A3 => n2070, ZN => 
                           n2571);
   U3319 : NAND2_X1 port map( A1 => n2595, A2 => n2572, ZN => n2574);
   U3320 : NOR2_X1 port map( A1 => n2719, A2 => n2573, ZN => n2572);
   U3321 : NAND2_X1 port map( A1 => n2376, A2 => n2575, ZN => n2573);
   U3322 : OAI21_X1 port map( B1 => n3215, B2 => n49, A => n2579, ZN => n2578);
   U3323 : AOI22_X1 port map( A1 => n3210, A2 => DRAM_ADDRESS_3_port, B1 => 
                           n3209, B2 => DataP_alu_out_W_3_port, ZN => n2579);
   U3324 : INV_X1 port map( A => n1635, ZN => n2580);
   U3325 : NAND2_X1 port map( A1 => n1564, A2 => n2747, ZN => n2581);
   U3326 : NAND2_X1 port map( A1 => n2584, A2 => n3721, ZN => n2582);
   U3327 : INV_X1 port map( A => n2096, ZN => n2584);
   U3328 : NAND2_X1 port map( A1 => n2587, A2 => n2108, ZN => n2586);
   U3329 : XNOR2_X1 port map( A => n2589, B => n2588, ZN => n2587);
   U3330 : NAND2_X1 port map( A1 => n1574, A2 => n2107, ZN => n2589);
   U3331 : NAND2_X1 port map( A1 => n2590, A2 => n2591, ZN => DataP_PC_reg_N29)
                           ;
   U3332 : NAND2_X1 port map( A1 => n2719, A2 => n2710, ZN => n2593);
   U3333 : XNOR2_X1 port map( A => n1594, B => DataP_alu_a_in_23_port, ZN => 
                           n3713);
   U3334 : OAI21_X1 port map( B1 => n2596, B2 => n2535, A => n2701, ZN => n3689
                           );
   U3335 : XNOR2_X1 port map( A => n2597, B => n2124, ZN => n2596);
   U3336 : NOR2_X1 port map( A1 => n3669, A2 => n2702, ZN => n2597);
   U3337 : OAI21_X1 port map( B1 => n2610, B2 => n3489, A => n2600, ZN => n3860
                           );
   U3338 : AOI21_X1 port map( B1 => n3486, B2 => n2601, A => n2235, ZN => n2600
                           );
   U3339 : NAND2_X1 port map( A1 => n3487, A2 => n2473, ZN => n2610);
   U3340 : NAND2_X1 port map( A1 => n3860, A2 => n3628, ZN => n3864);
   U3341 : INV_X1 port map( A => n3489, ZN => n2601);
   U3342 : NAND2_X1 port map( A1 => n2602, A2 => n3753, ZN => n2603);
   U3343 : AND2_X1 port map( A1 => n3766, A2 => n1588, ZN => n3753);
   U3344 : OAI211_X1 port map( C1 => n2604, C2 => n2607, A => n2603, B => n3686
                           , ZN => n2605);
   U3345 : OR2_X1 port map( A1 => n2606, A2 => n3687, ZN => n2604);
   U3346 : NAND2_X1 port map( A1 => n2605, A2 => n2608, ZN => n3716);
   U3347 : INV_X1 port map( A => n3776, ZN => n2608);
   U3348 : NAND2_X1 port map( A1 => n3688, A2 => n1717, ZN => n3776);
   U3349 : NAND2_X1 port map( A1 => n3671, A2 => n3778, ZN => n3688);
   U3350 : NAND3_X1 port map( A1 => n1745, A2 => n2609, A3 => n3634, ZN => 
                           n2725);
   U3351 : NAND3_X1 port map( A1 => n2610, A2 => n3488, A3 => n2222, ZN => 
                           n2609);
   U3352 : NAND2_X1 port map( A1 => n2430, A2 => n2613, ZN => n3887);
   U3353 : OAI21_X1 port map( B1 => n2385, B2 => n3722, A => n3885, ZN => n2613
                           );
   U3354 : AOI21_X1 port map( B1 => n3647, B2 => n2617, A => n2616, ZN => n2615
                           );
   U3355 : NAND2_X1 port map( A1 => n2730, A2 => n2734, ZN => n2616);
   U3356 : NAND2_X1 port map( A1 => n2618, A2 => n3909, ZN => n3212);
   U3357 : NAND2_X1 port map( A1 => n3295, A2 => n3296, ZN => n2618);
   U3358 : NAND2_X1 port map( A1 => n3293, A2 => n2629, ZN => n3295);
   U3359 : NAND2_X1 port map( A1 => n2085, A2 => n3258, ZN => n2781);
   U3360 : AND2_X1 port map( A1 => n3256, A2 => n3257, ZN => n2621);
   U3361 : NAND3_X1 port map( A1 => n2635, A2 => n2622, A3 => n2624, ZN => 
                           n2639);
   U3362 : NAND2_X1 port map( A1 => n2480, A2 => n2623, ZN => n2622);
   U3363 : XNOR2_X1 port map( A => n2779, B => n2383, ZN => n2623);
   U3364 : NAND2_X1 port map( A1 => n2483, A2 => DataP_opcode_W_1_port, ZN => 
                           n2624);
   U3365 : OAI211_X1 port map( C1 => DataP_opcode_W_0_port, C2 => 
                           DataP_opcode_W_4_port, A => DataP_opcode_W_2_port, B
                           => DataP_opcode_W_1_port, ZN => n2625);
   U3366 : OAI21_X1 port map( B1 => n2213, B2 => DataP_alu_b_in_20_port, A => 
                           n3663, ZN => n2630);
   U3367 : NAND2_X1 port map( A1 => n2152, A2 => n3664, ZN => n2631);
   U3368 : NAND4_X1 port map( A1 => n2634, A2 => n3292, A3 => n2633, A4 => 
                           n2632, ZN => n3402);
   U3369 : OR2_X1 port map( A1 => n3295, A2 => n1718, ZN => n2632);
   U3370 : AOI21_X1 port map( B1 => n3909, B2 => n2619, A => n2475, ZN => n2633
                           );
   U3371 : NAND2_X1 port map( A1 => n2635, A2 => DataP_opcode_W_5_port, ZN => 
                           n2638);
   U3372 : NAND4_X1 port map( A1 => n2640, A2 => n3244, A3 => n3243, A4 => 
                           n3242, ZN => n3289);
   U3373 : NOR2_X1 port map( A1 => n3241, A2 => n2641, ZN => n2640);
   U3374 : XNOR2_X1 port map( A => n2775, B => DataP_dest_M_3_port, ZN => n2641
                           );
   U3375 : AOI21_X1 port map( B1 => n3481, B2 => n1726, A => n2644, ZN => n2643
                           );
   U3376 : NAND2_X1 port map( A1 => n2646, A2 => n2645, ZN => n2644);
   U3377 : NAND2_X1 port map( A1 => n2393, A2 => n2738, ZN => n2645);
   U3378 : NAND2_X1 port map( A1 => n2735, A2 => n2736, ZN => n2646);
   U3379 : NAND2_X1 port map( A1 => n1713, A2 => n2393, ZN => n2647);
   U3380 : NAND2_X1 port map( A1 => n2648, A2 => n2649, ZN => n3632);
   U3381 : NAND2_X1 port map( A1 => n2685, A2 => n2651, ZN => n2648);
   U3382 : INV_X1 port map( A => DataP_alu_a_in_14_port, ZN => n2652);
   U3383 : NAND2_X1 port map( A1 => n2667, A2 => n2665, ZN => n2716);
   U3384 : NOR2_X1 port map( A1 => n3633, A2 => n2758, ZN => n2665);
   U3385 : NAND2_X1 port map( A1 => n2666, A2 => n3873, ZN => n3633);
   U3386 : NAND2_X1 port map( A1 => n3860, A2 => n1634, ZN => n2667);
   U3387 : NOR2_X1 port map( A1 => n3861, A2 => n3868, ZN => n3634);
   U3388 : NAND2_X1 port map( A1 => n3414, A2 => n2206, ZN => n3574);
   U3389 : NAND3_X1 port map( A1 => n2725, A2 => n2724, A3 => n3635, ZN => 
                           n2783);
   U3390 : NAND2_X1 port map( A1 => n2111, A2 => n2108, ZN => n2677);
   U3391 : NAND2_X1 port map( A1 => n3663, A2 => n3886, ZN => n2679);
   U3392 : NAND2_X1 port map( A1 => DataP_alu_b_in_6_port, A2 => n3886, ZN => 
                           n2680);
   U3393 : NAND2_X1 port map( A1 => n3841, A2 => n3886, ZN => n2686);
   U3394 : OAI211_X1 port map( C1 => n3215, C2 => n81, A => n2692, B => n2691, 
                           ZN => n2690);
   U3395 : NAND2_X1 port map( A1 => n2209, A2 => DRAM_ADDRESS_11_port, ZN => 
                           n2691);
   U3396 : AOI21_X1 port map( B1 => n2695, B2 => n2698, A => n2694, ZN => n2696
                           );
   U3397 : INV_X1 port map( A => n3686, ZN => n2694);
   U3398 : INV_X1 port map( A => n2759, ZN => n2695);
   U3399 : NAND4_X1 port map( A1 => n2700, A2 => n2223, A3 => n2394, A4 => 
                           n2698, ZN => n2697);
   U3400 : NOR2_X1 port map( A1 => n2699, A2 => n2607, ZN => n2698);
   U3401 : INV_X1 port map( A => n1723, ZN => n2699);
   U3402 : NAND3_X1 port map( A1 => n3889, A2 => n2129, A3 => n3902, ZN => 
                           n2704);
   U3403 : OAI21_X1 port map( B1 => n2709, B2 => n2708, A => n2707, ZN => 
                           DataP_PC_reg_N32);
   U3404 : INV_X1 port map( A => n2376, ZN => n2710);
   U3405 : NAND2_X1 port map( A1 => n1552, A2 => n1619, ZN => n2729);
   U3406 : NAND3_X1 port map( A1 => n2716, A2 => n2718, A3 => n2713, ZN => 
                           n2711);
   U3407 : NAND2_X1 port map( A1 => n2484, A2 => n2718, ZN => n2712);
   U3408 : AND2_X1 port map( A1 => n3712, A2 => n2714, ZN => n2713);
   U3409 : AOI21_X1 port map( B1 => n3635, B2 => n3636, A => n2715, ZN => n2714
                           );
   U3410 : INV_X1 port map( A => n3715, ZN => n2715);
   U3411 : OR2_X1 port map( A1 => DataP_alu_b_in_17_port, A2 => n2108, ZN => 
                           n2721);
   U3412 : NAND2_X1 port map( A1 => DataP_alu_b_in_26_port, A2 => n2535, ZN => 
                           n2722);
   U3413 : NOR2_X1 port map( A1 => n3693, A2 => n3694, ZN => n2723);
   U3414 : NAND2_X1 port map( A1 => n3716, A2 => n2726, ZN => n2728);
   U3415 : INV_X1 port map( A => n3718, ZN => n2727);
   U3416 : NAND2_X1 port map( A1 => n1600, A2 => n2535, ZN => n2734);
   U3417 : NAND2_X1 port map( A1 => n1573, A2 => n2128, ZN => n2739);
   U3418 : NAND2_X1 port map( A1 => n2141, A2 => n2128, ZN => n2740);
   U3419 : NAND2_X1 port map( A1 => n1736, A2 => n2535, ZN => n2757);
   U3420 : AND2_X1 port map( A1 => n1636, A2 => n2224, ZN => n2764);
   U3421 : AOI21_X1 port map( B1 => n3283, B2 => DataP_opcode_E_4_port, A => 
                           n17, ZN => n3285);
   U3422 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_0_port, ZN => 
                           n3308);
   U3423 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_3_port, ZN => 
                           n3310);
   U3424 : INV_X1 port map( A => n2782, ZN => n2771);
   U3425 : NAND2_X1 port map( A1 => n3221, A2 => DataP_B_s_8_port, ZN => n3350)
                           ;
   U3426 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_11_port, ZN => n3457
                           );
   U3427 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_2_port, ZN => n3314)
                           ;
   U3428 : NAND2_X1 port map( A1 => n3221, A2 => DataP_B_s_6_port, ZN => n3326)
                           ;
   U3429 : NAND2_X1 port map( A1 => n3221, A2 => DataP_B_s_9_port, ZN => n3263)
                           ;
   U3430 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_10_port, ZN => n3442
                           );
   U3431 : NAND2_X1 port map( A1 => n3220, A2 => DataP_B_s_4_port, ZN => n3318)
                           ;
   U3432 : NAND2_X1 port map( A1 => n3219, A2 => DataP_B_s_7_port, ZN => n3303)
                           ;
   U3433 : NAND2_X1 port map( A1 => n3220, A2 => DataP_B_s_5_port, ZN => n3322)
                           ;
   U3434 : OR2_X1 port map( A1 => n2773, A2 => n2450, ZN => n3320);
   U3435 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_5_port, ZN => 
                           n3319);
   U3436 : NAND2_X1 port map( A1 => n3763, A2 => n3667, ZN => n3686);
   U3437 : XNOR2_X1 port map( A => n2069, B => n2407, ZN => n3275);
   U3438 : XNOR2_X1 port map( A => n1638, B => n538, ZN => n3243);
   U3439 : NOR2_X1 port map( A1 => DataP_dest_M_4_port, A2 => n1621, ZN => 
                           n3249);
   U3440 : XNOR2_X1 port map( A => n2392, B => n1630, ZN => n3276);
   U3441 : XNOR2_X1 port map( A => n528, B => n536, ZN => n3242);
   U3442 : NAND2_X1 port map( A1 => n3238, A2 => DataP_opcode_W_5_port, ZN => 
                           n3239);
   U3443 : NAND2_X1 port map( A1 => n3226, A2 => DataP_alu_out_W_1_port, ZN => 
                           n3304);
   U3444 : XNOR2_X1 port map( A => n529, B => DataP_Rs1_1_port, ZN => n3269);
   U3445 : XNOR2_X1 port map( A => DataP_Rs2_1_port, B => n529, ZN => n3252);
   U3446 : XNOR2_X1 port map( A => n1628, B => n524, ZN => n3273);
   U3447 : XNOR2_X1 port map( A => DataP_dest_M_4_port, B => n540, ZN => n3241)
                           ;
   U3448 : AND2_X1 port map( A1 => n2220, A2 => n2167, ZN => n2784);
   U3449 : XNOR2_X1 port map( A => n2199, B => n2784, ZN => n3751);
   U3450 : XNOR2_X1 port map( A => DataP_add_D_1_port, B => n2429, ZN => n3277)
                           ;
   U3451 : XNOR2_X1 port map( A => DataP_add_D_1_port, B => DataP_Rs2_1_port, 
                           ZN => n3240);
   U3452 : XNOR2_X1 port map( A => DataP_dest_M_1_port, B => DataP_add_D_1_port
                           , ZN => n3244);
   U3453 : OAI21_X1 port map( B1 => DataP_opcode_W_1_port, B2 => 
                           DataP_opcode_W_2_port, A => DataP_opcode_W_4_port, 
                           ZN => n3238);
   U3454 : XNOR2_X1 port map( A => n3650, B => n2168, ZN => n3658);
   U3455 : NOR2_X1 port map( A1 => n21, A2 => DataP_opcode_E_0_port, ZN => 
                           n3282);
   U3456 : NAND2_X1 port map( A1 => n3537, A2 => n3199, ZN => n3554);
   U3457 : NAND2_X1 port map( A1 => n521, A2 => n520, ZN => n3283);
   U3458 : XNOR2_X1 port map( A => DataP_alu_a_in_5_port, B => 
                           lt_x_135_B_5_port, ZN => n3603);
   U3459 : INV_X1 port map( A => n2095, ZN => n3862);
   U3460 : NAND2_X1 port map( A1 => n3220, A2 => DataP_B_s_1_port, ZN => n3307)
                           ;
   U3461 : XNOR2_X1 port map( A => n1757, B => n523, ZN => n3274);
   U3462 : NAND2_X1 port map( A1 => n2780, A2 => n3258, ZN => n3549);
   U3463 : OAI21_X1 port map( B1 => n521, B2 => n3883, A => Rst, ZN => 
                           DataP_FORWARDING_BR_N12);
   U3464 : NAND2_X1 port map( A1 => n2248, A2 => n3272, ZN => n3294);
   U3465 : NOR2_X1 port map( A1 => DataP_opcode_M_2_port, A2 => 
                           DataP_opcode_M_1_port, ZN => n3247);
   U3466 : XNOR2_X1 port map( A => n2232, B => n3047, ZN => n3579);
   U3467 : OAI21_X1 port map( B1 => n521, B2 => n520, A => 
                           DataP_opcode_E_3_port, ZN => n3284);
   U3468 : OR2_X1 port map( A1 => n3293, A2 => n3291, ZN => n3292);
   U3469 : NAND2_X1 port map( A1 => n3416, A2 => n1716, ZN => n3410);
   U3470 : XNOR2_X1 port map( A => n2250, B => n1567, ZN => n3413);
   U3471 : NAND2_X1 port map( A1 => n2246, A2 => DataP_IMM_s_11_port, ZN => 
                           n3456);
   U3472 : NAND2_X1 port map( A1 => n1581, A2 => DataP_IMM_s_8_port, ZN => 
                           n3349);
   U3473 : NAND2_X1 port map( A1 => n3223, A2 => DataP_IMM_s_10_port, ZN => 
                           n3441);
   U3474 : NAND2_X1 port map( A1 => n3223, A2 => DataP_IMM_s_6_port, ZN => 
                           n3325);
   U3475 : NAND2_X1 port map( A1 => n2247, A2 => DataP_IMM_s_12_port, ZN => 
                           n3477);
   U3476 : OR2_X1 port map( A1 => n2773, A2 => n2477, ZN => n3261);
   U3477 : NAND2_X1 port map( A1 => n3222, A2 => DataP_IMM_s_4_port, ZN => 
                           n3317);
   U3478 : OR2_X1 port map( A1 => n2773, A2 => n2468, ZN => n3301);
   U3479 : OR2_X1 port map( A1 => n2771, A2 => n2466, ZN => n3316);
   U3480 : NAND2_X1 port map( A1 => n1581, A2 => DataP_IMM_s_2_port, ZN => 
                           n3313);
   U3481 : NAND2_X1 port map( A1 => n2247, A2 => DataP_IMM_s_5_port, ZN => 
                           n3321);
   U3482 : OR2_X1 port map( A1 => n2773, A2 => n2472, ZN => n3309);
   U3483 : NAND2_X1 port map( A1 => n3223, A2 => DataP_IMM_s_1_port, ZN => 
                           n3306);
   U3484 : OR2_X1 port map( A1 => n2773, A2 => n2469, ZN => n3305);
   U3485 : NAND4_X1 port map( A1 => n2201, A2 => n2918, A3 => n2126, A4 => 
                           n2916, ZN => n2853);
   U3486 : NOR2_X1 port map( A1 => n3204, A2 => n2853, ZN => n2810);
   U3487 : NAND2_X1 port map( A1 => n2231, A2 => n2916, ZN => n2785);
   U3488 : AOI22_X1 port map( A1 => n2103, A2 => n2232, B1 => 
                           DataP_alu_a_in_2_port, B2 => n2916, ZN => n2787);
   U3489 : AOI22_X1 port map( A1 => n2917, A2 => n2785, B1 => n2787, B2 => 
                           n2105, ZN => n2799);
   U3490 : NAND2_X1 port map( A1 => n2918, A2 => n2799, ZN => n2820);
   U3491 : AOI22_X1 port map( A1 => n2103, A2 => n1973, B1 => 
                           DataP_alu_a_in_4_port, B2 => n2916, ZN => n2786);
   U3492 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_5_port, B1 => 
                           DataP_alu_a_in_6_port, B2 => n2916, ZN => n2790);
   U3493 : AOI22_X1 port map( A1 => n2917, A2 => n2786, B1 => n2790, B2 => 
                           n2105, ZN => n2798);
   U3494 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_7_port, B1 => 
                           DataP_alu_a_in_8_port, B2 => n2916, ZN => n2789);
   U3495 : AOI22_X1 port map( A1 => n2103, A2 => n2207, B1 => 
                           DataP_alu_a_in_10_port, B2 => n2916, ZN => n2791);
   U3496 : AOI22_X1 port map( A1 => n2917, A2 => n2789, B1 => n2791, B2 => 
                           n2105, ZN => n2801);
   U3497 : AOI22_X1 port map( A1 => n3202, A2 => n2798, B1 => n2801, B2 => 
                           n3052, ZN => n2819);
   U3498 : AOI22_X1 port map( A1 => n3204, A2 => n2820, B1 => n2819, B2 => 
                           n2101, ZN => n2863);
   U3499 : AOI22_X1 port map( A1 => n2103, A2 => n2231, B1 => n2232, B2 => 
                           n2916, ZN => n2792);
   U3500 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_2_port, B1 => 
                           n1973, B2 => n2118, ZN => n2794);
   U3501 : AOI22_X1 port map( A1 => n2917, A2 => n2792, B1 => n2794, B2 => 
                           n2105, ZN => n2803);
   U3502 : NAND2_X1 port map( A1 => n2918, A2 => n2803, ZN => n2825);
   U3503 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_4_port, B1 => 
                           DataP_alu_a_in_5_port, B2 => n2916, ZN => n2793);
   U3504 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_6_port, B1 => 
                           DataP_alu_a_in_7_port, B2 => n2916, ZN => n2796);
   U3505 : AOI22_X1 port map( A1 => n2917, A2 => n2793, B1 => n2796, B2 => 
                           n2105, ZN => n2802);
   U3506 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_8_port, B1 => 
                           n2207, B2 => n2916, ZN => n2795);
   U3507 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_10_port, B1 => 
                           n2200, B2 => n2118, ZN => n2797);
   U3508 : AOI22_X1 port map( A1 => n2917, A2 => n2795, B1 => n2797, B2 => 
                           n2105, ZN => n2805);
   U3509 : AOI22_X1 port map( A1 => n3202, A2 => n2802, B1 => n2805, B2 => 
                           n3053, ZN => n2824);
   U3510 : AOI22_X1 port map( A1 => n2115, A2 => n2825, B1 => n2824, B2 => 
                           n2101, ZN => n2868);
   U3511 : NOR2_X1 port map( A1 => n3055, A2 => n2903, ZN => 
                           DataP_ALU_C_shifter_N29);
   U3512 : NOR2_X1 port map( A1 => n3050, A2 => n2785, ZN => n2788);
   U3513 : AOI22_X1 port map( A1 => n2917, A2 => n2787, B1 => n2786, B2 => 
                           n2105, ZN => n2807);
   U3514 : AOI22_X1 port map( A1 => n3202, A2 => n2788, B1 => n2807, B2 => 
                           n3052, ZN => n2831);
   U3515 : AOI22_X1 port map( A1 => n2917, A2 => n2790, B1 => n2789, B2 => 
                           n2105, ZN => n2806);
   U3516 : AOI22_X1 port map( A1 => n2103, A2 => n2200, B1 => 
                           DataP_alu_a_in_12_port, B2 => n2118, ZN => n2800);
   U3517 : AOI22_X1 port map( A1 => n3049, A2 => n2791, B1 => n2800, B2 => 
                           n2105, ZN => n2809);
   U3518 : AOI22_X1 port map( A1 => n3051, A2 => n2806, B1 => n2809, B2 => 
                           n3052, ZN => n2830);
   U3519 : AOI22_X1 port map( A1 => n2115, A2 => n2831, B1 => n2830, B2 => 
                           n2101, ZN => n2875);
   U3520 : NOR2_X1 port map( A1 => n2917, A2 => n2792, ZN => n2816);
   U3521 : AOI22_X1 port map( A1 => n2917, A2 => n2794, B1 => n2793, B2 => 
                           n2105, ZN => n2813);
   U3522 : AOI22_X1 port map( A1 => n3051, A2 => n2816, B1 => n2813, B2 => 
                           n3052, ZN => n2836);
   U3523 : AOI22_X1 port map( A1 => n2917, A2 => n2796, B1 => n2795, B2 => 
                           n2105, ZN => n2812);
   U3524 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_12_port, B1 => 
                           DataP_alu_a_in_13_port, B2 => n2118, ZN => n2804);
   U3525 : AOI22_X1 port map( A1 => n3050, A2 => n2797, B1 => n2804, B2 => 
                           n2105, ZN => n2815);
   U3526 : AOI22_X1 port map( A1 => n3202, A2 => n2812, B1 => n2815, B2 => 
                           n2919, ZN => n2835);
   U3527 : AOI22_X1 port map( A1 => n3204, A2 => n2836, B1 => n2835, B2 => 
                           n2101, ZN => n2882);
   U3528 : AOI22_X1 port map( A1 => n3202, A2 => n2799, B1 => n2798, B2 => 
                           n3053, ZN => n2841);
   U3529 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_13_port, B1 => 
                           DataP_alu_a_in_14_port, B2 => n2118, ZN => n2808);
   U3530 : AOI22_X1 port map( A1 => n2917, A2 => n2800, B1 => n2808, B2 => 
                           n2105, ZN => n2818);
   U3531 : AOI22_X1 port map( A1 => n3202, A2 => n2801, B1 => n2818, B2 => 
                           n3053, ZN => n2840);
   U3532 : AOI22_X1 port map( A1 => n2115, A2 => n2841, B1 => n2840, B2 => 
                           n2101, ZN => n2890);
   U3533 : NOR2_X1 port map( A1 => n3055, A2 => n2906, ZN => 
                           DataP_ALU_C_shifter_N32);
   U3534 : AOI22_X1 port map( A1 => n3202, A2 => n2803, B1 => n2802, B2 => 
                           n2919, ZN => n2846);
   U3535 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_14_port, B1 => 
                           DataP_alu_a_in_15_port, B2 => n2118, ZN => n2814);
   U3536 : AOI22_X1 port map( A1 => n2917, A2 => n2804, B1 => n2814, B2 => 
                           n2105, ZN => n2823);
   U3537 : AOI22_X1 port map( A1 => n3202, A2 => n2805, B1 => n2823, B2 => 
                           n3053, ZN => n2845);
   U3538 : AOI22_X1 port map( A1 => n2115, A2 => n2846, B1 => n2845, B2 => 
                           n2101, ZN => n2894);
   U3539 : NOR2_X1 port map( A1 => n3055, A2 => n2907, ZN => 
                           DataP_ALU_C_shifter_N33);
   U3540 : AOI22_X1 port map( A1 => n3202, A2 => n2807, B1 => n2806, B2 => 
                           n3053, ZN => n2852);
   U3541 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_15_port, B1 => 
                           DataP_alu_a_in_16_port, B2 => n2118, ZN => n2817);
   U3542 : AOI22_X1 port map( A1 => n3049, A2 => n2808, B1 => n2817, B2 => 
                           n2105, ZN => n2829);
   U3543 : AOI22_X1 port map( A1 => n3202, A2 => n2809, B1 => n2829, B2 => 
                           n3053, ZN => n2851);
   U3544 : AOI22_X1 port map( A1 => n2115, A2 => n2852, B1 => n2851, B2 => 
                           n2101, ZN => n2811);
   U3545 : MUX2_X1 port map( A => n2811, B => n2810, S => n2138, Z => 
                           DataP_ALU_C_shifter_N34);
   U3546 : AOI22_X1 port map( A1 => n3202, A2 => n2813, B1 => n2812, B2 => 
                           n2919, ZN => n2858);
   U3547 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_16_port, B1 => 
                           n1751, B2 => n2118, ZN => n2822);
   U3548 : AOI22_X1 port map( A1 => n3049, A2 => n2814, B1 => n2822, B2 => 
                           n2105, ZN => n2834);
   U3549 : AOI22_X1 port map( A1 => n3202, A2 => n2815, B1 => n2834, B2 => 
                           n2919, ZN => n2857);
   U3550 : NAND2_X1 port map( A1 => n2816, A2 => n3053, ZN => n2859);
   U3551 : NOR2_X1 port map( A1 => n3204, A2 => n2859, ZN => n2827);
   U3552 : AOI22_X1 port map( A1 => n2226, A2 => n1751, B1 => 
                           DataP_alu_a_in_18_port, B2 => n2118, ZN => n2828);
   U3553 : AOI22_X1 port map( A1 => n2917, A2 => n2817, B1 => n2828, B2 => 
                           n2105, ZN => n2839);
   U3554 : AOI22_X1 port map( A1 => n3202, A2 => n2818, B1 => n2839, B2 => 
                           n2919, ZN => n2862);
   U3555 : AOI22_X1 port map( A1 => n2115, A2 => n2819, B1 => n2862, B2 => 
                           n2101, ZN => n2821);
   U3556 : NOR2_X1 port map( A1 => n3204, A2 => n2820, ZN => n2884);
   U3557 : MUX2_X1 port map( A => n2821, B => n2884, S => n3055, Z => 
                           DataP_ALU_C_shifter_N36);
   U3558 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_18_port, B1 => 
                           DataP_alu_a_in_19_port, B2 => n2118, ZN => n2833);
   U3559 : AOI22_X1 port map( A1 => n2917, A2 => n2822, B1 => n2833, B2 => 
                           n2105, ZN => n2844);
   U3560 : AOI22_X1 port map( A1 => n3202, A2 => n2823, B1 => n2844, B2 => 
                           n2919, ZN => n2867);
   U3561 : AOI22_X1 port map( A1 => n2115, A2 => n2824, B1 => n2867, B2 => 
                           n2101, ZN => n2826);
   U3562 : NOR2_X1 port map( A1 => n3204, A2 => n2825, ZN => n2895);
   U3563 : MUX2_X1 port map( A => n2826, B => n2895, S => n3055, Z => 
                           DataP_ALU_C_shifter_N37);
   U3564 : NOR2_X1 port map( A1 => n3055, A2 => n2908, ZN => 
                           DataP_ALU_C_shifter_N19);
   U3565 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_19_port, B1 => 
                           DataP_alu_a_in_20_port, B2 => n2118, ZN => n2838);
   U3566 : AOI22_X1 port map( A1 => n3050, A2 => n2828, B1 => n2838, B2 => 
                           n2105, ZN => n2849);
   U3567 : AOI22_X1 port map( A1 => n3202, A2 => n2829, B1 => n2849, B2 => 
                           n2919, ZN => n2874);
   U3568 : AOI22_X1 port map( A1 => n2115, A2 => n2830, B1 => n2874, B2 => 
                           n2101, ZN => n2832);
   U3569 : NOR2_X1 port map( A1 => n3204, A2 => n2831, ZN => n2896);
   U3570 : MUX2_X1 port map( A => n2832, B => n2896, S => n3055, Z => 
                           DataP_ALU_C_shifter_N38);
   U3571 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_20_port, B1 => 
                           DataP_alu_a_in_21_port, B2 => n2118, ZN => n2843);
   U3572 : AOI22_X1 port map( A1 => n3050, A2 => n2833, B1 => n2843, B2 => 
                           n2105, ZN => n2856);
   U3573 : AOI22_X1 port map( A1 => n3202, A2 => n2834, B1 => n2856, B2 => 
                           n2919, ZN => n2881);
   U3574 : AOI22_X1 port map( A1 => n2115, A2 => n2835, B1 => n2881, B2 => 
                           n2101, ZN => n2837);
   U3575 : NOR2_X1 port map( A1 => n3204, A2 => n2836, ZN => n2897);
   U3576 : MUX2_X1 port map( A => n2837, B => n2897, S => n3055, Z => 
                           DataP_ALU_C_shifter_N39);
   U3577 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_21_port, B1 => 
                           DataP_alu_a_in_22_port, B2 => n2118, ZN => n2848);
   U3578 : AOI22_X1 port map( A1 => n2917, A2 => n2838, B1 => n2848, B2 => 
                           n2105, ZN => n2861);
   U3579 : AOI22_X1 port map( A1 => n3202, A2 => n2839, B1 => n2861, B2 => 
                           n2919, ZN => n2889);
   U3580 : AOI22_X1 port map( A1 => n2115, A2 => n2840, B1 => n2889, B2 => 
                           n2101, ZN => n2842);
   U3581 : NOR2_X1 port map( A1 => n3204, A2 => n2841, ZN => n2898);
   U3582 : MUX2_X1 port map( A => n2842, B => n2898, S => n3055, Z => 
                           DataP_ALU_C_shifter_N40);
   U3583 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_22_port, B1 => 
                           DataP_alu_a_in_23_port, B2 => n2118, ZN => n2855);
   U3584 : AOI22_X1 port map( A1 => n2917, A2 => n2843, B1 => n2855, B2 => 
                           n2105, ZN => n2865);
   U3585 : AOI22_X1 port map( A1 => n3202, A2 => n2844, B1 => n2865, B2 => 
                           n2919, ZN => n2893);
   U3586 : AOI22_X1 port map( A1 => n2115, A2 => n2845, B1 => n2893, B2 => 
                           n2101, ZN => n2847);
   U3587 : NOR2_X1 port map( A1 => n3204, A2 => n2846, ZN => n2899);
   U3588 : MUX2_X1 port map( A => n2847, B => n2899, S => n3055, Z => 
                           DataP_ALU_C_shifter_N41);
   U3589 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_23_port, B1 => 
                           DataP_alu_a_in_24_port, B2 => n2118, ZN => n2860);
   U3590 : AOI22_X1 port map( A1 => n2917, A2 => n2848, B1 => n2860, B2 => 
                           n2105, ZN => n2872);
   U3591 : AOI22_X1 port map( A1 => n3202, A2 => n2849, B1 => n2872, B2 => 
                           n2919, ZN => n2850);
   U3592 : AOI22_X1 port map( A1 => n2115, A2 => n2851, B1 => n2850, B2 => 
                           n2101, ZN => n2854);
   U3593 : AOI22_X1 port map( A1 => n2115, A2 => n2853, B1 => n2852, B2 => 
                           n2101, ZN => n2900);
   U3594 : MUX2_X1 port map( A => n2854, B => n2900, S => n2138, Z => 
                           DataP_ALU_C_shifter_N42);
   U3595 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_24_port, B1 => 
                           DataP_alu_a_in_25_port, B2 => n2118, ZN => n2864);
   U3596 : AOI22_X1 port map( A1 => n2917, A2 => n2855, B1 => n2864, B2 => 
                           n2105, ZN => n2879);
   U3597 : AOI22_X1 port map( A1 => n2115, A2 => n2859, B1 => n2858, B2 => 
                           n2101, ZN => n2901);
   U3598 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_25_port, B1 => 
                           DataP_alu_a_in_26_port, B2 => n2118, ZN => n2870);
   U3599 : AOI22_X1 port map( A1 => n2917, A2 => n2860, B1 => n2870, B2 => 
                           n2105, ZN => n2888);
   U3600 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_26_port, B1 => 
                           DataP_alu_a_in_27_port, B2 => n2118, ZN => n2877);
   U3601 : AOI22_X1 port map( A1 => n2917, A2 => n2864, B1 => n2877, B2 => 
                           n2105, ZN => n2892);
   U3602 : AOI22_X1 port map( A1 => n3202, A2 => n2865, B1 => n2892, B2 => 
                           n2918, ZN => n2866);
   U3603 : AOI22_X1 port map( A1 => n2115, A2 => n2867, B1 => n2866, B2 => 
                           n2101, ZN => n2869);
   U3604 : MUX2_X1 port map( A => n2869, B => n2868, S => n3055, Z => 
                           DataP_ALU_C_shifter_N45);
   U3605 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_27_port, B1 => 
                           DataP_alu_a_in_28_port, B2 => n2118, ZN => n2886);
   U3606 : AOI22_X1 port map( A1 => n2917, A2 => n2870, B1 => n2886, B2 => 
                           n2105, ZN => n2871);
   U3607 : AOI22_X1 port map( A1 => n3202, A2 => n2872, B1 => n2871, B2 => 
                           n2918, ZN => n2873);
   U3608 : AOI22_X1 port map( A1 => n2115, A2 => n2874, B1 => n2873, B2 => 
                           n2101, ZN => n2876);
   U3609 : MUX2_X1 port map( A => n2876, B => n2875, S => n3055, Z => 
                           DataP_ALU_C_shifter_N46);
   U3610 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_28_port, B1 => 
                           DataP_alu_a_in_29_port, B2 => n2118, ZN => n2891);
   U3611 : AOI22_X1 port map( A1 => n2917, A2 => n2877, B1 => n2891, B2 => 
                           n2105, ZN => n2878);
   U3612 : AOI22_X1 port map( A1 => n3051, A2 => n2879, B1 => n2878, B2 => 
                           n2918, ZN => n2880);
   U3613 : AOI22_X1 port map( A1 => n2115, A2 => n2881, B1 => n2880, B2 => 
                           n2101, ZN => n2883);
   U3614 : MUX2_X1 port map( A => n2883, B => n2882, S => n3055, Z => 
                           DataP_ALU_C_shifter_N47);
   U3615 : NOR2_X1 port map( A1 => n2138, A2 => n2909, ZN => 
                           DataP_ALU_C_shifter_N20);
   U3616 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_29_port, B1 => 
                           DataP_alu_a_in_30_port, B2 => n2118, ZN => n2885);
   U3617 : AOI22_X1 port map( A1 => n2917, A2 => n2886, B1 => n2885, B2 => 
                           n2105, ZN => n2887);
   U3618 : INV_X1 port map( A => n2126, ZN => n2917);
   U3619 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_15_port, B1 => 
                           DataP_alu_a_in_14_port, B2 => n2117, ZN => n2928);
   U3620 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_13_port, B1 => 
                           DataP_alu_a_in_12_port, B2 => n2117, ZN => n2931);
   U3621 : AOI22_X1 port map( A1 => n3049, A2 => n2928, B1 => n2931, B2 => 
                           n3047, ZN => n2939);
   U3622 : AOI22_X1 port map( A1 => n2103, A2 => n2200, B1 => 
                           DataP_alu_a_in_10_port, B2 => n2117, ZN => n2930);
   U3623 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_9_port, B1 => 
                           DataP_alu_a_in_8_port, B2 => n2117, ZN => n3000);
   U3624 : AOI22_X1 port map( A1 => n3050, A2 => n2930, B1 => n3000, B2 => 
                           n3047, ZN => n3017);
   U3625 : AOI22_X1 port map( A1 => n3051, A2 => n2939, B1 => n3017, B2 => 
                           n3053, ZN => n3038);
   U3626 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_7_port, B1 => 
                           DataP_alu_a_in_6_port, B2 => n2117, ZN => n2999);
   U3627 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_5_port, B1 => 
                           DataP_alu_a_in_4_port, B2 => n2117, ZN => n3002);
   U3628 : AOI22_X1 port map( A1 => n3049, A2 => n2999, B1 => n3002, B2 => 
                           n3047, ZN => n3016);
   U3629 : AOI22_X1 port map( A1 => n2103, A2 => n1973, B1 => 
                           DataP_alu_a_in_2_port, B2 => n2117, ZN => n3001);
   U3630 : AOI22_X1 port map( A1 => n2103, A2 => n2232, B1 => n2231, B2 => 
                           n2117, ZN => n2920);
   U3631 : AOI221_X1 port map( B1 => n3001, B2 => n3050, C1 => n2920, C2 => 
                           n3047, A => n3051, ZN => n2921);
   U3632 : AOI21_X1 port map( B1 => n3051, B2 => n3016, A => n2921, ZN => n2922
                           );
   U3633 : AOI22_X1 port map( A1 => n3204, A2 => n3038, B1 => n2922, B2 => 
                           n2101, ZN => n2923);
   U3634 : AOI22_X1 port map( A1 => n2226, A2 => DataP_alu_a_in_31_port, B1 => 
                           DataP_alu_a_in_30_port, B2 => n2117, ZN => n2932);
   U3635 : AOI22_X1 port map( A1 => n2226, A2 => DataP_alu_a_in_29_port, B1 => 
                           DataP_alu_a_in_28_port, B2 => n2117, ZN => n2934);
   U3636 : AOI22_X1 port map( A1 => n3049, A2 => n2932, B1 => n2934, B2 => 
                           n3201, ZN => n2982);
   U3637 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_27_port, B1 => 
                           DataP_alu_a_in_26_port, B2 => n2117, ZN => n2933);
   U3638 : AOI22_X1 port map( A1 => n2226, A2 => DataP_alu_a_in_25_port, B1 => 
                           DataP_alu_a_in_24_port, B2 => n2117, ZN => n2925);
   U3639 : AOI22_X1 port map( A1 => n3049, A2 => n2933, B1 => n2925, B2 => 
                           n3201, ZN => n2938);
   U3640 : AOI22_X1 port map( A1 => n3202, A2 => n2982, B1 => n2938, B2 => 
                           n3052, ZN => n2993);
   U3641 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_23_port, B1 => 
                           DataP_alu_a_in_22_port, B2 => n2117, ZN => n2924);
   U3642 : AOI22_X1 port map( A1 => n2226, A2 => DataP_alu_a_in_21_port, B1 => 
                           DataP_alu_a_in_20_port, B2 => n2117, ZN => n2927);
   U3643 : AOI22_X1 port map( A1 => n3050, A2 => n2924, B1 => n2927, B2 => 
                           n3047, ZN => n2937);
   U3644 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_19_port, B1 => 
                           DataP_alu_a_in_18_port, B2 => n2117, ZN => n2926);
   U3645 : AOI22_X1 port map( A1 => n2226, A2 => DataP_alu_a_in_17_port, B1 => 
                           DataP_alu_a_in_16_port, B2 => n2117, ZN => n2929);
   U3646 : AOI22_X1 port map( A1 => n3050, A2 => n2926, B1 => n2929, B2 => 
                           n3047, ZN => n2940);
   U3647 : AOI22_X1 port map( A1 => n3202, A2 => n2937, B1 => n2940, B2 => 
                           n3052, ZN => n3039);
   U3648 : AOI22_X1 port map( A1 => n2112, A2 => n2993, B1 => n3039, B2 => 
                           n2101, ZN => n2966);
   U3649 : MUX2_X1 port map( A => n2923, B => n2966, S => n3055, Z => 
                           DataP_ALU_C_shifter_N50);
   U3650 : AOI22_X1 port map( A1 => n3049, A2 => n2925, B1 => n2924, B2 => 
                           n3047, ZN => n2954);
   U3651 : AOI22_X1 port map( A1 => n3049, A2 => n2927, B1 => n2926, B2 => 
                           n3047, ZN => n2957);
   U3652 : AOI22_X1 port map( A1 => n3202, A2 => n2954, B1 => n2957, B2 => 
                           n3052, ZN => n2971);
   U3653 : AOI22_X1 port map( A1 => n3050, A2 => n2929, B1 => n2928, B2 => 
                           n3047, ZN => n2956);
   U3654 : AOI22_X1 port map( A1 => n3049, A2 => n2931, B1 => n2930, B2 => 
                           n3201, ZN => n3028);
   U3655 : AOI22_X1 port map( A1 => n3202, A2 => n2956, B1 => n3028, B2 => 
                           n3052, ZN => n3005);
   U3656 : AOI22_X1 port map( A1 => n2112, A2 => n2971, B1 => n3005, B2 => 
                           n2101, ZN => n2935);
   U3657 : NOR2_X1 port map( A1 => n3050, A2 => n2932, ZN => n2987);
   U3658 : AOI22_X1 port map( A1 => n3050, A2 => n2934, B1 => n2933, B2 => 
                           n3201, ZN => n2955);
   U3659 : AOI22_X1 port map( A1 => n3202, A2 => n2987, B1 => n2955, B2 => 
                           n3052, ZN => n2972);
   U3660 : NOR2_X1 port map( A1 => n2112, A2 => n2972, ZN => n2995);
   U3661 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_26_port, B1 => 
                           DataP_alu_a_in_25_port, B2 => n2117, ZN => n2943);
   U3662 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_24_port, B1 => 
                           DataP_alu_a_in_23_port, B2 => n2117, ZN => n2946);
   U3663 : AOI22_X1 port map( A1 => n3049, A2 => n2943, B1 => n2946, B2 => 
                           n3047, ZN => n2960);
   U3664 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_22_port, B1 => 
                           DataP_alu_a_in_21_port, B2 => n2117, ZN => n2945);
   U3665 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_20_port, B1 => 
                           DataP_alu_a_in_19_port, B2 => n2117, ZN => n2948);
   U3666 : AOI22_X1 port map( A1 => n3050, A2 => n2945, B1 => n2948, B2 => 
                           n3047, ZN => n2963);
   U3667 : AOI22_X1 port map( A1 => n3202, A2 => n2960, B1 => n2963, B2 => 
                           n3053, ZN => n2973);
   U3668 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_18_port, B1 => 
                           DataP_alu_a_in_17_port, B2 => n2117, ZN => n2947);
   U3669 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_16_port, B1 => 
                           DataP_alu_a_in_15_port, B2 => n2117, ZN => n2950);
   U3670 : AOI22_X1 port map( A1 => n3048, A2 => n2947, B1 => n2950, B2 => 
                           n3201, ZN => n2962);
   U3671 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_14_port, B1 => 
                           DataP_alu_a_in_13_port, B2 => n2117, ZN => n2949);
   U3672 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_12_port, B1 => 
                           n2200, B2 => n2117, ZN => n2975);
   U3673 : AOI22_X1 port map( A1 => n3048, A2 => n2949, B1 => n2975, B2 => 
                           n3201, ZN => n3034);
   U3674 : AOI22_X1 port map( A1 => n3202, A2 => n2962, B1 => n3034, B2 => 
                           n3053, ZN => n3014);
   U3675 : AOI22_X1 port map( A1 => n2112, A2 => n2973, B1 => n3014, B2 => 
                           n2101, ZN => n2936);
   U3676 : NAND2_X1 port map( A1 => DataP_alu_a_in_31_port, A2 => n2117, ZN => 
                           n2952);
   U3677 : NOR2_X1 port map( A1 => n3050, A2 => n2952, ZN => n2990);
   U3678 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_30_port, B1 => 
                           DataP_alu_a_in_29_port, B2 => n2117, ZN => n2951);
   U3679 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_28_port, B1 => 
                           DataP_alu_a_in_27_port, B2 => n2117, ZN => n2944);
   U3680 : AOI22_X1 port map( A1 => n3049, A2 => n2951, B1 => n2944, B2 => 
                           n3047, ZN => n2961);
   U3681 : AOI22_X1 port map( A1 => n3202, A2 => n2990, B1 => n2961, B2 => 
                           n3052, ZN => n2974);
   U3682 : NOR2_X1 port map( A1 => n2112, A2 => n2974, ZN => n2996);
   U3683 : MUX2_X1 port map( A => n2936, B => n2996, S => n3055, Z => 
                           DataP_ALU_C_shifter_N61);
   U3684 : NAND3_X1 port map( A1 => n2101, A2 => n3052, A3 => n2982, ZN => 
                           n2997);
   U3685 : AOI22_X1 port map( A1 => n3202, A2 => n2938, B1 => n2937, B2 => 
                           n3053, ZN => n2983);
   U3686 : AOI22_X1 port map( A1 => n3202, A2 => n2940, B1 => n2939, B2 => 
                           n3053, ZN => n3018);
   U3687 : AOI22_X1 port map( A1 => n2112, A2 => n2983, B1 => n3018, B2 => 
                           n2101, ZN => n2941);
   U3688 : NAND2_X1 port map( A1 => n2102, A2 => n2941, ZN => n2942);
   U3689 : AOI22_X1 port map( A1 => n3049, A2 => n2944, B1 => n2943, B2 => 
                           n3047, ZN => n2967);
   U3690 : AOI22_X1 port map( A1 => n3050, A2 => n2946, B1 => n2945, B2 => 
                           n3201, ZN => n2970);
   U3691 : AOI22_X1 port map( A1 => n3051, A2 => n2967, B1 => n2970, B2 => 
                           n3053, ZN => n2985);
   U3692 : AOI22_X1 port map( A1 => n3048, A2 => n2948, B1 => n2947, B2 => 
                           n3047, ZN => n2969);
   U3693 : AOI22_X1 port map( A1 => n3048, A2 => n2950, B1 => n2949, B2 => 
                           n3201, ZN => n2976);
   U3694 : AOI22_X1 port map( A1 => n3051, A2 => n2969, B1 => n2976, B2 => 
                           n3053, ZN => n3024);
   U3695 : AOI22_X1 port map( A1 => n2112, A2 => n2985, B1 => n3024, B2 => 
                           n2101, ZN => n2953);
   U3696 : AOI22_X1 port map( A1 => n3049, A2 => n2952, B1 => n2951, B2 => 
                           n3201, ZN => n2968);
   U3697 : NAND2_X1 port map( A1 => n3052, A2 => n2968, ZN => n2986);
   U3698 : NOR2_X1 port map( A1 => n2112, A2 => n2986, ZN => n2998);
   U3699 : NAND3_X1 port map( A1 => n2987, A2 => n2101, A3 => n3053, ZN => 
                           n3008);
   U3700 : AOI22_X1 port map( A1 => n3051, A2 => n2955, B1 => n2954, B2 => 
                           n3053, ZN => n2988);
   U3701 : AOI22_X1 port map( A1 => n3051, A2 => n2957, B1 => n2956, B2 => 
                           n3053, ZN => n3030);
   U3702 : AOI22_X1 port map( A1 => n2112, A2 => n2988, B1 => n3030, B2 => 
                           n2101, ZN => n2958);
   U3703 : NAND2_X1 port map( A1 => n3206, A2 => n2958, ZN => n2959);
   U3704 : OAI21_X1 port map( B1 => n2102, B2 => n3008, A => n2959, ZN => 
                           DataP_ALU_C_shifter_N64);
   U3705 : NAND3_X1 port map( A1 => n2990, A2 => n2101, A3 => n3052, ZN => 
                           n3009);
   U3706 : AOI22_X1 port map( A1 => n3051, A2 => n2961, B1 => n2960, B2 => 
                           n3053, ZN => n2991);
   U3707 : AOI22_X1 port map( A1 => n3051, A2 => n2963, B1 => n2962, B2 => 
                           n3053, ZN => n3035);
   U3708 : AOI22_X1 port map( A1 => n2115, A2 => n2991, B1 => n3035, B2 => 
                           n2101, ZN => n2964);
   U3709 : NAND2_X1 port map( A1 => n2102, A2 => n2964, ZN => n2965);
   U3710 : OAI21_X1 port map( B1 => n3206, B2 => n3009, A => n2965, ZN => 
                           DataP_ALU_C_shifter_N65);
   U3711 : AND2_X1 port map( A1 => n3206, A2 => n2966, ZN => 
                           DataP_ALU_C_shifter_N66);
   U3712 : AOI22_X1 port map( A1 => n3202, A2 => n2968, B1 => n2967, B2 => 
                           n3053, ZN => n2994);
   U3713 : AOI22_X1 port map( A1 => n3202, A2 => n2970, B1 => n2969, B2 => 
                           n3052, ZN => n3043);
   U3714 : AOI22_X1 port map( A1 => n3204, A2 => n2994, B1 => n3043, B2 => 
                           n2101, ZN => n2980);
   U3715 : AND2_X1 port map( A1 => n3206, A2 => n2980, ZN => 
                           DataP_ALU_C_shifter_N67);
   U3716 : AOI22_X1 port map( A1 => n3204, A2 => n2972, B1 => n2971, B2 => 
                           n2101, ZN => n3006);
   U3717 : AOI22_X1 port map( A1 => n2115, A2 => n2974, B1 => n2973, B2 => 
                           n2101, ZN => n3015);
   U3718 : AND2_X1 port map( A1 => n2102, A2 => n3015, ZN => 
                           DataP_ALU_C_shifter_N69);
   U3719 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_10_port, B1 => 
                           n2207, B2 => n2117, ZN => n3011);
   U3720 : AOI22_X1 port map( A1 => n3050, A2 => n2975, B1 => n3011, B2 => 
                           n3047, ZN => n3022);
   U3721 : AOI22_X1 port map( A1 => n3202, A2 => n2976, B1 => n3022, B2 => 
                           n3053, ZN => n3042);
   U3722 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_8_port, B1 => 
                           DataP_alu_a_in_7_port, B2 => n2117, ZN => n3010);
   U3723 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_6_port, B1 => 
                           DataP_alu_a_in_5_port, B2 => n2117, ZN => n3013);
   U3724 : AOI22_X1 port map( A1 => n3048, A2 => n3010, B1 => n3013, B2 => 
                           n3047, ZN => n3021);
   U3725 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_4_port, B1 => 
                           n1973, B2 => n2117, ZN => n3012);
   U3726 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_2_port, B1 => 
                           n2232, B2 => n2117, ZN => n2977);
   U3727 : AOI22_X1 port map( A1 => n3049, A2 => n3012, B1 => n2977, B2 => 
                           n3201, ZN => n2978);
   U3728 : AOI22_X1 port map( A1 => n3202, A2 => n3021, B1 => n2978, B2 => 
                           n3052, ZN => n2979);
   U3729 : AOI22_X1 port map( A1 => n3204, A2 => n3042, B1 => n2979, B2 => 
                           n2101, ZN => n2981);
   U3730 : MUX2_X1 port map( A => n2981, B => n2980, S => n3055, Z => 
                           DataP_ALU_C_shifter_N51);
   U3731 : NAND2_X1 port map( A1 => n3052, A2 => n2982, ZN => n2984);
   U3732 : AOI22_X1 port map( A1 => n3204, A2 => n2984, B1 => n2983, B2 => 
                           n2101, ZN => n3019);
   U3733 : AND2_X1 port map( A1 => n2102, A2 => n3019, ZN => 
                           DataP_ALU_C_shifter_N70);
   U3734 : AOI22_X1 port map( A1 => n3204, A2 => n2986, B1 => n2985, B2 => 
                           n2101, ZN => n3025);
   U3735 : AND2_X1 port map( A1 => n3206, A2 => n3025, ZN => 
                           DataP_ALU_C_shifter_N71);
   U3736 : NAND2_X1 port map( A1 => n2987, A2 => n3052, ZN => n2989);
   U3737 : AOI22_X1 port map( A1 => n3204, A2 => n2989, B1 => n2988, B2 => 
                           n2101, ZN => n3031);
   U3738 : AND2_X1 port map( A1 => n3206, A2 => n3031, ZN => 
                           DataP_ALU_C_shifter_N72);
   U3739 : NAND2_X1 port map( A1 => n2990, A2 => n3053, ZN => n2992);
   U3740 : AOI22_X1 port map( A1 => n3204, A2 => n2992, B1 => n2991, B2 => 
                           n2101, ZN => n3036);
   U3741 : AND2_X1 port map( A1 => n3206, A2 => n3036, ZN => 
                           DataP_ALU_C_shifter_N73);
   U3742 : NOR2_X1 port map( A1 => n2112, A2 => n2993, ZN => n3040);
   U3743 : AND2_X1 port map( A1 => n3040, A2 => n3206, ZN => 
                           DataP_ALU_C_shifter_N74);
   U3744 : NOR2_X1 port map( A1 => n2112, A2 => n2994, ZN => n3044);
   U3745 : AND2_X1 port map( A1 => n3044, A2 => n2102, ZN => 
                           DataP_ALU_C_shifter_N75);
   U3746 : AND2_X1 port map( A1 => n2995, A2 => n2102, ZN => 
                           DataP_ALU_C_shifter_N76);
   U3747 : AND2_X1 port map( A1 => n2996, A2 => n2102, ZN => 
                           DataP_ALU_C_shifter_N77);
   U3748 : NOR2_X1 port map( A1 => n3055, A2 => n2997, ZN => 
                           DataP_ALU_C_shifter_N78);
   U3749 : AND2_X1 port map( A1 => n2998, A2 => n2102, ZN => 
                           DataP_ALU_C_shifter_N79);
   U3750 : AOI22_X1 port map( A1 => n3048, A2 => n3000, B1 => n2999, B2 => 
                           n3201, ZN => n3027);
   U3751 : AOI22_X1 port map( A1 => n3048, A2 => n3002, B1 => n3001, B2 => 
                           n3047, ZN => n3003);
   U3752 : AOI22_X1 port map( A1 => n3202, A2 => n3027, B1 => n3003, B2 => 
                           n3052, ZN => n3004);
   U3753 : AOI22_X1 port map( A1 => n2115, A2 => n3005, B1 => n3004, B2 => 
                           n2101, ZN => n3007);
   U3754 : MUX2_X1 port map( A => n3007, B => n3006, S => n2138, Z => 
                           DataP_ALU_C_shifter_N52);
   U3755 : NOR2_X1 port map( A1 => n2138, A2 => n3008, ZN => 
                           DataP_ALU_C_shifter_N80);
   U3756 : NOR2_X1 port map( A1 => n3055, A2 => n3009, ZN => 
                           DataP_ALU_C_shifter_N81);
   U3757 : AOI22_X1 port map( A1 => n3049, A2 => n3011, B1 => n3010, B2 => 
                           n3047, ZN => n3033);
   U3758 : AOI22_X1 port map( A1 => n3051, A2 => n3022, B1 => n3021, B2 => 
                           n3052, ZN => n3023);
   U3759 : AOI22_X1 port map( A1 => n2112, A2 => n3024, B1 => n3023, B2 => 
                           n2101, ZN => n3026);
   U3760 : AOI22_X1 port map( A1 => n3051, A2 => n3028, B1 => n3027, B2 => 
                           n3052, ZN => n3029);
   U3761 : AOI22_X1 port map( A1 => n2112, A2 => n3030, B1 => n3029, B2 => 
                           n2101, ZN => n3032);
   U3762 : AOI22_X1 port map( A1 => n2112, A2 => n3039, B1 => n3038, B2 => 
                           n2101, ZN => n3041);
   U3763 : AOI22_X1 port map( A1 => n2112, A2 => n3043, B1 => n3042, B2 => 
                           n2101, ZN => n3045);
   U3764 : MUX2_X1 port map( A => n3045, B => n3044, S => n3055, Z => 
                           DataP_ALU_C_shifter_N59);
   U3765 : INV_X1 port map( A => n3200, ZN => n3049);
   U3766 : INV_X1 port map( A => n3200, ZN => n3050);
   U3767 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_31_port, B1 => 
                           DataP_alu_a_in_30_port, B2 => n3199, ZN => n3060);
   U3768 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_29_port, B1 => 
                           DataP_alu_a_in_28_port, B2 => n3199, ZN => n3062);
   U3769 : AOI22_X1 port map( A1 => n3048, A2 => n3060, B1 => n3062, B2 => 
                           n3047, ZN => n3073);
   U3770 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_27_port, B1 => 
                           DataP_alu_a_in_26_port, B2 => n3199, ZN => n3061);
   U3771 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_25_port, B1 => 
                           DataP_alu_a_in_24_port, B2 => n3199, ZN => n3064);
   U3772 : AOI22_X1 port map( A1 => n3048, A2 => n3061, B1 => n3064, B2 => 
                           n3201, ZN => n3075);
   U3773 : AOI22_X1 port map( A1 => n3202, A2 => n3073, B1 => n3075, B2 => 
                           n3053, ZN => n3126);
   U3774 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_23_port, B1 => 
                           DataP_alu_a_in_22_port, B2 => n3199, ZN => n3063);
   U3775 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_21_port, B1 => 
                           DataP_alu_a_in_20_port, B2 => n3199, ZN => n3066);
   U3776 : AOI22_X1 port map( A1 => n3048, A2 => n3063, B1 => n3066, B2 => 
                           n3047, ZN => n3074);
   U3777 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_19_port, B1 => 
                           DataP_alu_a_in_18_port, B2 => n3199, ZN => n3065);
   U3778 : AOI22_X1 port map( A1 => n2103, A2 => n1751, B1 => 
                           DataP_alu_a_in_16_port, B2 => n3199, ZN => n3068);
   U3779 : AOI22_X1 port map( A1 => n3048, A2 => n3065, B1 => n3068, B2 => 
                           n3047, ZN => n3077);
   U3780 : AOI22_X1 port map( A1 => n3203, A2 => n3074, B1 => n3077, B2 => 
                           n2918, ZN => n3189);
   U3781 : AOI22_X1 port map( A1 => n3205, A2 => n3126, B1 => n3189, B2 => 
                           n2101, ZN => n3101);
   U3782 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_15_port, B1 => 
                           DataP_alu_a_in_14_port, B2 => n3199, ZN => n3067);
   U3783 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_13_port, B1 => 
                           DataP_alu_a_in_12_port, B2 => n3199, ZN => n3070);
   U3784 : AOI22_X1 port map( A1 => n3049, A2 => n3067, B1 => n3070, B2 => 
                           n3201, ZN => n3076);
   U3785 : AOI22_X1 port map( A1 => n2103, A2 => n2200, B1 => 
                           DataP_alu_a_in_10_port, B2 => n2916, ZN => n3069);
   U3786 : AOI22_X1 port map( A1 => n2103, A2 => n2207, B1 => 
                           DataP_alu_a_in_8_port, B2 => n2916, ZN => n3141);
   U3787 : AOI22_X1 port map( A1 => n3048, A2 => n3069, B1 => n3141, B2 => 
                           n3047, ZN => n3162);
   U3788 : AOI22_X1 port map( A1 => n3203, A2 => n3076, B1 => n3162, B2 => 
                           n2918, ZN => n3188);
   U3789 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_7_port, B1 => 
                           DataP_alu_a_in_6_port, B2 => n3199, ZN => n3140);
   U3790 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_5_port, B1 => 
                           DataP_alu_a_in_4_port, B2 => n2916, ZN => n3143);
   U3791 : AOI22_X1 port map( A1 => n3050, A2 => n3140, B1 => n3143, B2 => 
                           n3047, ZN => n3161);
   U3792 : AOI22_X1 port map( A1 => n2103, A2 => n1973, B1 => 
                           DataP_alu_a_in_2_port, B2 => n3199, ZN => n3142);
   U3793 : AOI22_X1 port map( A1 => n2103, A2 => n2232, B1 => n2201, B2 => 
                           n2916, ZN => n3056);
   U3794 : AOI221_X1 port map( B1 => n3142, B2 => n3050, C1 => n3056, C2 => 
                           n3047, A => n3202, ZN => n3057);
   U3795 : AOI21_X1 port map( B1 => n3202, B2 => n3161, A => n3057, ZN => n3058
                           );
   U3796 : AOI22_X1 port map( A1 => n3205, A2 => n3188, B1 => n3058, B2 => 
                           n2101, ZN => n3059);
   U3797 : MUX2_X1 port map( A => n3101, B => n3059, S => n3206, Z => 
                           DataP_ALU_C_shifter_N82);
   U3798 : AOI22_X1 port map( A1 => n3050, A2 => n2073, B1 => n3060, B2 => 
                           n3047, ZN => n3090);
   U3799 : AOI22_X1 port map( A1 => n3048, A2 => n3062, B1 => n3061, B2 => 
                           n3047, ZN => n3092);
   U3800 : AOI22_X1 port map( A1 => n3203, A2 => n3090, B1 => n3092, B2 => 
                           n2918, ZN => n3107);
   U3801 : NAND2_X1 port map( A1 => n3204, A2 => DataP_alu_a_in_31_port, ZN => 
                           n3128);
   U3802 : OAI21_X1 port map( B1 => n3205, B2 => n3107, A => n3128, ZN => n3132
                           );
   U3803 : AOI22_X1 port map( A1 => n3049, A2 => n3064, B1 => n3063, B2 => 
                           n3047, ZN => n3091);
   U3804 : AOI22_X1 port map( A1 => n3049, A2 => n3066, B1 => n3065, B2 => 
                           n3201, ZN => n3094);
   U3805 : AOI22_X1 port map( A1 => n3202, A2 => n3091, B1 => n3094, B2 => 
                           n2918, ZN => n3106);
   U3806 : AOI22_X1 port map( A1 => n3050, A2 => n3068, B1 => n3067, B2 => 
                           n3047, ZN => n3093);
   U3807 : AOI22_X1 port map( A1 => n3048, A2 => n3070, B1 => n3069, B2 => 
                           n3201, ZN => n3176);
   U3808 : AOI22_X1 port map( A1 => n3202, A2 => n3093, B1 => n3176, B2 => 
                           n2918, ZN => n3146);
   U3809 : AOI22_X1 port map( A1 => n3205, A2 => n3106, B1 => n3146, B2 => 
                           n2101, ZN => n3071);
   U3810 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_30_port, B1 => 
                           DataP_alu_a_in_29_port, B2 => n2916, ZN => n3079);
   U3811 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_28_port, B1 => 
                           DataP_alu_a_in_27_port, B2 => n3199, ZN => n3081);
   U3812 : AOI22_X1 port map( A1 => n3050, A2 => n3079, B1 => n3081, B2 => 
                           n3047, ZN => n3097);
   U3813 : NOR2_X1 port map( A1 => n3052, A2 => n2073, ZN => n3089);
   U3814 : AOI21_X1 port map( B1 => n2919, B2 => n3097, A => n3089, ZN => n3109
                           );
   U3815 : OAI21_X1 port map( B1 => n3205, B2 => n3109, A => n3128, ZN => n3134
                           );
   U3816 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_26_port, B1 => 
                           DataP_alu_a_in_25_port, B2 => n2916, ZN => n3080);
   U3817 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_24_port, B1 => 
                           DataP_alu_a_in_23_port, B2 => n3199, ZN => n3083);
   U3818 : AOI22_X1 port map( A1 => n3048, A2 => n3080, B1 => n3083, B2 => 
                           n3047, ZN => n3096);
   U3819 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_22_port, B1 => 
                           DataP_alu_a_in_21_port, B2 => n3199, ZN => n3082);
   U3820 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_20_port, B1 => 
                           DataP_alu_a_in_19_port, B2 => n3199, ZN => n3085);
   U3821 : AOI22_X1 port map( A1 => n3049, A2 => n3082, B1 => n3085, B2 => 
                           n3047, ZN => n3099);
   U3822 : AOI22_X1 port map( A1 => n3202, A2 => n3096, B1 => n3099, B2 => 
                           n2919, ZN => n3108);
   U3823 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_18_port, B1 => 
                           n1751, B2 => n3199, ZN => n3084);
   U3824 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_16_port, B1 => 
                           DataP_alu_a_in_15_port, B2 => n2916, ZN => n3087);
   U3825 : AOI22_X1 port map( A1 => n3050, A2 => n3084, B1 => n3087, B2 => 
                           n3047, ZN => n3098);
   U3826 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_14_port, B1 => 
                           DataP_alu_a_in_13_port, B2 => n3199, ZN => n3086);
   U3827 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_12_port, B1 => 
                           n2200, B2 => n2916, ZN => n3110);
   U3828 : AOI22_X1 port map( A1 => n3048, A2 => n3086, B1 => n3110, B2 => 
                           n3047, ZN => n3183);
   U3829 : AOI22_X1 port map( A1 => n3202, A2 => n3098, B1 => n3183, B2 => 
                           n2919, ZN => n3157);
   U3830 : AOI22_X1 port map( A1 => n3205, A2 => n3108, B1 => n3157, B2 => 
                           n2101, ZN => n3072);
   U3831 : MUX2_X1 port map( A => n3134, B => n3072, S => n3206, Z => 
                           DataP_ALU_C_shifter_N93);
   U3832 : AOI21_X1 port map( B1 => n2919, B2 => n3073, A => n3089, ZN => n3119
                           );
   U3833 : OAI21_X1 port map( B1 => n3205, B2 => n3119, A => n3128, ZN => n3136
                           );
   U3834 : AOI22_X1 port map( A1 => n3202, A2 => n3075, B1 => n3074, B2 => 
                           n2918, ZN => n3118);
   U3835 : AOI22_X1 port map( A1 => n3202, A2 => n3077, B1 => n3076, B2 => 
                           n2918, ZN => n3164);
   U3836 : AOI22_X1 port map( A1 => n3205, A2 => n3118, B1 => n3164, B2 => 
                           n2101, ZN => n3078);
   U3837 : AOI22_X1 port map( A1 => n3050, A2 => n2073, B1 => n3079, B2 => 
                           n3047, ZN => n3103);
   U3838 : AOI21_X1 port map( B1 => n2918, B2 => n3103, A => n3089, ZN => n3121
                           );
   U3839 : OAI21_X1 port map( B1 => n3204, B2 => n3121, A => n3128, ZN => n3138
                           );
   U3840 : AOI22_X1 port map( A1 => n3050, A2 => n3081, B1 => n3080, B2 => 
                           n3047, ZN => n3102);
   U3841 : AOI22_X1 port map( A1 => n3050, A2 => n3083, B1 => n3082, B2 => 
                           n3047, ZN => n3105);
   U3842 : AOI22_X1 port map( A1 => n3202, A2 => n3102, B1 => n3105, B2 => 
                           n3052, ZN => n3120);
   U3843 : AOI22_X1 port map( A1 => n3048, A2 => n3085, B1 => n3084, B2 => 
                           n3047, ZN => n3104);
   U3844 : AOI22_X1 port map( A1 => n3048, A2 => n3087, B1 => n3086, B2 => 
                           n3047, ZN => n3111);
   U3845 : AOI22_X1 port map( A1 => n3202, A2 => n3104, B1 => n3111, B2 => 
                           n3052, ZN => n3171);
   U3846 : AOI22_X1 port map( A1 => n3205, A2 => n3120, B1 => n3171, B2 => 
                           n2101, ZN => n3088);
   U3847 : AOI21_X1 port map( B1 => n3053, B2 => n3090, A => n3089, ZN => n3123
                           );
   U3848 : OAI21_X1 port map( B1 => n3204, B2 => n3123, A => n3128, ZN => n3150
                           );
   U3849 : AOI22_X1 port map( A1 => n3202, A2 => n3092, B1 => n3091, B2 => 
                           n2919, ZN => n3122);
   U3850 : AOI22_X1 port map( A1 => n3202, A2 => n3094, B1 => n3093, B2 => 
                           n2918, ZN => n3178);
   U3851 : AOI22_X1 port map( A1 => n3205, A2 => n3122, B1 => n3178, B2 => 
                           n2101, ZN => n3095);
   U3852 : MUX2_X1 port map( A => n3150, B => n3095, S => n2102, Z => 
                           DataP_ALU_C_shifter_N96);
   U3853 : NAND2_X1 port map( A1 => n3055, A2 => DataP_alu_a_in_31_port, ZN => 
                           n3131);
   U3854 : AOI22_X1 port map( A1 => n3202, A2 => n3097, B1 => n3096, B2 => 
                           n2918, ZN => n3124);
   U3855 : AOI22_X1 port map( A1 => n3202, A2 => n3099, B1 => n3098, B2 => 
                           n3053, ZN => n3185);
   U3856 : AOI221_X1 port map( B1 => n3124, B2 => n3204, C1 => n3185, C2 => 
                           n2101, A => n3055, ZN => n3100);
   U3857 : OR2_X1 port map( A1 => n3195, A2 => n3100, ZN => 
                           DataP_ALU_C_shifter_N97);
   U3858 : AOI22_X1 port map( A1 => n3202, A2 => n3103, B1 => n3102, B2 => 
                           n3052, ZN => n3129);
   U3859 : AOI22_X1 port map( A1 => n3202, A2 => n3105, B1 => n3104, B2 => 
                           n3052, ZN => n3192);
   U3860 : MUX2_X1 port map( A => n3129, B => n3192, S => n2101, Z => n3117);
   U3861 : OAI21_X1 port map( B1 => n3055, B2 => n3117, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N99);
   U3862 : MUX2_X1 port map( A => n3107, B => n3106, S => n2101, Z => n3149);
   U3863 : OAI21_X1 port map( B1 => n3055, B2 => n3149, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N100);
   U3864 : MUX2_X1 port map( A => n3109, B => n3108, S => n2101, Z => n3160);
   U3865 : OAI21_X1 port map( B1 => n3055, B2 => n3160, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N101);
   U3866 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_10_port, B1 => 
                           n2207, B2 => n2916, ZN => n3152);
   U3867 : AOI22_X1 port map( A1 => n3049, A2 => n3110, B1 => n3152, B2 => 
                           n3047, ZN => n3169);
   U3868 : AOI22_X1 port map( A1 => n3202, A2 => n3111, B1 => n3169, B2 => 
                           n2919, ZN => n3191);
   U3869 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_8_port, B1 => 
                           DataP_alu_a_in_7_port, B2 => n3199, ZN => n3151);
   U3870 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_6_port, B1 => 
                           DataP_alu_a_in_5_port, B2 => n3199, ZN => n3154);
   U3871 : AOI22_X1 port map( A1 => n3049, A2 => n3151, B1 => n3154, B2 => 
                           n3047, ZN => n3168);
   U3872 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_4_port, B1 => 
                           n1973, B2 => n3199, ZN => n3153);
   U3873 : AOI22_X1 port map( A1 => n2103, A2 => DataP_alu_a_in_2_port, B1 => 
                           n2232, B2 => n3199, ZN => n3112);
   U3874 : AOI22_X1 port map( A1 => n3048, A2 => n3153, B1 => n3112, B2 => 
                           n3201, ZN => n3113);
   U3875 : AOI22_X1 port map( A1 => n3202, A2 => n3168, B1 => n3113, B2 => 
                           n3052, ZN => n3114);
   U3876 : AOI22_X1 port map( A1 => n3205, A2 => n3191, B1 => n3114, B2 => 
                           n2101, ZN => n3115);
   U3877 : NAND2_X1 port map( A1 => n2102, A2 => n3115, ZN => n3116);
   U3878 : OAI21_X1 port map( B1 => n2102, B2 => n3117, A => n3116, ZN => 
                           DataP_ALU_C_shifter_N83);
   U3879 : MUX2_X1 port map( A => n3119, B => n3118, S => n2101, Z => n3167);
   U3880 : OAI21_X1 port map( B1 => n3055, B2 => n3167, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N102);
   U3881 : MUX2_X1 port map( A => n3121, B => n3120, S => n2101, Z => n3174);
   U3882 : OAI21_X1 port map( B1 => n3055, B2 => n3174, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N103);
   U3883 : MUX2_X1 port map( A => n3123, B => n3122, S => n2101, Z => n3181);
   U3884 : OAI21_X1 port map( B1 => n2138, B2 => n3181, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N104);
   U3885 : OAI21_X1 port map( B1 => n3205, B2 => n3124, A => n3128, ZN => n3125
                           );
   U3886 : OAI21_X1 port map( B1 => n3055, B2 => n3196, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N105);
   U3887 : OAI21_X1 port map( B1 => n3205, B2 => n3126, A => n3128, ZN => n3127
                           );
   U3888 : OAI21_X1 port map( B1 => n3055, B2 => n3197, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N106);
   U3889 : OAI21_X1 port map( B1 => n3205, B2 => n3129, A => n3128, ZN => n3130
                           );
   U3890 : OAI21_X1 port map( B1 => n2138, B2 => n3198, A => n3131, ZN => 
                           DataP_ALU_C_shifter_N107);
   U3891 : AOI21_X1 port map( B1 => n3206, B2 => n3132, A => n3195, ZN => n3133
                           );
   U3892 : AOI21_X1 port map( B1 => n2102, B2 => n3134, A => n3195, ZN => n3135
                           );
   U3893 : AOI21_X1 port map( B1 => n3206, B2 => n3136, A => n3195, ZN => n3137
                           );
   U3894 : AOI21_X1 port map( B1 => n2102, B2 => n3138, A => n3195, ZN => n3139
                           );
   U3895 : AOI22_X1 port map( A1 => n3048, A2 => n3141, B1 => n3140, B2 => 
                           n3047, ZN => n3175);
   U3896 : AOI22_X1 port map( A1 => n3050, A2 => n3143, B1 => n3142, B2 => 
                           n3047, ZN => n3144);
   U3897 : AOI22_X1 port map( A1 => n3202, A2 => n3175, B1 => n3144, B2 => 
                           n2919, ZN => n3145);
   U3898 : AOI22_X1 port map( A1 => n3205, A2 => n3146, B1 => n3145, B2 => 
                           n2101, ZN => n3147);
   U3899 : NAND2_X1 port map( A1 => n2102, A2 => n3147, ZN => n3148);
   U3900 : OAI21_X1 port map( B1 => n3206, B2 => n3149, A => n3148, ZN => 
                           DataP_ALU_C_shifter_N84);
   U3901 : AOI22_X1 port map( A1 => n3048, A2 => n3152, B1 => n3151, B2 => 
                           n3047, ZN => n3182);
   U3902 : AOI22_X1 port map( A1 => n3049, A2 => n3154, B1 => n3153, B2 => 
                           n3047, ZN => n3155);
   U3903 : AOI22_X1 port map( A1 => n3202, A2 => n3182, B1 => n3155, B2 => 
                           n3052, ZN => n3156);
   U3904 : AOI22_X1 port map( A1 => n3205, A2 => n3157, B1 => n3156, B2 => 
                           n2101, ZN => n3158);
   U3905 : NAND2_X1 port map( A1 => n2102, A2 => n3158, ZN => n3159);
   U3906 : AOI22_X1 port map( A1 => n3202, A2 => n3162, B1 => n3161, B2 => 
                           n2919, ZN => n3163);
   U3907 : AOI22_X1 port map( A1 => n3205, A2 => n3164, B1 => n3163, B2 => 
                           n2101, ZN => n3165);
   U3908 : NAND2_X1 port map( A1 => n2102, A2 => n3165, ZN => n3166);
   U3909 : AOI22_X1 port map( A1 => n3202, A2 => n3169, B1 => n3168, B2 => 
                           n2918, ZN => n3170);
   U3910 : AOI22_X1 port map( A1 => n3205, A2 => n3171, B1 => n3170, B2 => 
                           n2101, ZN => n3172);
   U3911 : NAND2_X1 port map( A1 => n2102, A2 => n3172, ZN => n3173);
   U3912 : AOI22_X1 port map( A1 => n3202, A2 => n3176, B1 => n3175, B2 => 
                           n3052, ZN => n3177);
   U3913 : AOI22_X1 port map( A1 => n3205, A2 => n3178, B1 => n3177, B2 => 
                           n2101, ZN => n3179);
   U3914 : NAND2_X1 port map( A1 => n2102, A2 => n3179, ZN => n3180);
   U3915 : AOI22_X1 port map( A1 => n3203, A2 => n3183, B1 => n3182, B2 => 
                           n2918, ZN => n3184);
   U3916 : AOI22_X1 port map( A1 => n3204, A2 => n3185, B1 => n3184, B2 => 
                           n2101, ZN => n3186);
   U3917 : NAND2_X1 port map( A1 => n2102, A2 => n3186, ZN => n3187);
   U3918 : AOI22_X1 port map( A1 => n3205, A2 => n3192, B1 => n3191, B2 => 
                           n2101, ZN => n3193);
   U3919 : NAND2_X1 port map( A1 => n3206, A2 => n3193, ZN => n3194);
   U3920 : INV_X1 port map( A => n3054, ZN => n3204);
   U3921 : INV_X1 port map( A => n2072, ZN => n3209);
   U3922 : MUX2_X1 port map( A => n3247, B => DataP_opcode_M_2_port, S => 
                           DataP_opcode_M_4_port, Z => n3248);
   U3923 : XOR2_X1 port map( A => n1625, B => n524, Z => n3267);
   U3924 : XOR2_X1 port map( A => n1621, B => n523, Z => n3266);
   U3925 : NAND3_X1 port map( A1 => n3268, A2 => n3267, A3 => n3266, ZN => 
                           n3271);
   U3926 : MUX2_X1 port map( A => DataP_opcode_E_0_port, B => 
                           DataP_opcode_E_3_port, S => DataP_opcode_E_1_port, Z
                           => n3280);
   U3927 : MUX2_X1 port map( A => n3282, B => n3281, S => DataP_opcode_E_4_port
                           , Z => n3287);
   U3928 : NAND3_X1 port map( A1 => n3407, A2 => n443, A3 => 
                           ALU_OPCODE_i_3_port, ZN => n3408);
   U3929 : NAND3_X1 port map( A1 => ALU_OPCODE_i_0_port, A2 => 
                           ALU_OPCODE_i_3_port, A3 => n3431, ZN => n3892);
   U3930 : MUX2_X1 port map( A => n3459, B => n3448, S => n2108, Z => n3447);
   U3931 : NAND3_X1 port map( A1 => n2200, A2 => n3886, A3 => n2151, ZN => 
                           n3490);
   U3932 : NAND3_X1 port map( A1 => n3563, A2 => ALU_OPCODE_i_3_port, A3 => 
                           n2395, ZN => n3570);
   U3933 : XOR2_X1 port map( A => n1741, B => n3576, Z => n3582);
   U3934 : XOR2_X1 port map( A => n1740, B => n3587, Z => n3594);
   U3935 : NAND3_X1 port map( A1 => DataP_alu_a_in_15_port, A2 => n3886, A3 => 
                           DataP_alu_b_in_15_port, ZN => n3637);
   U3936 : NAND3_X1 port map( A1 => n3639, A2 => n2371, A3 => n2230, ZN => 
                           n3640);
   U3937 : NAND3_X1 port map( A1 => n3656, A2 => n3655, A3 => n3654, ZN => 
                           n3657);
   U3938 : MUX2_X1 port map( A => n3670, B => n2122, S => n3886, Z => n3671);
   U3939 : NAND3_X1 port map( A1 => n3692, A2 => n2122, A3 => n2124, ZN => 
                           n3693);
   U3940 : MUX2_X1 port map( A => n2120, B => n3723, S => n2108, Z => n3816);
   U3941 : XOR2_X1 port map( A => n3729, B => n1596, Z => n3737);
   U3942 : NAND3_X1 port map( A1 => n3735, A2 => n3734, A3 => n3733, ZN => 
                           n3736);
   U3943 : NAND3_X1 port map( A1 => n3745, A2 => n3744, A3 => n3743, ZN => 
                           n3746);
   U3944 : XOR2_X1 port map( A => n3767, B => n3753, Z => n3761);
   U3945 : NAND3_X1 port map( A1 => n3759, A2 => n3758, A3 => n3757, ZN => 
                           n3760);
   U3946 : NAND3_X1 port map( A1 => n3794, A2 => n3793, A3 => n3792, ZN => 
                           n3795);
   U3947 : NAND3_X1 port map( A1 => n3804, A2 => n3803, A3 => n3802, ZN => 
                           n3805);
   U3948 : NAND3_X1 port map( A1 => n3814, A2 => n3813, A3 => n3812, ZN => 
                           n3815);
   U3949 : MUX2_X1 port map( A => n3839, B => n3856, S => DataP_alu_a_in_8_port
                           , Z => n3842);
   U3950 : NAND3_X1 port map( A1 => DataP_alu_a_in_13_port, A2 => n3890, A3 => 
                           n2141, ZN => n3870);
   U3951 : MUX2_X1 port map( A => n3887, B => n3898, S => n3886, Z => n3889);
   U3952 : NAND3_X1 port map( A1 => n3893, A2 => n3892, A3 => n3891, ZN => 
                           n3895);
   U3953 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_30_port, B1 => 
                           DataP_pc_out_30_port, B2 => n3233, ZN => n3968);
   U3954 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_28_port, B1 => 
                           DataP_pc_out_28_port, B2 => n3233, ZN => n3952);
   U3955 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_26_port, B1 => 
                           DataP_pc_out_26_port, B2 => n3233, ZN => n3953);
   U3956 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_24_port, B1 => 
                           DataP_pc_out_24_port, B2 => n3233, ZN => n3963);
   U3957 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_22_port, B1 => 
                           DataP_pc_out_22_port, B2 => n3233, ZN => n3962);
   U3958 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_20_port, B1 => 
                           DataP_pc_out_20_port, B2 => n3233, ZN => n3959);
   U3959 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_18_port, B1 => 
                           DataP_pc_out_18_port, B2 => n3233, ZN => n3964);
   U3960 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_16_port, B1 => 
                           DataP_pc_out_16_port, B2 => n3233, ZN => n3958);
   U3961 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_14_port, B1 => DataP_pc_out_14_port, 
                           B2 => n3233, ZN => n3957);
   U3962 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_12_port, B1 => DataP_pc_out_12_port, 
                           B2 => n3233, ZN => n3965);
   U3963 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_10_port, B1 => 
                           DataP_pc_out_10_port, B2 => n3233, ZN => n3973);
   U3964 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_8_port, B1 => IRAM_ADDRESS_6_port, B2 
                           => n3233, ZN => n3935);
   U3965 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_6_port, B1 => IRAM_ADDRESS_4_port, B2 
                           => n3233, ZN => n3941);
   U3966 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_4_port, B1 => IRAM_ADDRESS_2_port, B2 
                           => n3233, ZN => n3948);
   U3967 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_2_port, B1 => IRAM_ADDRESS_0_port, B2 
                           => n3233, ZN => DataP_NPC_add_N3);
   U3968 : AOI22_X1 port map( A1 => DataP_npc_mux_sel, A2 => 
                           DataP_npc_pre_3_port, B1 => IRAM_ADDRESS_1_port, B2 
                           => n3233, ZN => n3950);
   U3969 : NOR2_X1 port map( A1 => DataP_NPC_add_N3, A2 => n3950, ZN => n3949);
   U3970 : INV_X1 port map( A => n3949, ZN => n3947);
   U3971 : NOR2_X1 port map( A1 => n3948, A2 => n3947, ZN => n3946);
   U3972 : OAI221_X1 port map( B1 => n2132, B2 => IRAM_ADDRESS_3_port, C1 => 
                           n3233, C2 => DataP_npc_pre_5_port, A => n3946, ZN =>
                           n3942);
   U3973 : NOR2_X1 port map( A1 => n3941, A2 => n3942, ZN => n3940);
   U3974 : OAI221_X1 port map( B1 => n2132, B2 => IRAM_ADDRESS_5_port, C1 => 
                           n3233, C2 => DataP_npc_pre_7_port, A => n3940, ZN =>
                           n3936);
   U3975 : NOR2_X1 port map( A1 => n3935, A2 => n3936, ZN => n3934);
   U3976 : OAI221_X1 port map( B1 => n2132, B2 => IRAM_ADDRESS_7_port, C1 => 
                           n3233, C2 => DataP_npc_pre_9_port, A => n3934, ZN =>
                           n3972);
   U3977 : NOR2_X1 port map( A1 => n3973, A2 => n3972, ZN => n3930);
   U3978 : MUX2_X1 port map( A => DataP_pc_out_11_port, B => 
                           DataP_npc_pre_11_port, S => n2132, Z => n3969);
   U3979 : NAND2_X1 port map( A1 => n3930, A2 => n3969, ZN => n3929);
   U3980 : NOR2_X1 port map( A1 => n3965, A2 => n3929, ZN => n3928);
   U3981 : MUX2_X1 port map( A => DataP_pc_out_13_port, B => 
                           DataP_npc_pre_13_port, S => n2132, Z => n3960);
   U3982 : NAND2_X1 port map( A1 => n3928, A2 => n3960, ZN => n3927);
   U3983 : NOR2_X1 port map( A1 => n3957, A2 => n3927, ZN => n3926);
   U3984 : MUX2_X1 port map( A => DataP_pc_out_15_port, B => 
                           DataP_npc_pre_15_port, S => n2132, Z => n3956);
   U3985 : NAND2_X1 port map( A1 => n3926, A2 => n3956, ZN => n3925);
   U3986 : NOR2_X1 port map( A1 => n3958, A2 => n3925, ZN => n3924);
   U3987 : MUX2_X1 port map( A => DataP_pc_out_17_port, B => 
                           DataP_npc_pre_17_port, S => n2132, Z => n3966);
   U3988 : NAND2_X1 port map( A1 => n3924, A2 => n3966, ZN => n3923);
   U3989 : NOR2_X1 port map( A1 => n3964, A2 => n3923, ZN => n3922);
   U3990 : MUX2_X1 port map( A => DataP_pc_out_19_port, B => 
                           DataP_npc_pre_19_port, S => n2132, Z => n3961);
   U3991 : NAND2_X1 port map( A1 => n3922, A2 => n3961, ZN => n3921);
   U3992 : NOR2_X1 port map( A1 => n3959, A2 => n3921, ZN => n3920);
   U3993 : MUX2_X1 port map( A => DataP_pc_out_21_port, B => 
                           DataP_npc_pre_21_port, S => n2132, Z => n3970);
   U3994 : NAND2_X1 port map( A1 => n3920, A2 => n3970, ZN => n3919);
   U3995 : NOR2_X1 port map( A1 => n3962, A2 => n3919, ZN => n3918);
   U3996 : MUX2_X1 port map( A => DataP_pc_out_23_port, B => 
                           DataP_npc_pre_23_port, S => n2132, Z => n3971);
   U3997 : NAND2_X1 port map( A1 => n3918, A2 => n3971, ZN => n3917);
   U3998 : NOR2_X1 port map( A1 => n3963, A2 => n3917, ZN => n3916);
   U3999 : MUX2_X1 port map( A => DataP_pc_out_25_port, B => 
                           DataP_npc_pre_25_port, S => n2132, Z => n3954);
   U4000 : NAND2_X1 port map( A1 => n3916, A2 => n3954, ZN => n3915);
   U4001 : NOR2_X1 port map( A1 => n3953, A2 => n3915, ZN => n3914);
   U4002 : MUX2_X1 port map( A => DataP_pc_out_27_port, B => 
                           DataP_npc_pre_27_port, S => n2132, Z => n3955);
   U4003 : NAND2_X1 port map( A1 => n3914, A2 => n3955, ZN => n3913);
   U4004 : NOR2_X1 port map( A1 => n3952, A2 => n3913, ZN => n3912);
   U4005 : MUX2_X1 port map( A => DataP_pc_out_29_port, B => 
                           DataP_npc_pre_29_port, S => n2132, Z => n3967);
   U4006 : NAND2_X1 port map( A1 => n3912, A2 => n3967, ZN => n3911);
   U4007 : NOR2_X1 port map( A1 => n3968, A2 => n3911, ZN => n3951);
   U4008 : AOI21_X1 port map( B1 => n3968, B2 => n3911, A => n3951, ZN => 
                           DataP_NPC_add_N31);
   U4009 : XOR2_X1 port map( A => n3912, B => n3967, Z => DataP_NPC_add_N30);
   U4010 : AOI21_X1 port map( B1 => n3952, B2 => n3913, A => n3912, ZN => 
                           DataP_NPC_add_N29);
   U4011 : XOR2_X1 port map( A => n3914, B => n3955, Z => DataP_NPC_add_N28);
   U4012 : AOI21_X1 port map( B1 => n3953, B2 => n3915, A => n3914, ZN => 
                           DataP_NPC_add_N27);
   U4013 : XOR2_X1 port map( A => n3916, B => n3954, Z => DataP_NPC_add_N26);
   U4014 : AOI21_X1 port map( B1 => n3963, B2 => n3917, A => n3916, ZN => 
                           DataP_NPC_add_N25);
   U4015 : XOR2_X1 port map( A => n3918, B => n3971, Z => DataP_NPC_add_N24);
   U4016 : AOI21_X1 port map( B1 => n3962, B2 => n3919, A => n3918, ZN => 
                           DataP_NPC_add_N23);
   U4017 : XOR2_X1 port map( A => n3920, B => n3970, Z => DataP_NPC_add_N22);
   U4018 : AOI21_X1 port map( B1 => n3959, B2 => n3921, A => n3920, ZN => 
                           DataP_NPC_add_N21);
   U4019 : XOR2_X1 port map( A => n3922, B => n3961, Z => DataP_NPC_add_N20);
   U4020 : AOI21_X1 port map( B1 => n3964, B2 => n3923, A => n3922, ZN => 
                           DataP_NPC_add_N19);
   U4021 : XOR2_X1 port map( A => n3924, B => n3966, Z => DataP_NPC_add_N18);
   U4022 : AOI21_X1 port map( B1 => n3958, B2 => n3925, A => n3924, ZN => 
                           DataP_NPC_add_N17);
   U4023 : XOR2_X1 port map( A => n3926, B => n3956, Z => DataP_NPC_add_N16);
   U4024 : AOI21_X1 port map( B1 => n3957, B2 => n3927, A => n3926, ZN => 
                           DataP_NPC_add_N15);
   U4025 : XOR2_X1 port map( A => n3928, B => n3960, Z => DataP_NPC_add_N14);
   U4026 : AOI21_X1 port map( B1 => n3965, B2 => n3929, A => n3928, ZN => 
                           DataP_NPC_add_N13);
   U4027 : XOR2_X1 port map( A => n3930, B => n3969, Z => DataP_NPC_add_N12);
   U4028 : AOI21_X1 port map( B1 => n3973, B2 => n3972, A => n3930, ZN => 
                           DataP_NPC_add_N11);
   U4029 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_9_port, B1 => 
                           IRAM_ADDRESS_7_port, B2 => n3233, ZN => n3933);
   U4030 : INV_X1 port map( A => n3934, ZN => n3932);
   U4031 : INV_X1 port map( A => n3972, ZN => n3931);
   U4032 : AOI21_X1 port map( B1 => n3933, B2 => n3932, A => n3931, ZN => 
                           DataP_NPC_add_N10);
   U4033 : AOI21_X1 port map( B1 => n3935, B2 => n3936, A => n3934, ZN => 
                           DataP_NPC_add_N9);
   U4034 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_7_port, B1 => 
                           IRAM_ADDRESS_5_port, B2 => n3233, ZN => n3939);
   U4035 : INV_X1 port map( A => n3940, ZN => n3938);
   U4036 : INV_X1 port map( A => n3936, ZN => n3937);
   U4037 : AOI21_X1 port map( B1 => n3939, B2 => n3938, A => n3937, ZN => 
                           DataP_NPC_add_N8);
   U4038 : AOI21_X1 port map( B1 => n3941, B2 => n3942, A => n3940, ZN => 
                           DataP_NPC_add_N7);
   U4039 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_5_port, B1 => 
                           IRAM_ADDRESS_3_port, B2 => n3233, ZN => n3945);
   U4040 : INV_X1 port map( A => n3946, ZN => n3944);
   U4041 : INV_X1 port map( A => n3942, ZN => n3943);
   U4042 : AOI21_X1 port map( B1 => n3945, B2 => n3944, A => n3943, ZN => 
                           DataP_NPC_add_N6);
   U4043 : AOI21_X1 port map( B1 => n3948, B2 => n3947, A => n3946, ZN => 
                           DataP_NPC_add_N5);
   U4044 : AOI21_X1 port map( B1 => n3950, B2 => DataP_NPC_add_N3, A => n3949, 
                           ZN => DataP_NPC_add_N4);
   U4045 : AOI22_X1 port map( A1 => n2132, A2 => DataP_npc_pre_31_port, B1 => 
                           DataP_pc_out_31_port, B2 => n3233, ZN => n3974);
   U4046 : XNOR2_X1 port map( A => n3974, B => n3951, ZN => DataP_NPC_add_N32);
   n4224 <= '0';
   n1546 <= '1';
   U4049 : NAND2_X1 port map( A1 => n514, A2 => n515, ZN => n4155);
   U4050 : NAND2_X1 port map( A1 => IR_CU_28, A2 => n516, ZN => n3980);
   U4051 : NOR2_X1 port map( A1 => n4155, A2 => n3980, ZN => n607);
   U4052 : NAND2_X1 port map( A1 => IR_CU_27, A2 => n497, ZN => n4151);
   U4053 : NOR2_X1 port map( A1 => n514, A2 => n515, ZN => n4176);
   U4054 : NAND3_X1 port map( A1 => IR_CU_31, A2 => n4176, A3 => n1960, ZN => 
                           n4012);
   U4055 : NOR2_X1 port map( A1 => IR_CU_27, A2 => n497, ZN => n3996);
   U4056 : INV_X1 port map( A => n4176, ZN => n4177);
   U4057 : NOR2_X1 port map( A1 => n3980, A2 => n4177, ZN => n4013);
   U4058 : NOR3_X1 port map( A1 => IR_CU_27, A2 => n4155, A3 => n516, ZN => 
                           n4046);
   U4059 : AOI22_X1 port map( A1 => IR_CU_31, A2 => n4166, B1 => n2374, B2 => 
                           n504, ZN => n3975);
   U4060 : NAND2_X1 port map( A1 => n515, A2 => n1960, ZN => n4044);
   U4061 : NOR3_X1 port map( A1 => n514, A2 => n2377, A3 => n3980, ZN => n3995)
                           ;
   U4062 : AOI22_X1 port map( A1 => n4055, A2 => n607, B1 => n4052, B2 => n3995
                           , ZN => n3997);
   U4063 : NAND3_X1 port map( A1 => n4166, A2 => n16, A3 => n2377, ZN => n4156)
                           ;
   U4064 : OAI211_X1 port map( C1 => n3975, C2 => n4044, A => n3997, B => n4156
                           , ZN => n3976);
   U4065 : AOI211_X1 port map( C1 => n3996, C2 => n4013, A => n4046, B => n3976
                           , ZN => n3987);
   U4066 : NOR4_X1 port map( A1 => IR_CU_8_port, A2 => IR_CU_6_port, A3 => 
                           IR_CU_7_port, A4 => IR_CU_9_port, ZN => n3977);
   U4067 : NAND3_X1 port map( A1 => n4153, A2 => n484, A3 => n3977, ZN => n3989
                           );
   U4068 : NOR2_X1 port map( A1 => n479, A2 => n3989, ZN => n4023);
   U4069 : NAND2_X1 port map( A1 => IR_CU_5_port, A2 => n4023, ZN => n4001);
   U4070 : NOR3_X1 port map( A1 => n477, A2 => n2375, A3 => n4001, ZN => n3985)
                           ;
   U4071 : NOR3_X1 port map( A1 => n478, A2 => n3989, A3 => n2399, ZN => n4003)
                           ;
   U4072 : NAND2_X1 port map( A1 => n4003, A2 => n476, ZN => n4005);
   U4073 : OAI21_X1 port map( B1 => n476, B2 => n479, A => n2375, ZN => n3978);
   U4074 : OAI211_X1 port map( C1 => n479, C2 => n2375, A => n3978, B => n477, 
                           ZN => n3979);
   U4075 : NAND2_X1 port map( A1 => IR_CU_5_port, A2 => n480, ZN => n4035);
   U4076 : AOI221_X1 port map( B1 => n3989, B2 => n4005, C1 => n3979, C2 => 
                           n4005, A => n4035, ZN => n3984);
   U4077 : INV_X1 port map( A => n3985, ZN => n4032);
   U4078 : NOR3_X1 port map( A1 => n3994, A2 => n4155, A3 => n4151, ZN => n4020
                           );
   U4079 : INV_X1 port map( A => n3980, ZN => n3981);
   U4080 : NAND3_X1 port map( A1 => n514, A2 => n3981, A3 => n2377, ZN => n4016
                           );
   U4081 : NAND4_X1 port map( A1 => n4003, A2 => IR_CU_1_port, A3 => n480, A4 
                           => n482, ZN => n4026);
   U4082 : OAI21_X1 port map( B1 => n504, B2 => n4016, A => n4026, ZN => n4000)
                           ;
   U4083 : AOI211_X1 port map( C1 => n4055, C2 => n3995, A => n4020, B => n4000
                           , ZN => n3983);
   U4084 : NAND3_X1 port map( A1 => n4166, A2 => n4176, A3 => n1960, ZN => 
                           n3982);
   U4085 : OAI211_X1 port map( C1 => n4032, C2 => n476, A => n3983, B => n3982,
                           ZN => n3991);
   U4086 : AOI211_X1 port map( C1 => n3985, C2 => IR_CU_4_port, A => n3984, B 
                           => n3991, ZN => n3986);
   U4087 : OAI211_X1 port map( C1 => n4151, C2 => n4012, A => n3987, B => n3986
                           , ZN => CU_I_aluOpcode_i_0_port);
   U4088 : INV_X1 port map( A => n3994, ZN => n4168);
   U4089 : NAND2_X1 port map( A1 => n4168, A2 => IR_CU_27, ZN => n4154);
   U4090 : NOR2_X1 port map( A1 => IR_CU_1_port, A2 => n478, ZN => n3988);
   U4091 : AOI22_X1 port map( A1 => IR_CU_1_port, A2 => n478, B1 => n3988, B2 
                           => n476, ZN => n4002);
   U4092 : NOR3_X1 port map( A1 => n4002, A2 => n4035, A3 => n3989, ZN => n3990
                           );
   U4093 : AOI21_X1 port map( B1 => n4013, B2 => n4055, A => n3990, ZN => n3993
                           );
   U4094 : NOR3_X1 port map( A1 => IR_CU_1_port, A2 => n478, A3 => n4001, ZN =>
                           n4031);
   U4095 : NOR2_X1 port map( A1 => n516, A2 => n1960, ZN => n4174);
   U4096 : NAND2_X1 port map( A1 => n4176, A2 => n4174, ZN => n4027);
   U4097 : AOI211_X1 port map( C1 => n4031, C2 => n476, A => n3991, B => n4006,
                           ZN => n3992);
   U4098 : OAI211_X1 port map( C1 => n514, C2 => n4154, A => n3993, B => n3992,
                           ZN => CU_I_aluOpcode_i_1_port);
   U4099 : INV_X1 port map( A => n4166, ZN => n4048);
   U4100 : NOR3_X1 port map( A1 => n3994, A2 => n4155, A3 => n4048, ZN => n4019
                           );
   U4101 : NOR3_X1 port map( A1 => n3994, A2 => n4036, A3 => n4177, ZN => n4030
                           );
   U4102 : INV_X1 port map( A => n3995, ZN => n3998);
   U4103 : INV_X1 port map( A => n3996, ZN => n4170);
   U4104 : OAI21_X1 port map( B1 => n3998, B2 => n4170, A => n3997, ZN => n3999
                           );
   U4105 : NOR4_X1 port map( A1 => n4019, A2 => n4030, A3 => n4000, A4 => n3999
                           , ZN => n4011);
   U4106 : NOR3_X1 port map( A1 => n4002, A2 => n4001, A3 => n480, ZN => n4009)
                           ;
   U4107 : NAND3_X1 port map( A1 => n478, A2 => n4023, A3 => n476, ZN => n4034)
                           ;
   U4108 : NAND2_X1 port map( A1 => n4003, A2 => IR_CU_0_port, ZN => n4004);
   U4109 : AOI211_X1 port map( C1 => n4034, C2 => n4004, A => IR_CU_1_port, B 
                           => n4035, ZN => n4008);
   U4110 : NOR3_X1 port map( A1 => IR_CU_4_port, A2 => n477, A3 => n4005, ZN =>
                           n4007);
   U4111 : NOR4_X1 port map( A1 => n4009, A2 => n4008, A3 => n4007, A4 => n4006
                           , ZN => n4010);
   U4112 : OAI211_X1 port map( C1 => n504, C2 => n4012, A => n4011, B => n4010,
                           ZN => CU_I_aluOpcode_i_2_port);
   U4113 : AOI211_X1 port map( C1 => IR_CU_31, C2 => n1960, A => n4177, B => 
                           n4170, ZN => n4018);
   U4114 : NAND2_X1 port map( A1 => n4055, A2 => n4013, ZN => n4015);
   U4115 : NAND2_X1 port map( A1 => n607, A2 => n504, ZN => n4014);
   U4116 : OAI211_X1 port map( C1 => n4048, C2 => n4016, A => n4015, B => n4014
                           , ZN => n4017);
   U4117 : NOR4_X1 port map( A1 => n4020, A2 => n4019, A3 => n4018, A4 => n4017
                           , ZN => n4025);
   U4118 : OAI211_X1 port map( C1 => n2375, C2 => n480, A => IR_CU_5_port, B =>
                           IR_CU_0_port, ZN => n4021);
   U4119 : OAI21_X1 port map( B1 => n478, B2 => n4035, A => n4021, ZN => n4022)
                           ;
   U4120 : NAND3_X1 port map( A1 => n4023, A2 => n477, A3 => n4022, ZN => n4024
                           );
   U4121 : OAI211_X1 port map( C1 => n476, C2 => n4026, A => n4025, B => n4024,
                           ZN => CU_I_aluOpcode_i_3_port);
   U4122 : OAI211_X1 port map( C1 => n516, C2 => n2374, A => n1960, B => n2377,
                           ZN => n4028);
   U4123 : AOI22_X1 port map( A1 => IR_CU_27, A2 => n4028, B1 => n4027, B2 => 
                           n504, ZN => n4029);
   U4124 : AOI211_X1 port map( C1 => n4031, C2 => IR_CU_4_port, A => n4030, B 
                           => n4029, ZN => n4033);
   U4125 : OAI211_X1 port map( C1 => n4035, C2 => n4034, A => n4033, B => n4032
                           , ZN => CU_I_aluOpcode_i_4_port);
   U4126 : OAI211_X1 port map( C1 => IR_CU_26, C2 => n2377, A => IR_CU_28, B =>
                           IR_CU_27, ZN => n4038);
   U4127 : NOR3_X1 port map( A1 => n515, A2 => n1960, A3 => n4036, ZN => n4037)
                           ;
   U4128 : AOI21_X1 port map( B1 => n2374, B2 => n4038, A => n4037, ZN => n4056
                           );
   U4129 : NOR3_X1 port map( A1 => n515, A2 => n2374, A3 => n504, ZN => n4058);
   U4130 : INV_X1 port map( A => n4044, ZN => n4039);
   U4131 : AOI22_X1 port map( A1 => IR_CU_28, A2 => n4058, B1 => n4055, B2 => 
                           n4039, ZN => n4040);
   U4132 : AOI22_X1 port map( A1 => IR_CU_28, A2 => IR_CU_27, B1 => n504, B2 =>
                           n1960, ZN => n4043);
   U4133 : NAND2_X1 port map( A1 => n4176, A2 => n4043, ZN => n4059);
   U4134 : OAI221_X1 port map( B1 => IR_CU_31, B2 => n4056, C1 => IR_CU_31, C2 
                           => n4040, A => n4059, ZN => n4045);
   U4135 : AOI21_X1 port map( B1 => n4168, B2 => n4166, A => n4045, ZN => n1372
                           );
   U4136 : AOI21_X1 port map( B1 => IR_CU_26, B2 => n1960, A => n504, ZN => 
                           n4042);
   U4137 : INV_X1 port map( A => n4155, ZN => n4173);
   U4138 : NAND2_X1 port map( A1 => IR_CU_31, A2 => n4173, ZN => n4041);
   U4139 : OAI21_X1 port map( B1 => n4042, B2 => n4041, A => n1372, ZN => 
                           CU_I_cw_0_port);
   U4140 : AND3_X1 port map( A1 => n4173, A2 => n4043, A3 => n516, ZN => 
                           CU_I_cw_10_port);
   U4141 : AOI21_X1 port map( B1 => n4151, B2 => n4049, A => n4046, ZN => n4061
                           );
   U4142 : INV_X1 port map( A => n4061, ZN => CU_I_cw_6_port);
   U4143 : OR2_X1 port map( A1 => n4045, A2 => CU_I_cw_6_port, ZN => 
                           CU_I_cw_1_port);
   U4144 : NAND2_X1 port map( A1 => n4049, A2 => n2374, ZN => n4051);
   U4145 : AOI22_X1 port map( A1 => n4049, A2 => n4055, B1 => n4046, B2 => 
                           n1960, ZN => n4047);
   U4146 : OAI21_X1 port map( B1 => n4048, B2 => n4051, A => n4047, ZN => 
                           CU_I_cw_3_port);
   U4147 : NAND2_X1 port map( A1 => n4173, A2 => n4174, ZN => n4053);
   U4148 : OAI211_X1 port map( C1 => n2374, C2 => n497, A => n4049, B => n504, 
                           ZN => n4050);
   U4149 : OAI21_X1 port map( B1 => n4170, B2 => n4053, A => n4050, ZN => 
                           CU_I_cw_4_port);
   U4150 : INV_X1 port map( A => n4053, ZN => n4054);
   U4151 : AOI21_X1 port map( B1 => n4055, B2 => n4054, A => CU_I_cw_7_port, ZN
                           => n1358);
   U4152 : INV_X1 port map( A => n4056, ZN => n4057);
   U4153 : AOI221_X1 port map( B1 => n4058, B2 => n516, C1 => n4057, C2 => n516
                           , A => CU_I_cw_10_port, ZN => n4060);
   U4154 : NAND3_X1 port map( A1 => n443, A2 => ALU_OPCODE_i_2_port, A3 => 
                           ALU_OPCODE_i_1_port, ZN => n4101);
   U4155 : NOR4_X1 port map( A1 => DataP_alu_out_W_12_port, A2 => 
                           DataP_alu_out_W_11_port, A3 => 
                           DataP_alu_out_W_10_port, A4 => 
                           DataP_alu_out_W_0_port, ZN => n4065);
   U4156 : NOR4_X1 port map( A1 => DataP_alu_out_W_15_port, A2 => 
                           DataP_alu_out_W_14_port, A3 => 
                           DataP_alu_out_W_13_port, A4 => 
                           DataP_alu_out_W_16_port, ZN => n4064);
   U4157 : NOR4_X1 port map( A1 => DataP_alu_out_W_17_port, A2 => 
                           DataP_alu_out_W_19_port, A3 => 
                           DataP_alu_out_W_18_port, A4 => 
                           DataP_alu_out_W_1_port, ZN => n4063);
   U4158 : NOR4_X1 port map( A1 => DataP_alu_out_W_23_port, A2 => 
                           DataP_alu_out_W_21_port, A3 => 
                           DataP_alu_out_W_20_port, A4 => 
                           DataP_alu_out_W_22_port, ZN => n4062);
   U4159 : NAND4_X1 port map( A1 => n4065, A2 => n4064, A3 => n4063, A4 => 
                           n4062, ZN => n4098);
   U4160 : INV_X1 port map( A => DataP_FWD_MUX_BR_S_0_port, ZN => n4070);
   U4161 : NAND2_X1 port map( A1 => n4070, A2 => DataP_FWD_MUX_BR_S_1_port, ZN 
                           => n4079);
   U4162 : INV_X1 port map( A => n4079, ZN => n4097);
   U4163 : NOR4_X1 port map( A1 => DataP_alu_out_W_27_port, A2 => 
                           DataP_alu_out_W_26_port, A3 => 
                           DataP_alu_out_W_25_port, A4 => 
                           DataP_alu_out_W_24_port, ZN => n4069);
   U4164 : NOR4_X1 port map( A1 => DataP_alu_out_W_30_port, A2 => 
                           DataP_alu_out_W_29_port, A3 => 
                           DataP_alu_out_W_28_port, A4 => 
                           DataP_alu_out_W_2_port, ZN => n4068);
   U4165 : NOR4_X1 port map( A1 => DataP_alu_out_W_31_port, A2 => 
                           DataP_alu_out_W_5_port, A3 => DataP_alu_out_W_4_port
                           , A4 => DataP_alu_out_W_3_port, ZN => n4067);
   U4166 : NOR4_X1 port map( A1 => DataP_alu_out_W_9_port, A2 => 
                           DataP_alu_out_W_8_port, A3 => DataP_alu_out_W_7_port
                           , A4 => DataP_alu_out_W_6_port, ZN => n4066);
   U4167 : NAND4_X1 port map( A1 => n4069, A2 => n4068, A3 => n4067, A4 => 
                           n4066, ZN => n4096);
   U4168 : NOR2_X1 port map( A1 => DataP_FWD_MUX_BR_S_1_port, A2 => n4070, ZN 
                           => n4094);
   U4169 : NOR4_X1 port map( A1 => DataP_A_s_27_port, A2 => DataP_A_s_26_port, 
                           A3 => DataP_A_s_25_port, A4 => DataP_A_s_24_port, ZN
                           => n4074);
   U4170 : NOR4_X1 port map( A1 => DataP_A_s_30_port, A2 => DataP_A_s_29_port, 
                           A3 => DataP_A_s_28_port, A4 => DataP_A_s_2_port, ZN 
                           => n4073);
   U4171 : NOR4_X1 port map( A1 => DataP_A_s_31_port, A2 => DataP_A_s_5_port, 
                           A3 => DataP_A_s_4_port, A4 => DataP_A_s_3_port, ZN 
                           => n4072);
   U4172 : NOR4_X1 port map( A1 => DataP_A_s_9_port, A2 => DataP_A_s_8_port, A3
                           => DataP_A_s_7_port, A4 => DataP_A_s_6_port, ZN => 
                           n4071);
   U4173 : NAND4_X1 port map( A1 => n4074, A2 => n4073, A3 => n4072, A4 => 
                           n4071, ZN => n4081);
   U4174 : NOR4_X1 port map( A1 => DataP_A_s_12_port, A2 => DataP_A_s_11_port, 
                           A3 => DataP_A_s_10_port, A4 => DataP_A_s_0_port, ZN 
                           => n4078);
   U4175 : NOR4_X1 port map( A1 => DataP_A_s_15_port, A2 => DataP_A_s_14_port, 
                           A3 => DataP_A_s_13_port, A4 => DataP_A_s_16_port, ZN
                           => n4077);
   U4176 : NOR4_X1 port map( A1 => DataP_A_s_17_port, A2 => DataP_A_s_19_port, 
                           A3 => DataP_A_s_18_port, A4 => DataP_A_s_1_port, ZN 
                           => n4076);
   U4177 : NOR4_X1 port map( A1 => DataP_A_s_23_port, A2 => DataP_A_s_21_port, 
                           A3 => DataP_A_s_20_port, A4 => DataP_A_s_22_port, ZN
                           => n4075);
   U4178 : NAND4_X1 port map( A1 => n4078, A2 => n4077, A3 => n4076, A4 => 
                           n4075, ZN => n4080);
   U4179 : OAI21_X1 port map( B1 => n4081, B2 => n4080, A => n4079, ZN => n4093
                           );
   U4180 : NOR4_X1 port map( A1 => DRAM_ADDRESS_11_port, A2 => 
                           DRAM_ADDRESS_10_port, A3 => DRAM_ADDRESS_1_port, A4 
                           => DRAM_ADDRESS_0_port, ZN => n4085);
   U4181 : NOR4_X1 port map( A1 => DRAM_ADDRESS_5_port, A2 => 
                           DRAM_ADDRESS_4_port, A3 => DRAM_ADDRESS_3_port, A4 
                           => DRAM_ADDRESS_2_port, ZN => n4084);
   U4182 : NOR4_X1 port map( A1 => DRAM_ADDRESS_9_port, A2 => 
                           DRAM_ADDRESS_8_port, A3 => DRAM_ADDRESS_7_port, A4 
                           => DRAM_ADDRESS_6_port, ZN => n4083);
   U4183 : NOR4_X1 port map( A1 => DataP_alu_out_M_15_port, A2 => 
                           DataP_alu_out_M_14_port, A3 => 
                           DataP_alu_out_M_13_port, A4 => 
                           DataP_alu_out_M_12_port, ZN => n4082);
   U4184 : NAND4_X1 port map( A1 => n4085, A2 => n4084, A3 => n4083, A4 => 
                           n4082, ZN => n4091);
   U4185 : NOR4_X1 port map( A1 => DataP_alu_out_M_16_port, A2 => 
                           DataP_alu_out_M_17_port, A3 => 
                           DataP_alu_out_M_19_port, A4 => 
                           DataP_alu_out_M_18_port, ZN => n4089);
   U4186 : NOR4_X1 port map( A1 => DataP_alu_out_M_23_port, A2 => 
                           DataP_alu_out_M_21_port, A3 => 
                           DataP_alu_out_M_20_port, A4 => 
                           DataP_alu_out_M_22_port, ZN => n4088);
   U4187 : NOR4_X1 port map( A1 => DataP_alu_out_M_27_port, A2 => 
                           DataP_alu_out_M_26_port, A3 => 
                           DataP_alu_out_M_25_port, A4 => 
                           DataP_alu_out_M_24_port, ZN => n4087);
   U4188 : NOR4_X1 port map( A1 => DataP_alu_out_M_31_port, A2 => 
                           DataP_alu_out_M_30_port, A3 => 
                           DataP_alu_out_M_29_port, A4 => 
                           DataP_alu_out_M_28_port, ZN => n4086);
   U4189 : NAND4_X1 port map( A1 => n4089, A2 => n4088, A3 => n4087, A4 => 
                           n4086, ZN => n4090);
   U4190 : OAI21_X1 port map( B1 => n4091, B2 => n4090, A => n4094, ZN => n4092
                           );
   U4191 : OAI21_X1 port map( B1 => n4094, B2 => n4093, A => n4092, ZN => n4095
                           );
   U4192 : AOI221_X1 port map( B1 => n4098, B2 => n4097, C1 => n4096, C2 => 
                           n4097, A => n4095, ZN => n4099);
   U4193 : XNOR2_X1 port map( A => DataP_pr_E, B => n4099, ZN => n4183);
   U4194 : NAND2_X1 port map( A1 => BR_EN_i, A2 => ALU_OPCODE_i_3_port, ZN => 
                           n4182);
   U4195 : NAND2_X1 port map( A1 => ALU_OPCODE_i_1_port, A2 => 
                           ALU_OPCODE_i_0_port, ZN => n4100);
   U4196 : INV_X1 port map( A => DataP_npc_8_port, ZN => n4214);
   U4197 : INV_X1 port map( A => DataP_npc_9_port, ZN => n4213);
   U4198 : OAI22_X1 port map( A1 => n341, A2 => n4111, B1 => n4110, B2 => n4213
                           , ZN => DataP_PC_reg_N11);
   U4199 : INV_X1 port map( A => DataP_npc_10_port, ZN => n4212);
   U4200 : OAI22_X1 port map( A1 => n340, A2 => n4111, B1 => n4110, B2 => n4212
                           , ZN => DataP_PC_reg_N12);
   U4201 : INV_X1 port map( A => DataP_npc_11_port, ZN => n4211);
   U4202 : OAI22_X1 port map( A1 => n2386, A2 => n4111, B1 => n4110, B2 => 
                           n4211, ZN => DataP_PC_reg_N13);
   U4203 : INV_X1 port map( A => DataP_npc_12_port, ZN => n4210);
   U4204 : OAI22_X1 port map( A1 => n337, A2 => n4111, B1 => n4110, B2 => n4210
                           , ZN => DataP_PC_reg_N14);
   U4205 : NAND3_X1 port map( A1 => n2434, A2 => n4107, A3 => n4106, ZN => 
                           n4105);
   U4206 : INV_X1 port map( A => DataP_npc_0_port, ZN => n4223);
   U4207 : OAI22_X1 port map( A1 => n296, A2 => n4111, B1 => n4110, B2 => n4223
                           , ZN => DataP_PC_reg_N2);
   U4208 : INV_X1 port map( A => DataP_npc_1_port, ZN => n4221);
   U4209 : OAI22_X1 port map( A1 => n358, A2 => n4111, B1 => n4110, B2 => n4221
                           , ZN => DataP_PC_reg_N3);
   U4210 : INV_X1 port map( A => DataP_npc_2_port, ZN => n4220);
   U4211 : OAI22_X1 port map( A1 => n357, A2 => n4111, B1 => n4110, B2 => n4220
                           , ZN => DataP_PC_reg_N4);
   U4212 : INV_X1 port map( A => DataP_npc_3_port, ZN => n4219);
   U4213 : INV_X1 port map( A => DataP_npc_4_port, ZN => n4218);
   U4214 : INV_X1 port map( A => DataP_npc_5_port, ZN => n4217);
   U4215 : OAI22_X1 port map( A1 => n354, A2 => n4111, B1 => n4110, B2 => n4217
                           , ZN => DataP_PC_reg_N7);
   U4216 : INV_X1 port map( A => DataP_npc_6_port, ZN => n4216);
   U4217 : INV_X1 port map( A => DataP_npc_7_port, ZN => n4215);
   U4218 : OAI22_X1 port map( A1 => n350, A2 => n4111, B1 => n4110, B2 => n4215
                           , ZN => DataP_PC_reg_N9);
   U4219 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_0_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_0_port, ZN => n4112);
   U4220 : OAI21_X1 port map( B1 => n2521, B2 => n4146, A => n4112, ZN => 
                           DataP_WB_0_port);
   U4221 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_10_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_10_port, ZN => n4113)
                           ;
   U4222 : OAI21_X1 port map( B1 => n2503, B2 => n4146, A => n4113, ZN => 
                           DataP_WB_10_port);
   U4223 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_11_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_11_port, ZN => n4114)
                           ;
   U4224 : OAI21_X1 port map( B1 => n2518, B2 => n4146, A => n4114, ZN => 
                           DataP_WB_11_port);
   U4225 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_12_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_12_port, ZN => n4115)
                           ;
   U4226 : OAI21_X1 port map( B1 => n2492, B2 => n4146, A => n4115, ZN => 
                           DataP_WB_12_port);
   U4227 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_13_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_13_port, ZN => n4116)
                           ;
   U4228 : OAI21_X1 port map( B1 => n2504, B2 => n4146, A => n4116, ZN => 
                           DataP_WB_13_port);
   U4229 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_14_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_14_port, ZN => n4117)
                           ;
   U4230 : OAI21_X1 port map( B1 => n2497, B2 => n4146, A => n4117, ZN => 
                           DataP_WB_14_port);
   U4231 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_15_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_15_port, ZN => n4118)
                           ;
   U4232 : OAI21_X1 port map( B1 => n2516, B2 => n4146, A => n4118, ZN => 
                           DataP_WB_15_port);
   U4233 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_16_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_16_port, ZN => n4119)
                           ;
   U4234 : OAI21_X1 port map( B1 => n2511, B2 => n4146, A => n4119, ZN => 
                           DataP_WB_16_port);
   U4235 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_17_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_17_port, ZN => n4120)
                           ;
   U4236 : OAI21_X1 port map( B1 => n2493, B2 => n4146, A => n4120, ZN => 
                           DataP_WB_17_port);
   U4237 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_18_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_18_port, ZN => n4121)
                           ;
   U4238 : OAI21_X1 port map( B1 => n2505, B2 => n4146, A => n4121, ZN => 
                           DataP_WB_18_port);
   U4239 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_19_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_19_port, ZN => n4122)
                           ;
   U4240 : OAI21_X1 port map( B1 => n2498, B2 => n4146, A => n4122, ZN => 
                           DataP_WB_19_port);
   U4241 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_1_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_1_port, ZN => n4123);
   U4242 : OAI21_X1 port map( B1 => n2522, B2 => n4146, A => n4123, ZN => 
                           DataP_WB_1_port);
   U4243 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_20_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_20_port, ZN => n4124)
                           ;
   U4244 : OAI21_X1 port map( B1 => n2506, B2 => n4146, A => n4124, ZN => 
                           DataP_WB_20_port);
   U4245 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_21_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_21_port, ZN => n4125)
                           ;
   U4246 : OAI21_X1 port map( B1 => n2499, B2 => n4146, A => n4125, ZN => 
                           DataP_WB_21_port);
   U4247 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_22_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_22_port, ZN => n4126)
                           ;
   U4248 : OAI21_X1 port map( B1 => n2512, B2 => n4146, A => n4126, ZN => 
                           DataP_WB_22_port);
   U4249 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_23_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_23_port, ZN => n4127)
                           ;
   U4250 : OAI21_X1 port map( B1 => n2494, B2 => n4146, A => n4127, ZN => 
                           DataP_WB_23_port);
   U4251 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_24_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_24_port, ZN => n4128)
                           ;
   U4252 : OAI21_X1 port map( B1 => n2513, B2 => n4146, A => n4128, ZN => 
                           DataP_WB_24_port);
   U4253 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_25_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_25_port, ZN => n4129)
                           ;
   U4254 : OAI21_X1 port map( B1 => n2507, B2 => n4146, A => n4129, ZN => 
                           DataP_WB_25_port);
   U4255 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_26_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_26_port, ZN => n4130)
                           ;
   U4256 : OAI21_X1 port map( B1 => n2500, B2 => n4146, A => n4130, ZN => 
                           DataP_WB_26_port);
   U4257 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_27_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_27_port, ZN => n4131)
                           ;
   U4258 : OAI21_X1 port map( B1 => n2495, B2 => n4146, A => n4131, ZN => 
                           DataP_WB_27_port);
   U4259 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_28_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_28_port, ZN => n4132)
                           ;
   U4260 : OAI21_X1 port map( B1 => n2508, B2 => n4146, A => n4132, ZN => 
                           DataP_WB_28_port);
   U4261 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_29_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_29_port, ZN => n4133)
                           ;
   U4262 : OAI21_X1 port map( B1 => n2501, B2 => n4146, A => n4133, ZN => 
                           DataP_WB_29_port);
   U4263 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_2_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_2_port, ZN => n4134);
   U4264 : OAI21_X1 port map( B1 => n2514, B2 => n4146, A => n4134, ZN => 
                           DataP_WB_2_port);
   U4265 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_30_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_30_port, ZN => n4135)
                           ;
   U4266 : OAI21_X1 port map( B1 => n2496, B2 => n4146, A => n4135, ZN => 
                           DataP_WB_30_port);
   U4267 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_31_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_31_port, ZN => n4136)
                           ;
   U4268 : OAI21_X1 port map( B1 => n2517, B2 => n4146, A => n4136, ZN => 
                           DataP_WB_31_port);
   U4269 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_3_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_3_port, ZN => n4137);
   U4270 : OAI21_X1 port map( B1 => n2523, B2 => n4146, A => n4137, ZN => 
                           DataP_WB_3_port);
   U4271 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_4_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_4_port, ZN => n4138);
   U4272 : OAI21_X1 port map( B1 => n2509, B2 => n4146, A => n4138, ZN => 
                           DataP_WB_4_port);
   U4273 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_5_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_5_port, ZN => n4139);
   U4274 : OAI21_X1 port map( B1 => n2520, B2 => n4146, A => n4139, ZN => 
                           DataP_WB_5_port);
   U4275 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_6_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_6_port, ZN => n4140);
   U4276 : OAI21_X1 port map( B1 => n2515, B2 => n4146, A => n4140, ZN => 
                           DataP_WB_6_port);
   U4277 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_7_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_7_port, ZN => n4141);
   U4278 : OAI21_X1 port map( B1 => n2510, B2 => n4146, A => n4141, ZN => 
                           DataP_WB_7_port);
   U4279 : AOI22_X1 port map( A1 => n4144, A2 => DataP_LMD_out_8_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_8_port, ZN => n4142);
   U4280 : OAI21_X1 port map( B1 => n2502, B2 => n4146, A => n4142, ZN => 
                           DataP_WB_8_port);
   U4281 : AOI22_X1 port map( A1 => n3229, A2 => DataP_LMD_out_9_port, B1 => 
                           n4143, B2 => DataP_link_addr_W_9_port, ZN => n4145);
   U4282 : OAI21_X1 port map( B1 => n2519, B2 => n4146, A => n4145, ZN => 
                           DataP_WB_9_port);
   U4283 : INV_X1 port map( A => n16, ZN => n4152);
   U4284 : AOI211_X1 port map( C1 => n607, C2 => n504, A => CU_I_cw_7_port, B 
                           => n4153, ZN => n4150);
   U4285 : OAI211_X1 port map( C1 => n4152, C2 => n4151, A => Rst, B => n4150, 
                           ZN => n4164);
   U4286 : AND2_X1 port map( A1 => Rst, A2 => n4153, ZN => n4162);
   U4287 : NOR2_X1 port map( A1 => n4155, A2 => n4154, ZN => n4165);
   U4288 : NAND2_X1 port map( A1 => Rst, A2 => n4165, ZN => n4179);
   U4289 : OAI22_X1 port map( A1 => n497, A2 => n4179, B1 => n4156, B2 => n4164
                           , ZN => n4161);
   U4290 : AOI21_X1 port map( B1 => n4162, B2 => DataP_IR1_11_port, A => n4161,
                           ZN => n4157);
   U4291 : OAI21_X1 port map( B1 => n485, B2 => n4164, A => n4157, ZN => 
                           DataP_dest_D_0_port);
   U4292 : AOI21_X1 port map( B1 => n4162, B2 => DataP_IR1_12_port, A => n4161,
                           ZN => n4158);
   U4293 : OAI21_X1 port map( B1 => n486, B2 => n4164, A => n4158, ZN => 
                           DataP_dest_D_1_port);
   U4294 : AOI21_X1 port map( B1 => n4162, B2 => DataP_IR1_13_port, A => n4161,
                           ZN => n4159);
   U4295 : OAI21_X1 port map( B1 => n487, B2 => n4164, A => n4159, ZN => 
                           DataP_dest_D_2_port);
   U4296 : AOI21_X1 port map( B1 => n4162, B2 => DataP_IR1_14_port, A => n4161,
                           ZN => n4160);
   U4297 : OAI21_X1 port map( B1 => n488, B2 => n4164, A => n4160, ZN => 
                           DataP_dest_D_3_port);
   U4298 : AOI21_X1 port map( B1 => n4162, B2 => DataP_IR1_15_port, A => n4161,
                           ZN => n4163);
   U4299 : OAI21_X1 port map( B1 => n489, B2 => n4164, A => n4163, ZN => 
                           DataP_dest_D_4_port);
   U4300 : NAND2_X1 port map( A1 => IR_CU_28, A2 => n4166, ZN => n4171);
   U4301 : OAI21_X1 port map( B1 => n515, B2 => IR_CU_27, A => n2374, ZN => 
                           n4167);
   U4302 : AOI22_X1 port map( A1 => n4168, A2 => n497, B1 => n1960, B2 => n4167
                           , ZN => n4169);
   U4303 : OAI221_X1 port map( B1 => n514, B2 => n4171, C1 => n2374, C2 => 
                           n4170, A => n4169, ZN => n4172);
   U4304 : AOI211_X1 port map( C1 => IR_CU_27, C2 => n4174, A => n4173, B => 
                           n4172, ZN => n4175);
   U4305 : OAI221_X1 port map( B1 => IR_CU_31, B2 => n4177, C1 => n516, C2 => 
                           n4176, A => n4175, ZN => n4178);
   U4306 : NAND4_X1 port map( A1 => Rst, A2 => DataP_IR1_15_port, A3 => n4181, 
                           A4 => n4178, ZN => n4180);
   U4307 : OAI21_X1 port map( B1 => n485, B2 => n4179, A => n4180, ZN => 
                           DataP_imm_out_16_port);
   U4308 : OAI21_X1 port map( B1 => n486, B2 => n4179, A => n4180, ZN => 
                           DataP_imm_out_17_port);
   U4309 : OAI21_X1 port map( B1 => n487, B2 => n4179, A => n4180, ZN => 
                           DataP_imm_out_18_port);
   U4310 : OAI21_X1 port map( B1 => n488, B2 => n4179, A => n4180, ZN => 
                           DataP_imm_out_19_port);
   U4311 : OAI21_X1 port map( B1 => n489, B2 => n4179, A => n4180, ZN => 
                           DataP_imm_out_20_port);
   U4312 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_21_port, ZN => n4189);
   U4313 : OAI21_X1 port map( B1 => n4181, B2 => n4189, A => n4180, ZN => 
                           DataP_imm_out_21_port);
   U4314 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_22_port, ZN => n4188);
   U4315 : OAI21_X1 port map( B1 => n4181, B2 => n4188, A => n4180, ZN => 
                           DataP_imm_out_22_port);
   U4316 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_23_port, ZN => n4187);
   U4317 : OAI21_X1 port map( B1 => n4181, B2 => n4187, A => n4180, ZN => 
                           DataP_imm_out_23_port);
   U4318 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_24_port, ZN => n4186);
   U4319 : OAI21_X1 port map( B1 => n4181, B2 => n4186, A => n4180, ZN => 
                           DataP_imm_out_24_port);
   U4320 : NAND2_X1 port map( A1 => Rst, A2 => DataP_IR1_25_port, ZN => n4185);
   U4321 : OAI21_X1 port map( B1 => n4181, B2 => n4185, A => n4180, ZN => 
                           DataP_imm_out_31_port);
   U4322 : MUX2_X1 port map( A => DataP_pc_out_0, B => DataP_npc_pre_0_port, S 
                           => n2132, Z => DataP_NPC_add_N1);
   U4323 : MUX2_X1 port map( A => DataP_pc_out_1, B => DataP_npc_pre_1_port, S 
                           => n2132, Z => DataP_NPC_add_N2);
   U4324 : MUX2_X1 port map( A => DataP_link_addr_D_31_port, B => 
                           DataP_link_addr_F_31_port, S => n3230, Z => n1481);
   U4325 : MUX2_X1 port map( A => DataP_link_addr_D_0_port, B => 
                           DataP_link_addr_F_0_port, S => n3230, Z => n1480);
   U4326 : MUX2_X1 port map( A => DataP_link_addr_D_1_port, B => 
                           DataP_link_addr_F_1_port, S => n3230, Z => n1479);
   U4327 : MUX2_X1 port map( A => DataP_link_addr_D_2_port, B => 
                           DataP_link_addr_F_2_port, S => n3230, Z => n1478);
   U4328 : MUX2_X1 port map( A => DataP_link_addr_D_3_port, B => 
                           DataP_link_addr_F_3_port, S => n3230, Z => n1477);
   U4329 : MUX2_X1 port map( A => DataP_link_addr_D_4_port, B => 
                           DataP_link_addr_F_4_port, S => n3230, Z => n1476);
   U4330 : MUX2_X1 port map( A => DataP_link_addr_D_5_port, B => 
                           DataP_link_addr_F_5_port, S => n3230, Z => n1475);
   U4331 : MUX2_X1 port map( A => DataP_link_addr_D_6_port, B => 
                           DataP_link_addr_F_6_port, S => n3230, Z => n1474);
   U4332 : MUX2_X1 port map( A => DataP_link_addr_D_7_port, B => 
                           DataP_link_addr_F_7_port, S => n3230, Z => n1473);
   U4333 : MUX2_X1 port map( A => DataP_link_addr_D_8_port, B => 
                           DataP_link_addr_F_8_port, S => n3230, Z => n1472);
   U4334 : MUX2_X1 port map( A => DataP_link_addr_D_9_port, B => 
                           DataP_link_addr_F_9_port, S => n3230, Z => n1471);
   U4335 : MUX2_X1 port map( A => DataP_link_addr_D_10_port, B => 
                           DataP_link_addr_F_10_port, S => n3230, Z => n1470);
   U4336 : MUX2_X1 port map( A => DataP_link_addr_D_11_port, B => 
                           DataP_link_addr_F_11_port, S => n3231, Z => n1469);
   U4337 : MUX2_X1 port map( A => DataP_link_addr_D_12_port, B => 
                           DataP_link_addr_F_12_port, S => n3231, Z => n1468);
   U4338 : MUX2_X1 port map( A => DataP_link_addr_D_13_port, B => 
                           DataP_link_addr_F_13_port, S => n3231, Z => n1467);
   U4339 : MUX2_X1 port map( A => DataP_link_addr_D_14_port, B => 
                           DataP_link_addr_F_14_port, S => n3231, Z => n1466);
   U4340 : MUX2_X1 port map( A => DataP_link_addr_D_15_port, B => 
                           DataP_link_addr_F_15_port, S => n3231, Z => n1465);
   U4341 : MUX2_X1 port map( A => DataP_link_addr_D_16_port, B => 
                           DataP_link_addr_F_16_port, S => n3231, Z => n1464);
   U4342 : MUX2_X1 port map( A => DataP_link_addr_D_17_port, B => 
                           DataP_link_addr_F_17_port, S => n3231, Z => n1463);
   U4343 : MUX2_X1 port map( A => DataP_link_addr_D_18_port, B => 
                           DataP_link_addr_F_18_port, S => n3231, Z => n1462);
   U4344 : MUX2_X1 port map( A => DataP_link_addr_D_19_port, B => 
                           DataP_link_addr_F_19_port, S => n3231, Z => n1461);
   U4345 : MUX2_X1 port map( A => DataP_link_addr_D_20_port, B => 
                           DataP_link_addr_F_20_port, S => n3231, Z => n1460);
   U4346 : MUX2_X1 port map( A => DataP_link_addr_D_21_port, B => 
                           DataP_link_addr_F_21_port, S => n3231, Z => n1459);
   U4347 : MUX2_X1 port map( A => DataP_link_addr_D_22_port, B => 
                           DataP_link_addr_F_22_port, S => n3231, Z => n1458);
   U4348 : MUX2_X1 port map( A => DataP_link_addr_D_23_port, B => 
                           DataP_link_addr_F_23_port, S => n3230, Z => n1457);
   U4349 : MUX2_X1 port map( A => DataP_link_addr_D_24_port, B => 
                           DataP_link_addr_F_24_port, S => n3231, Z => n1456);
   U4350 : MUX2_X1 port map( A => DataP_link_addr_D_25_port, B => 
                           DataP_link_addr_F_25_port, S => n3230, Z => n1455);
   U4351 : MUX2_X1 port map( A => DataP_link_addr_D_26_port, B => 
                           DataP_link_addr_F_26_port, S => n3231, Z => n1454);
   U4352 : MUX2_X1 port map( A => DataP_link_addr_D_27_port, B => 
                           DataP_link_addr_F_27_port, S => n3230, Z => n1453);
   U4353 : MUX2_X1 port map( A => DataP_link_addr_D_28_port, B => 
                           DataP_link_addr_F_28_port, S => n3231, Z => n1452);
   U4354 : MUX2_X1 port map( A => DataP_link_addr_D_29_port, B => 
                           DataP_link_addr_F_29_port, S => n3230, Z => n1451);
   U4355 : MUX2_X1 port map( A => DataP_link_addr_D_30_port, B => 
                           DataP_link_addr_F_30_port, S => n3231, Z => n1450);
   U4356 : MUX2_X1 port map( A => DataP_pr_D, B => DataP_prediction, S => n3230
                           , Z => n1449);
   U4357 : NAND2_X1 port map( A1 => DataP_npc_31_port, A2 => n3232, ZN => n163)
                           ;
   U4358 : AOI21_X1 port map( B1 => n4191, B2 => n2104, A => n3235, ZN => n162)
                           ;
   U4359 : NAND2_X1 port map( A1 => DataP_npc_30_port, A2 => n3232, ZN => n159)
                           ;
   U4360 : AOI21_X1 port map( B1 => n4192, B2 => n2104, A => n3235, ZN => n158)
                           ;
   U4361 : NAND2_X1 port map( A1 => DataP_npc_29_port, A2 => n3232, ZN => n155)
                           ;
   U4362 : AOI21_X1 port map( B1 => n4193, B2 => n2104, A => n3235, ZN => n154)
                           ;
   U4363 : NAND2_X1 port map( A1 => DataP_npc_28_port, A2 => n3232, ZN => n151)
                           ;
   U4364 : AOI21_X1 port map( B1 => n4194, B2 => n2104, A => n3235, ZN => n150)
                           ;
   U4365 : NAND2_X1 port map( A1 => DataP_npc_27_port, A2 => n3232, ZN => n147)
                           ;
   U4366 : AOI21_X1 port map( B1 => n4195, B2 => n2104, A => n3235, ZN => n146)
                           ;
   U4367 : NAND2_X1 port map( A1 => DataP_npc_26_port, A2 => n3232, ZN => n143)
                           ;
   U4368 : AOI21_X1 port map( B1 => n4196, B2 => n2104, A => n3235, ZN => n142)
                           ;
   U4369 : NAND2_X1 port map( A1 => DataP_npc_25_port, A2 => n3232, ZN => n139)
                           ;
   U4370 : AOI21_X1 port map( B1 => n4197, B2 => n2104, A => n3235, ZN => n138)
                           ;
   U4371 : NAND2_X1 port map( A1 => DataP_npc_24_port, A2 => n3232, ZN => n135)
                           ;
   U4372 : AOI21_X1 port map( B1 => n4198, B2 => n2104, A => n3235, ZN => n134)
                           ;
   U4373 : NAND2_X1 port map( A1 => DataP_npc_23_port, A2 => n3232, ZN => n131)
                           ;
   U4374 : AOI21_X1 port map( B1 => n4199, B2 => n2104, A => n3235, ZN => n130)
                           ;
   U4375 : NAND2_X1 port map( A1 => DataP_npc_22_port, A2 => n3232, ZN => n127)
                           ;
   U4376 : AOI21_X1 port map( B1 => n4200, B2 => n2104, A => n3235, ZN => n126)
                           ;
   U4377 : NAND2_X1 port map( A1 => DataP_npc_21_port, A2 => n4222, ZN => n123)
                           ;
   U4378 : AOI21_X1 port map( B1 => n4201, B2 => n2104, A => n3235, ZN => n122)
                           ;
   U4379 : NAND2_X1 port map( A1 => DataP_npc_20_port, A2 => n4222, ZN => n119)
                           ;
   U4380 : AOI21_X1 port map( B1 => n4202, B2 => n2104, A => n3236, ZN => n118)
                           ;
   U4381 : NAND2_X1 port map( A1 => DataP_npc_19_port, A2 => n4222, ZN => n115)
                           ;
   U4382 : AOI21_X1 port map( B1 => n4203, B2 => n2104, A => n3235, ZN => n114)
                           ;
   U4383 : NAND2_X1 port map( A1 => DataP_npc_18_port, A2 => n3232, ZN => n111)
                           ;
   U4384 : AOI21_X1 port map( B1 => n4204, B2 => n2104, A => n3235, ZN => n110)
                           ;
   U4385 : NAND2_X1 port map( A1 => DataP_npc_17_port, A2 => n4222, ZN => n107)
                           ;
   U4386 : AOI21_X1 port map( B1 => n4205, B2 => n2104, A => n3235, ZN => n106)
                           ;
   U4387 : NAND2_X1 port map( A1 => DataP_npc_16_port, A2 => n3232, ZN => n103)
                           ;
   U4388 : AOI21_X1 port map( B1 => n4206, B2 => n2104, A => n3236, ZN => n102)
                           ;
   U4389 : NAND2_X1 port map( A1 => DataP_npc_15_port, A2 => n4222, ZN => n99);
   U4390 : AOI21_X1 port map( B1 => n4207, B2 => n2104, A => n3236, ZN => n98);
   U4391 : NAND2_X1 port map( A1 => DataP_npc_14_port, A2 => n3232, ZN => n95);
   U4392 : AOI21_X1 port map( B1 => n4208, B2 => n2104, A => n3236, ZN => n94);
   U4393 : NAND2_X1 port map( A1 => DataP_npc_13_port, A2 => n4222, ZN => n91);
   U4394 : AOI21_X1 port map( B1 => n4209, B2 => n2104, A => n3236, ZN => n90);
   U4395 : NAND2_X1 port map( A1 => DataP_npc_12_port, A2 => n4222, ZN => n87);
   U4396 : AOI21_X1 port map( B1 => n4210, B2 => n2104, A => n3236, ZN => n86);
   U4397 : NAND2_X1 port map( A1 => DataP_npc_11_port, A2 => n4222, ZN => n83);
   U4398 : AOI21_X1 port map( B1 => n4211, B2 => n2104, A => n3236, ZN => n82);
   U4399 : NAND2_X1 port map( A1 => DataP_npc_10_port, A2 => n4222, ZN => n79);
   U4400 : AOI21_X1 port map( B1 => n4212, B2 => n2104, A => n3236, ZN => n78);
   U4401 : NAND2_X1 port map( A1 => DataP_npc_9_port, A2 => n4222, ZN => n75);
   U4402 : AOI21_X1 port map( B1 => n4213, B2 => n2104, A => n3236, ZN => n74);
   U4403 : NAND2_X1 port map( A1 => DataP_npc_8_port, A2 => n4222, ZN => n71);
   U4404 : AOI21_X1 port map( B1 => n4214, B2 => n2104, A => n3236, ZN => n70);
   U4405 : NAND2_X1 port map( A1 => DataP_npc_7_port, A2 => n3232, ZN => n67);
   U4406 : AOI21_X1 port map( B1 => n4215, B2 => n2104, A => n3236, ZN => n66);
   U4407 : NAND2_X1 port map( A1 => DataP_npc_6_port, A2 => n3232, ZN => n63);
   U4408 : AOI21_X1 port map( B1 => n4216, B2 => n2104, A => n3236, ZN => n62);
   U4409 : NAND2_X1 port map( A1 => DataP_npc_5_port, A2 => n3232, ZN => n59);
   U4410 : AOI21_X1 port map( B1 => n4217, B2 => n2104, A => n3236, ZN => n58);
   U4411 : NAND2_X1 port map( A1 => DataP_npc_4_port, A2 => n3232, ZN => n55);
   U4412 : AOI21_X1 port map( B1 => n4218, B2 => n2104, A => n3236, ZN => n54);
   U4413 : NAND2_X1 port map( A1 => DataP_npc_3_port, A2 => n3232, ZN => n51);
   U4414 : AOI21_X1 port map( B1 => n4219, B2 => n2104, A => n3236, ZN => n50);
   U4415 : NAND2_X1 port map( A1 => DataP_npc_2_port, A2 => n3232, ZN => n47);
   U4416 : AOI21_X1 port map( B1 => n4220, B2 => n2104, A => n3236, ZN => n46);
   U4417 : NAND2_X1 port map( A1 => DataP_npc_1_port, A2 => n3232, ZN => n43);
   U4418 : AOI21_X1 port map( B1 => n4221, B2 => n2104, A => n3236, ZN => n42);
   U4419 : NAND2_X1 port map( A1 => DataP_npc_0_port, A2 => n3232, ZN => n39);
   U4420 : AOI21_X1 port map( B1 => n4223, B2 => n2104, A => n3235, ZN => n38);

end SYN_structural;
