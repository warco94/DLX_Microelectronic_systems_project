

    module dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11 ( 
        Clk, Rst, OPCODE_IN, FUNC_IN, MUXA_SEL, MUXB_SEL, BR_EN, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), DRAM_RW, DRAM_EN, DRAM_SEL, WB_MUX_SEL, RF_WE );
  input [5:0] OPCODE_IN;
  input [10:0] FUNC_IN;
  output [2:0] DRAM_SEL;
  output [1:0] WB_MUX_SEL;
  input Clk, Rst;
  output MUXA_SEL, MUXB_SEL, BR_EN, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , DRAM_RW, DRAM_EN,
         RF_WE;
  wire   n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n138, n139, n140, n141;
  wire   [4:0] ALU_OPCODE;
  wire   [10:0] cw;
  wire   [7:0] cw1;
  wire   [2:0] cw2;
  wire   [4:0] aluOpcode_i;

  DFFR_X1 \aluOpcode1_reg[4]  ( .D(aluOpcode_i[4]), .CK(Clk), .RN(n4), .Q(
        ALU_OPCODE[4]) );
  DFFR_X1 \aluOpcode1_reg[3]  ( .D(aluOpcode_i[3]), .CK(Clk), .RN(n6), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode1_reg[2]  ( .D(aluOpcode_i[2]), .CK(Clk), .RN(n6), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \cw1_reg[10]  ( .D(cw[10]), .CK(Clk), .RN(n5), .Q(MUXA_SEL) );
  DFFR_X1 \cw1_reg[9]  ( .D(cw[9]), .CK(Clk), .RN(n5), .Q(MUXB_SEL) );
  DFFR_X1 \cw1_reg[8]  ( .D(cw[8]), .CK(Clk), .RN(n5), .Q(BR_EN) );
  SDFFR_X1 \cw1_reg[7]  ( .D(n110), .SI(1'b0), .SE(n47), .CK(Clk), .RN(n6), 
        .Q(cw1[7]) );
  DFFR_X1 \cw1_reg[6]  ( .D(n12), .CK(Clk), .RN(n5), .Q(cw1[6]) );
  DFFR_X1 \cw1_reg[5]  ( .D(cw[5]), .CK(Clk), .RN(n5), .Q(cw1[5]) );
  DFFR_X1 \cw1_reg[4]  ( .D(cw[4]), .CK(Clk), .RN(n5), .Q(cw1[4]) );
  DFFR_X1 \cw1_reg[3]  ( .D(cw[3]), .CK(Clk), .RN(n5), .Q(cw1[3]) );
  DFFR_X1 \cw1_reg[2]  ( .D(n11), .CK(Clk), .RN(n5), .Q(cw1[2]) );
  DFFR_X1 \cw1_reg[1]  ( .D(cw[1]), .CK(Clk), .RN(n5), .Q(cw1[1]) );
  DFFR_X1 \cw1_reg[0]  ( .D(cw[0]), .CK(Clk), .RN(n4), .Q(cw1[0]) );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(Clk), .RN(n4), .Q(DRAM_RW) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(Clk), .RN(n4), .Q(DRAM_EN) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(Clk), .RN(n4), .Q(DRAM_SEL[2]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(Clk), .RN(n4), .Q(DRAM_SEL[1]) );
  DFFR_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(Clk), .RN(n4), .Q(DRAM_SEL[0]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(Clk), .RN(n4), .Q(cw2[2]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(Clk), .RN(n4), .Q(cw2[1]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(Clk), .RN(n4), .Q(cw2[0]) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .CK(Clk), .RN(n4), .Q(WB_MUX_SEL[1]) );
  DFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .CK(Clk), .RN(n4), .Q(WB_MUX_SEL[0]) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .CK(Clk), .RN(n5), .Q(RF_WE) );
  NAND3_X1 U132 ( .A1(n52), .A2(n28), .A3(n30), .ZN(n49) );
  XOR2_X1 U133 ( .A(n31), .B(OPCODE_IN[2]), .Z(n42) );
  OAI33_X1 U134 ( .A1(n45), .A2(n3), .A3(OPCODE_IN[2]), .B1(n62), .B2(n31), 
        .B3(n24), .ZN(n61) );
  NAND3_X1 U135 ( .A1(OPCODE_IN[2]), .A2(n3), .A3(n30), .ZN(n64) );
  NAND3_X1 U136 ( .A1(n31), .A2(n27), .A3(n52), .ZN(n58) );
  NAND3_X1 U137 ( .A1(n91), .A2(n140), .A3(n16), .ZN(n80) );
  NAND3_X1 U138 ( .A1(n103), .A2(n33), .A3(n19), .ZN(n102) );
  OAI33_X1 U139 ( .A1(n92), .A2(FUNC_IN[1]), .A3(n104), .B1(n105), .B2(n106), 
        .B3(n37), .ZN(n96) );
  NAND3_X1 U140 ( .A1(n30), .A2(n20), .A3(n25), .ZN(n88) );
  NAND3_X1 U141 ( .A1(n77), .A2(n141), .A3(n15), .ZN(n113) );
  NAND3_X1 U142 ( .A1(n101), .A2(n100), .A3(n127), .ZN(n126) );
  NAND3_X1 U143 ( .A1(n15), .A2(FUNC_IN[4]), .A3(n78), .ZN(n127) );
  NAND3_X1 U144 ( .A1(n128), .A2(n22), .A3(n32), .ZN(n100) );
  NAND3_X1 U145 ( .A1(n26), .A2(n30), .A3(n19), .ZN(n101) );
  NAND3_X1 U146 ( .A1(OPCODE_IN[2]), .A2(n3), .A3(OPCODE_IN[3]), .ZN(n121) );
  NAND3_X1 U147 ( .A1(n3), .A2(n20), .A3(n103), .ZN(n73) );
  NAND3_X1 U148 ( .A1(n3), .A2(n20), .A3(n128), .ZN(n72) );
  NAND3_X1 U149 ( .A1(n128), .A2(n22), .A3(n33), .ZN(n66) );
  NAND3_X1 U150 ( .A1(n3), .A2(n20), .A3(n26), .ZN(n90) );
  NAND3_X1 U151 ( .A1(n17), .A2(n141), .A3(n109), .ZN(n112) );
  OAI33_X1 U152 ( .A1(n141), .A2(n108), .A3(n139), .B1(n86), .B2(FUNC_IN[3]), 
        .B3(FUNC_IN[2]), .ZN(n135) );
  NAND3_X1 U153 ( .A1(OPCODE_IN[3]), .A2(OPCODE_IN[2]), .A3(n19), .ZN(n111) );
  DFFR_X1 \aluOpcode1_reg[0]  ( .D(aluOpcode_i[0]), .CK(Clk), .RN(n5), .Q(
        ALU_OPCODE[0]) );
  DFFR_X1 \aluOpcode1_reg[1]  ( .D(aluOpcode_i[1]), .CK(Clk), .RN(n5), .Q(
        ALU_OPCODE[1]) );
  OR2_X1 U4 ( .A1(n47), .A2(n32), .ZN(n2) );
  NOR2_X1 U5 ( .A1(n32), .A2(n33), .ZN(n74) );
  OAI21_X1 U6 ( .B1(n45), .B2(n72), .A(n100), .ZN(n70) );
  INV_X1 U7 ( .A(n57), .ZN(n19) );
  INV_X1 U8 ( .A(n72), .ZN(n9) );
  INV_X1 U9 ( .A(n45), .ZN(n30) );
  OAI21_X1 U10 ( .B1(n45), .B2(n46), .A(n2), .ZN(cw[5]) );
  NAND2_X1 U11 ( .A1(n26), .A2(n52), .ZN(n46) );
  OR4_X1 U12 ( .A1(n98), .A2(n99), .A3(n89), .A4(n70), .ZN(n97) );
  AND3_X1 U13 ( .A1(n120), .A2(n46), .A3(n130), .ZN(n129) );
  INV_X1 U14 ( .A(n56), .ZN(n23) );
  INV_X1 U15 ( .A(n90), .ZN(n7) );
  AND2_X1 U16 ( .A1(n51), .A2(n47), .ZN(n130) );
  INV_X1 U17 ( .A(n88), .ZN(n10) );
  NOR2_X1 U18 ( .A1(n20), .A2(n3), .ZN(n52) );
  NOR4_X1 U19 ( .A1(n28), .A2(n60), .A3(n27), .A4(n48), .ZN(n75) );
  NOR3_X1 U20 ( .A1(n48), .A2(n62), .A3(n57), .ZN(n84) );
  OAI221_X1 U21 ( .B1(n112), .B2(n116), .C1(n45), .C2(n90), .A(n117), .ZN(n98)
         );
  NAND2_X1 U22 ( .A1(n37), .A2(n35), .ZN(n116) );
  NOR2_X1 U23 ( .A1(n21), .A2(n84), .ZN(n117) );
  INV_X1 U24 ( .A(n65), .ZN(n21) );
  OAI221_X1 U25 ( .B1(n86), .B2(n87), .C1(n74), .C2(n90), .A(n66), .ZN(n99) );
  NOR3_X1 U26 ( .A1(n60), .A2(n42), .A3(n27), .ZN(n56) );
  NAND4_X1 U27 ( .A1(n113), .A2(n88), .A3(n18), .A4(n114), .ZN(aluOpcode_i[1])
         );
  INV_X1 U28 ( .A(n118), .ZN(n18) );
  AOI211_X1 U29 ( .C1(n32), .C2(n9), .A(n115), .B(n98), .ZN(n114) );
  NAND2_X1 U30 ( .A1(n31), .A2(n34), .ZN(n45) );
  OAI211_X1 U31 ( .C1(n45), .C2(n111), .A(n8), .B(n132), .ZN(n115) );
  INV_X1 U32 ( .A(n99), .ZN(n8) );
  AOI221_X1 U33 ( .B1(n9), .B2(n33), .C1(n133), .C2(n78), .A(n83), .ZN(n132)
         );
  NOR2_X1 U34 ( .A1(n105), .A2(n141), .ZN(n133) );
  INV_X1 U35 ( .A(n110), .ZN(n32) );
  NOR3_X1 U36 ( .A1(n141), .A2(n86), .A3(n87), .ZN(n85) );
  INV_X1 U37 ( .A(n50), .ZN(n33) );
  NAND2_X1 U38 ( .A1(n128), .A2(n52), .ZN(n47) );
  NAND2_X1 U39 ( .A1(n20), .A2(n24), .ZN(n57) );
  NAND2_X1 U40 ( .A1(n103), .A2(n52), .ZN(n51) );
  INV_X1 U41 ( .A(n3), .ZN(n24) );
  OAI211_X1 U42 ( .C1(n34), .C2(n51), .A(n58), .B(n53), .ZN(cw[0]) );
  INV_X1 U43 ( .A(n121), .ZN(n25) );
  INV_X1 U44 ( .A(n62), .ZN(n26) );
  INV_X1 U45 ( .A(n86), .ZN(n17) );
  NAND2_X1 U46 ( .A1(n19), .A2(n128), .ZN(n120) );
  NAND4_X1 U47 ( .A1(n65), .A2(n66), .A3(n67), .A4(n68), .ZN(aluOpcode_i[4])
         );
  AOI211_X1 U48 ( .C1(n36), .C2(n69), .A(n70), .B(n71), .ZN(n68) );
  AOI21_X1 U49 ( .B1(n15), .B2(n138), .A(n75), .ZN(n67) );
  AOI21_X1 U50 ( .B1(n72), .B2(n73), .A(n74), .ZN(n71) );
  INV_X1 U51 ( .A(n111), .ZN(n13) );
  AND3_X1 U52 ( .A1(n19), .A2(n103), .A3(n32), .ZN(n83) );
  NAND4_X1 U53 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(aluOpcode_i[3])
         );
  OAI21_X1 U54 ( .B1(n25), .B2(n9), .A(n29), .ZN(n79) );
  AOI21_X1 U55 ( .B1(n7), .B2(n33), .A(n89), .ZN(n81) );
  NOR4_X1 U56 ( .A1(n10), .A2(n83), .A3(n84), .A4(n85), .ZN(n82) );
  INV_X1 U57 ( .A(n60), .ZN(n22) );
  NAND2_X1 U58 ( .A1(n101), .A2(n102), .ZN(n89) );
  INV_X1 U59 ( .A(n105), .ZN(n15) );
  NAND2_X1 U60 ( .A1(n122), .A2(n123), .ZN(aluOpcode_i[0]) );
  AOI221_X1 U61 ( .B1(n33), .B2(n124), .C1(n29), .C2(n125), .A(n126), .ZN(n123) );
  AOI211_X1 U62 ( .C1(n13), .C2(n32), .A(n131), .B(n115), .ZN(n122) );
  NAND2_X1 U63 ( .A1(n130), .A2(n73), .ZN(n124) );
  INV_X1 U64 ( .A(n108), .ZN(n16) );
  OAI22_X1 U65 ( .A1(n119), .A2(n92), .B1(n120), .B2(n74), .ZN(n118) );
  OR2_X1 U66 ( .A1(n106), .A2(n86), .ZN(n119) );
  INV_X1 U67 ( .A(n39), .ZN(n12) );
  INV_X1 U68 ( .A(n53), .ZN(n11) );
  AOI21_X1 U69 ( .B1(n141), .B2(n77), .A(n78), .ZN(n106) );
  INV_X1 U70 ( .A(n48), .ZN(n29) );
  INV_X1 U71 ( .A(n92), .ZN(n36) );
  NOR2_X1 U72 ( .A1(OPCODE_IN[2]), .A2(OPCODE_IN[3]), .ZN(n103) );
  NOR2_X1 U73 ( .A1(n27), .A2(OPCODE_IN[2]), .ZN(n128) );
  NOR3_X1 U74 ( .A1(FUNC_IN[0]), .A2(FUNC_IN[2]), .A3(n108), .ZN(n69) );
  NAND2_X1 U75 ( .A1(OPCODE_IN[2]), .A2(n27), .ZN(n62) );
  NAND4_X1 U76 ( .A1(n19), .A2(n103), .A3(n136), .A4(n137), .ZN(n86) );
  NOR4_X1 U77 ( .A1(FUNC_IN[9]), .A2(FUNC_IN[8]), .A3(FUNC_IN[7]), .A4(
        FUNC_IN[6]), .ZN(n137) );
  NOR2_X1 U78 ( .A1(FUNC_IN[10]), .A2(n45), .ZN(n136) );
  INV_X1 U79 ( .A(OPCODE_IN[1]), .ZN(n31) );
  INV_X1 U80 ( .A(OPCODE_IN[2]), .ZN(n28) );
  NOR3_X1 U81 ( .A1(n43), .A2(OPCODE_IN[5]), .A3(OPCODE_IN[3]), .ZN(cw[8]) );
  AOI22_X1 U82 ( .A1(n44), .A2(OPCODE_IN[2]), .B1(OPCODE_IN[1]), .B2(n28), 
        .ZN(n43) );
  NOR2_X1 U83 ( .A1(n3), .A2(OPCODE_IN[1]), .ZN(n44) );
  INV_X1 U84 ( .A(OPCODE_IN[3]), .ZN(n27) );
  AOI21_X1 U85 ( .B1(n20), .B2(n59), .A(n56), .ZN(n53) );
  OAI21_X1 U86 ( .B1(n50), .B2(OPCODE_IN[2]), .A(n54), .ZN(n59) );
  NAND4_X1 U87 ( .A1(n30), .A2(OPCODE_IN[3]), .A3(n22), .A4(OPCODE_IN[2]), 
        .ZN(n65) );
  NAND2_X1 U88 ( .A1(OPCODE_IN[1]), .A2(n34), .ZN(n110) );
  OAI221_X1 U89 ( .B1(n47), .B2(n50), .C1(OPCODE_IN[1]), .C2(n51), .A(n49), 
        .ZN(cw[3]) );
  OAI221_X1 U90 ( .B1(n46), .B2(n48), .C1(OPCODE_IN[1]), .C2(n47), .A(n49), 
        .ZN(cw[4]) );
  NAND2_X1 U91 ( .A1(OPCODE_IN[0]), .A2(n31), .ZN(n48) );
  INV_X1 U92 ( .A(OPCODE_IN[5]), .ZN(n20) );
  OAI22_X1 U93 ( .A1(n129), .A2(n45), .B1(n134), .B2(n92), .ZN(n131) );
  AOI21_X1 U94 ( .B1(n135), .B2(n140), .A(n14), .ZN(n134) );
  INV_X1 U95 ( .A(n112), .ZN(n14) );
  OAI21_X1 U96 ( .B1(n63), .B2(n27), .A(n64), .ZN(n41) );
  AOI211_X1 U97 ( .C1(n34), .C2(n24), .A(n28), .B(n31), .ZN(n63) );
  NAND2_X1 U98 ( .A1(OPCODE_IN[0]), .A2(OPCODE_IN[1]), .ZN(n50) );
  OAI211_X1 U99 ( .C1(OPCODE_IN[5]), .C2(n54), .A(n23), .B(n39), .ZN(cw[1]) );
  OAI211_X1 U100 ( .C1(OPCODE_IN[5]), .C2(n38), .A(n23), .B(n39), .ZN(cw[9])
         );
  AOI21_X1 U101 ( .B1(n40), .B2(n27), .A(n41), .ZN(n38) );
  OAI22_X1 U102 ( .A1(n31), .A2(n24), .B1(n3), .B2(n42), .ZN(n40) );
  OAI21_X1 U103 ( .B1(OPCODE_IN[5]), .B2(n121), .A(n129), .ZN(n125) );
  NOR2_X1 U104 ( .A1(n41), .A2(n61), .ZN(n54) );
  NAND2_X1 U105 ( .A1(n3), .A2(OPCODE_IN[5]), .ZN(n60) );
  NOR3_X1 U106 ( .A1(n57), .A2(OPCODE_IN[3]), .A3(n42), .ZN(cw[10]) );
  INV_X1 U107 ( .A(OPCODE_IN[0]), .ZN(n34) );
  NAND2_X1 U108 ( .A1(n52), .A2(n55), .ZN(n39) );
  OAI22_X1 U109 ( .A1(OPCODE_IN[3]), .A2(OPCODE_IN[1]), .B1(OPCODE_IN[2]), 
        .B2(n32), .ZN(n55) );
  NAND2_X1 U110 ( .A1(FUNC_IN[5]), .A2(n16), .ZN(n105) );
  OAI22_X1 U111 ( .A1(n92), .A2(n141), .B1(n93), .B2(n139), .ZN(n91) );
  AOI21_X1 U112 ( .B1(FUNC_IN[0]), .B2(FUNC_IN[5]), .A(n36), .ZN(n93) );
  NAND2_X1 U113 ( .A1(FUNC_IN[3]), .A2(n17), .ZN(n108) );
  OR4_X1 U114 ( .A1(n94), .A2(n95), .A3(n96), .A4(n97), .ZN(aluOpcode_i[2]) );
  AOI21_X1 U115 ( .B1(n110), .B2(n48), .A(n111), .ZN(n95) );
  NOR3_X1 U116 ( .A1(n112), .A2(FUNC_IN[4]), .A3(n140), .ZN(n94) );
  NOR2_X1 U117 ( .A1(n107), .A2(n69), .ZN(n104) );
  AND3_X1 U118 ( .A1(FUNC_IN[0]), .A2(n17), .A3(n109), .ZN(n107) );
  BUF_X1 U119 ( .A(OPCODE_IN[4]), .Z(n3) );
  NOR2_X1 U120 ( .A1(n140), .A2(FUNC_IN[2]), .ZN(n78) );
  NOR2_X1 U121 ( .A1(n139), .A2(FUNC_IN[1]), .ZN(n77) );
  INV_X1 U122 ( .A(FUNC_IN[0]), .ZN(n141) );
  NAND4_X1 U123 ( .A1(n109), .A2(FUNC_IN[1]), .A3(n37), .A4(n35), .ZN(n87) );
  NOR2_X1 U124 ( .A1(n139), .A2(FUNC_IN[3]), .ZN(n109) );
  NAND2_X1 U125 ( .A1(FUNC_IN[5]), .A2(n37), .ZN(n92) );
  INV_X1 U126 ( .A(n76), .ZN(n138) );
  AOI21_X1 U127 ( .B1(n77), .B2(FUNC_IN[4]), .A(n78), .ZN(n76) );
  INV_X1 U128 ( .A(FUNC_IN[1]), .ZN(n140) );
  INV_X1 U129 ( .A(FUNC_IN[4]), .ZN(n37) );
  INV_X1 U130 ( .A(FUNC_IN[2]), .ZN(n139) );
  INV_X1 U131 ( .A(FUNC_IN[5]), .ZN(n35) );
  BUF_X1 U154 ( .A(Rst), .Z(n5) );
  BUF_X1 U155 ( .A(Rst), .Z(n4) );
  BUF_X1 U156 ( .A(Rst), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n54, n63, n64, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n41, n42, n44, n45, n46, n47, n48, n49;

  INV_X1 U1 ( .A(SEL), .ZN(n49) );
  INV_X1 U2 ( .A(n49), .ZN(n32) );
  INV_X1 U3 ( .A(n49), .ZN(n29) );
  INV_X1 U4 ( .A(n49), .ZN(n7) );
  INV_X1 U5 ( .A(n49), .ZN(n10) );
  INV_X1 U6 ( .A(n49), .ZN(n26) );
  INV_X1 U7 ( .A(n49), .ZN(n23) );
  INV_X1 U8 ( .A(n49), .ZN(n20) );
  NAND2_X1 U9 ( .A1(B[31]), .A2(n49), .ZN(n15) );
  INV_X1 U10 ( .A(n47), .ZN(n4) );
  INV_X1 U11 ( .A(SEL), .ZN(n47) );
  INV_X1 U12 ( .A(SEL), .ZN(n46) );
  NAND2_X1 U13 ( .A1(A[0]), .A2(n1), .ZN(n2) );
  NAND2_X1 U14 ( .A1(B[0]), .A2(n49), .ZN(n3) );
  NAND2_X1 U15 ( .A1(n2), .A2(n3), .ZN(Y[0]) );
  INV_X1 U16 ( .A(n49), .ZN(n1) );
  NAND2_X1 U17 ( .A1(A[22]), .A2(n4), .ZN(n5) );
  NAND2_X1 U18 ( .A1(B[22]), .A2(n47), .ZN(n6) );
  NAND2_X1 U19 ( .A1(n5), .A2(n6), .ZN(Y[22]) );
  NAND2_X1 U20 ( .A1(A[26]), .A2(n7), .ZN(n8) );
  NAND2_X1 U21 ( .A1(B[26]), .A2(n49), .ZN(n9) );
  NAND2_X1 U22 ( .A1(n8), .A2(n9), .ZN(Y[26]) );
  NAND2_X1 U23 ( .A1(A[23]), .A2(n10), .ZN(n11) );
  NAND2_X1 U24 ( .A1(B[23]), .A2(n49), .ZN(n12) );
  NAND2_X1 U25 ( .A1(n11), .A2(n12), .ZN(Y[23]) );
  NAND2_X1 U26 ( .A1(A[31]), .A2(n13), .ZN(n14) );
  NAND2_X1 U27 ( .A1(n14), .A2(n15), .ZN(Y[31]) );
  INV_X1 U28 ( .A(n49), .ZN(n13) );
  NAND2_X1 U29 ( .A1(A[30]), .A2(n4), .ZN(n16) );
  NAND2_X1 U30 ( .A1(B[30]), .A2(n46), .ZN(n17) );
  NAND2_X1 U31 ( .A1(n16), .A2(n17), .ZN(Y[30]) );
  NAND2_X1 U32 ( .A1(A[29]), .A2(n42), .ZN(n18) );
  NAND2_X1 U33 ( .A1(B[29]), .A2(n47), .ZN(n19) );
  NAND2_X1 U34 ( .A1(n18), .A2(n19), .ZN(Y[29]) );
  NAND2_X1 U35 ( .A1(A[28]), .A2(n20), .ZN(n21) );
  NAND2_X1 U36 ( .A1(B[28]), .A2(n49), .ZN(n22) );
  NAND2_X1 U37 ( .A1(n21), .A2(n22), .ZN(Y[28]) );
  NAND2_X1 U38 ( .A1(A[21]), .A2(n23), .ZN(n24) );
  NAND2_X1 U39 ( .A1(B[21]), .A2(n49), .ZN(n25) );
  NAND2_X1 U40 ( .A1(n24), .A2(n25), .ZN(Y[21]) );
  NAND2_X1 U41 ( .A1(A[20]), .A2(n26), .ZN(n27) );
  NAND2_X1 U42 ( .A1(B[20]), .A2(n49), .ZN(n28) );
  NAND2_X1 U43 ( .A1(n27), .A2(n28), .ZN(Y[20]) );
  NAND2_X1 U44 ( .A1(A[25]), .A2(n29), .ZN(n30) );
  NAND2_X1 U45 ( .A1(B[25]), .A2(n49), .ZN(n31) );
  NAND2_X1 U46 ( .A1(n30), .A2(n31), .ZN(Y[25]) );
  NAND2_X1 U47 ( .A1(A[24]), .A2(n32), .ZN(n33) );
  NAND2_X1 U48 ( .A1(B[24]), .A2(n49), .ZN(n41) );
  NAND2_X1 U49 ( .A1(n33), .A2(n41), .ZN(Y[24]) );
  MUX2_X1 U50 ( .A(A[27]), .B(B[27]), .S(n49), .Z(Y[27]) );
  INV_X1 U51 ( .A(n49), .ZN(n44) );
  INV_X1 U52 ( .A(n48), .ZN(n42) );
  INV_X1 U53 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U54 ( .A1(n42), .A2(A[9]), .B1(B[9]), .B2(n48), .ZN(n34) );
  INV_X1 U55 ( .A(n35), .ZN(Y[8]) );
  AOI22_X1 U56 ( .A1(A[8]), .A2(n42), .B1(B[8]), .B2(n47), .ZN(n35) );
  INV_X1 U57 ( .A(n64), .ZN(Y[10]) );
  AOI22_X1 U58 ( .A1(A[10]), .A2(n42), .B1(B[10]), .B2(n46), .ZN(n64) );
  INV_X1 U59 ( .A(n63), .ZN(Y[11]) );
  AOI22_X1 U60 ( .A1(A[11]), .A2(n42), .B1(B[11]), .B2(n48), .ZN(n63) );
  INV_X1 U61 ( .A(n36), .ZN(Y[7]) );
  AOI22_X1 U62 ( .A1(A[7]), .A2(n42), .B1(B[7]), .B2(n47), .ZN(n36) );
  INV_X1 U63 ( .A(n37), .ZN(Y[6]) );
  AOI22_X1 U64 ( .A1(A[6]), .A2(n42), .B1(B[6]), .B2(n47), .ZN(n37) );
  INV_X1 U65 ( .A(n39), .ZN(Y[4]) );
  AOI22_X1 U66 ( .A1(A[4]), .A2(n42), .B1(B[4]), .B2(n46), .ZN(n39) );
  INV_X1 U67 ( .A(n38), .ZN(Y[5]) );
  AOI22_X1 U68 ( .A1(A[5]), .A2(n42), .B1(B[5]), .B2(n46), .ZN(n38) );
  INV_X1 U69 ( .A(n54), .ZN(Y[1]) );
  AOI22_X1 U70 ( .A1(A[1]), .A2(n42), .B1(B[1]), .B2(n48), .ZN(n54) );
  INV_X1 U71 ( .A(n43), .ZN(Y[2]) );
  AOI22_X1 U72 ( .A1(A[2]), .A2(n42), .B1(B[2]), .B2(n47), .ZN(n43) );
  INV_X1 U73 ( .A(n40), .ZN(Y[3]) );
  AOI22_X1 U74 ( .A1(A[3]), .A2(n42), .B1(B[3]), .B2(n46), .ZN(n40) );
  INV_X1 U75 ( .A(n49), .ZN(n45) );
  INV_X1 U76 ( .A(SEL), .ZN(n48) );
  MUX2_X1 U77 ( .A(B[12]), .B(A[12]), .S(n42), .Z(Y[12]) );
  MUX2_X1 U78 ( .A(B[13]), .B(A[13]), .S(n45), .Z(Y[13]) );
  MUX2_X1 U79 ( .A(B[14]), .B(A[14]), .S(n45), .Z(Y[14]) );
  MUX2_X1 U80 ( .A(B[15]), .B(A[15]), .S(n44), .Z(Y[15]) );
  MUX2_X1 U81 ( .A(B[16]), .B(A[16]), .S(n44), .Z(Y[16]) );
  MUX2_X1 U82 ( .A(B[17]), .B(A[17]), .S(n44), .Z(Y[17]) );
  MUX2_X1 U83 ( .A(B[18]), .B(A[18]), .S(n44), .Z(Y[18]) );
  MUX2_X1 U84 ( .A(B[19]), .B(A[19]), .S(n44), .Z(Y[19]) );
endmodule


module register_e_N32 ( D, clk, rst, O );
  input [31:0] D;
  output [31:0] O;
  input clk, rst;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3;

  DFF_X1 \O_reg[10]  ( .D(N12), .CK(clk), .Q(O[10]) );
  DFF_X1 \O_reg[9]  ( .D(N11), .CK(clk), .Q(O[9]) );
  DFF_X1 \O_reg[4]  ( .D(N6), .CK(clk), .Q(O[4]) );
  DFF_X1 \O_reg[8]  ( .D(N10), .CK(clk), .Q(O[8]) );
  DFF_X1 \O_reg[15]  ( .D(N17), .CK(clk), .Q(O[15]) );
  DFF_X1 \O_reg[14]  ( .D(N16), .CK(clk), .Q(O[14]) );
  DFF_X1 \O_reg[13]  ( .D(N15), .CK(clk), .Q(O[13]) );
  DFF_X1 \O_reg[3]  ( .D(N5), .CK(clk), .Q(O[3]) );
  DFF_X1 \O_reg[12]  ( .D(N14), .CK(clk), .Q(O[12]) );
  DFF_X1 \O_reg[28]  ( .D(N30), .CK(clk), .Q(O[28]) );
  DFF_X1 \O_reg[7]  ( .D(N9), .CK(clk), .Q(O[7]) );
  DFF_X1 \O_reg[1]  ( .D(N3), .CK(clk), .Q(O[1]) );
  DFF_X1 \O_reg[6]  ( .D(N8), .CK(clk), .Q(O[6]) );
  DFF_X1 \O_reg[5]  ( .D(N7), .CK(clk), .Q(O[5]) );
  DFF_X1 \O_reg[22]  ( .D(N24), .CK(clk), .Q(O[22]) );
  DFF_X1 \O_reg[21]  ( .D(N23), .CK(clk), .Q(O[21]) );
  DFF_X1 \O_reg[20]  ( .D(N22), .CK(clk), .Q(O[20]) );
  DFF_X1 \O_reg[11]  ( .D(N13), .CK(clk), .Q(O[11]) );
  DFF_X1 \O_reg[16]  ( .D(N18), .CK(clk), .Q(O[16]) );
  DFF_X1 \O_reg[0]  ( .D(N2), .CK(clk), .Q(O[0]) );
  DFF_X1 \O_reg[2]  ( .D(N4), .CK(clk), .Q(O[2]) );
  DFF_X1 \O_reg[19]  ( .D(N21), .CK(clk), .Q(O[19]) );
  DFF_X1 \O_reg[18]  ( .D(N20), .CK(clk), .Q(O[18]) );
  DFF_X1 \O_reg[17]  ( .D(N19), .CK(clk), .Q(O[17]) );
  DFF_X1 \O_reg[30]  ( .D(N32), .CK(clk), .Q(O[30]) );
  DFF_X1 \O_reg[29]  ( .D(N31), .CK(clk), .Q(O[29]) );
  DFF_X1 \O_reg[23]  ( .D(N25), .CK(clk), .Q(O[23]) );
  DFF_X1 \O_reg[26]  ( .D(N28), .CK(clk), .Q(O[26]) );
  DFF_X1 \O_reg[25]  ( .D(N27), .CK(clk), .Q(O[25]) );
  DFF_X1 \O_reg[24]  ( .D(N26), .CK(clk), .Q(O[24]) );
  DFF_X1 \O_reg[31]  ( .D(N33), .CK(clk), .Q(O[31]) );
  DFF_X1 \O_reg[27]  ( .D(N29), .CK(clk), .Q(O[27]) );
  BUF_X1 U3 ( .A(rst), .Z(n1) );
  BUF_X1 U4 ( .A(rst), .Z(n2) );
  BUF_X1 U5 ( .A(rst), .Z(n3) );
  AND2_X1 U6 ( .A1(D[9]), .A2(n1), .ZN(N11) );
  AND2_X1 U7 ( .A1(D[8]), .A2(n1), .ZN(N10) );
  AND2_X1 U8 ( .A1(D[10]), .A2(n1), .ZN(N12) );
  AND2_X1 U9 ( .A1(D[11]), .A2(n1), .ZN(N13) );
  AND2_X1 U10 ( .A1(n1), .A2(D[7]), .ZN(N9) );
  AND2_X1 U11 ( .A1(D[6]), .A2(n1), .ZN(N8) );
  AND2_X1 U12 ( .A1(D[4]), .A2(n1), .ZN(N6) );
  AND2_X1 U13 ( .A1(D[5]), .A2(n1), .ZN(N7) );
  AND2_X1 U14 ( .A1(D[1]), .A2(n1), .ZN(N3) );
  AND2_X1 U15 ( .A1(D[2]), .A2(n1), .ZN(N4) );
  AND2_X1 U16 ( .A1(D[3]), .A2(n1), .ZN(N5) );
  AND2_X1 U17 ( .A1(D[0]), .A2(n2), .ZN(N2) );
  AND2_X1 U18 ( .A1(D[12]), .A2(n1), .ZN(N14) );
  AND2_X1 U19 ( .A1(D[13]), .A2(n3), .ZN(N15) );
  AND2_X1 U20 ( .A1(D[14]), .A2(n3), .ZN(N16) );
  AND2_X1 U21 ( .A1(D[15]), .A2(n3), .ZN(N17) );
  AND2_X1 U22 ( .A1(D[16]), .A2(n3), .ZN(N18) );
  AND2_X1 U23 ( .A1(D[17]), .A2(n2), .ZN(N19) );
  AND2_X1 U24 ( .A1(D[18]), .A2(n2), .ZN(N20) );
  AND2_X1 U25 ( .A1(D[19]), .A2(n2), .ZN(N21) );
  AND2_X1 U26 ( .A1(D[20]), .A2(n2), .ZN(N22) );
  AND2_X1 U27 ( .A1(D[21]), .A2(n2), .ZN(N23) );
  AND2_X1 U28 ( .A1(D[22]), .A2(n2), .ZN(N24) );
  AND2_X1 U29 ( .A1(D[23]), .A2(n2), .ZN(N25) );
  AND2_X1 U30 ( .A1(D[24]), .A2(n2), .ZN(N26) );
  AND2_X1 U31 ( .A1(D[25]), .A2(n2), .ZN(N27) );
  AND2_X1 U32 ( .A1(D[26]), .A2(n2), .ZN(N28) );
  AND2_X1 U33 ( .A1(D[27]), .A2(n2), .ZN(N29) );
  AND2_X1 U34 ( .A1(D[28]), .A2(n2), .ZN(N30) );
  AND2_X1 U35 ( .A1(D[29]), .A2(n2), .ZN(N31) );
  AND2_X1 U36 ( .A1(D[30]), .A2(n2), .ZN(N32) );
  AND2_X1 U37 ( .A1(D[31]), .A2(n2), .ZN(N33) );
endmodule


module branch_predictor_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module branch_predictor_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X1 U1 ( .A1(A[6]), .A2(n2), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[5]), .A2(n3), .ZN(n2) );
  NAND2_X1 U3 ( .A1(A[30]), .A2(n27), .ZN(n57) );
  AND2_X1 U4 ( .A1(A[4]), .A2(n4), .ZN(n3) );
  AND2_X1 U5 ( .A1(A[3]), .A2(A[2]), .ZN(n4) );
  AND2_X1 U6 ( .A1(A[7]), .A2(n1), .ZN(n5) );
  AND2_X1 U7 ( .A1(A[8]), .A2(n5), .ZN(n6) );
  AND2_X1 U8 ( .A1(A[9]), .A2(n6), .ZN(n7) );
  AND2_X1 U9 ( .A1(A[10]), .A2(n7), .ZN(n8) );
  AND2_X1 U10 ( .A1(A[11]), .A2(n8), .ZN(n9) );
  AND2_X1 U11 ( .A1(A[12]), .A2(n9), .ZN(n10) );
  AND2_X1 U12 ( .A1(A[13]), .A2(n10), .ZN(n11) );
  AND2_X1 U13 ( .A1(A[14]), .A2(n11), .ZN(n12) );
  AND2_X1 U14 ( .A1(A[15]), .A2(n12), .ZN(n13) );
  AND2_X1 U15 ( .A1(A[16]), .A2(n13), .ZN(n14) );
  AND2_X1 U16 ( .A1(A[17]), .A2(n14), .ZN(n15) );
  AND2_X1 U17 ( .A1(A[18]), .A2(n15), .ZN(n16) );
  AND2_X1 U18 ( .A1(A[19]), .A2(n16), .ZN(n17) );
  AND2_X1 U19 ( .A1(A[20]), .A2(n17), .ZN(n18) );
  AND2_X1 U20 ( .A1(A[21]), .A2(n18), .ZN(n19) );
  AND2_X1 U21 ( .A1(A[22]), .A2(n19), .ZN(n20) );
  AND2_X1 U22 ( .A1(A[23]), .A2(n20), .ZN(n21) );
  AND2_X1 U23 ( .A1(A[24]), .A2(n21), .ZN(n22) );
  AND2_X1 U24 ( .A1(A[25]), .A2(n22), .ZN(n23) );
  AND2_X1 U25 ( .A1(A[26]), .A2(n23), .ZN(n24) );
  AND2_X1 U26 ( .A1(A[27]), .A2(n24), .ZN(n25) );
  AND2_X1 U27 ( .A1(A[28]), .A2(n25), .ZN(n26) );
  AND2_X1 U28 ( .A1(A[29]), .A2(n26), .ZN(n27) );
  XOR2_X1 U29 ( .A(A[6]), .B(n2), .Z(SUM[6]) );
  XOR2_X1 U30 ( .A(A[7]), .B(n1), .Z(SUM[7]) );
  XOR2_X1 U31 ( .A(A[8]), .B(n5), .Z(SUM[8]) );
  XOR2_X1 U32 ( .A(A[9]), .B(n6), .Z(SUM[9]) );
  XOR2_X1 U33 ( .A(A[10]), .B(n7), .Z(SUM[10]) );
  XOR2_X1 U34 ( .A(A[11]), .B(n8), .Z(SUM[11]) );
  XOR2_X1 U35 ( .A(A[12]), .B(n9), .Z(SUM[12]) );
  XOR2_X1 U36 ( .A(A[13]), .B(n10), .Z(SUM[13]) );
  XOR2_X1 U37 ( .A(A[15]), .B(n12), .Z(SUM[15]) );
  XOR2_X1 U38 ( .A(A[16]), .B(n13), .Z(SUM[16]) );
  XOR2_X1 U39 ( .A(A[17]), .B(n14), .Z(SUM[17]) );
  XOR2_X1 U40 ( .A(A[18]), .B(n15), .Z(SUM[18]) );
  XOR2_X1 U41 ( .A(A[19]), .B(n16), .Z(SUM[19]) );
  XOR2_X1 U42 ( .A(A[20]), .B(n17), .Z(SUM[20]) );
  XOR2_X1 U43 ( .A(A[21]), .B(n18), .Z(SUM[21]) );
  XOR2_X1 U44 ( .A(A[22]), .B(n19), .Z(SUM[22]) );
  XOR2_X1 U45 ( .A(A[23]), .B(n20), .Z(SUM[23]) );
  XOR2_X1 U46 ( .A(A[24]), .B(n21), .Z(SUM[24]) );
  XOR2_X1 U47 ( .A(A[25]), .B(n22), .Z(SUM[25]) );
  XOR2_X1 U48 ( .A(A[26]), .B(n23), .Z(SUM[26]) );
  XOR2_X1 U49 ( .A(A[14]), .B(n11), .Z(SUM[14]) );
  XOR2_X1 U50 ( .A(A[27]), .B(n24), .Z(SUM[27]) );
  XOR2_X1 U51 ( .A(A[28]), .B(n25), .Z(SUM[28]) );
  XOR2_X1 U52 ( .A(A[29]), .B(n26), .Z(SUM[29]) );
  XOR2_X1 U53 ( .A(A[30]), .B(n27), .Z(SUM[30]) );
  XNOR2_X1 U54 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  INV_X1 U55 ( .A(A[2]), .ZN(SUM[2]) );
  XOR2_X1 U56 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U57 ( .A(A[4]), .B(n4), .Z(SUM[4]) );
  XOR2_X1 U58 ( .A(A[5]), .B(n3), .Z(SUM[5]) );
endmodule


module branch_predictor_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module branch_predictor_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module branch_predictor ( RST, PC_IN, PC_FAIL, IR_IN, IR_FAIL, WRONG_PRE, 
        RIGHT_PRE, NPC_OUT, LINK_ADD, SEL, TAKEN );
  input [31:0] PC_IN;
  input [31:0] PC_FAIL;
  input [31:0] IR_IN;
  input [15:0] IR_FAIL;
  output [31:0] NPC_OUT;
  output [31:0] LINK_ADD;
  input RST, WRONG_PRE, RIGHT_PRE;
  output SEL, TAKEN;
  wire   \CACHE_mem[0][1] , \CACHE_mem[0][0] , \CACHE_mem[1][1] ,
         \CACHE_mem[1][0] , \CACHE_mem[2][1] , \CACHE_mem[2][0] ,
         \CACHE_mem[3][1] , \CACHE_mem[3][0] , \CACHE_mem[4][1] ,
         \CACHE_mem[4][0] , \CACHE_mem[5][1] , \CACHE_mem[5][0] ,
         \CACHE_mem[6][1] , \CACHE_mem[6][0] , \CACHE_mem[7][1] ,
         \CACHE_mem[7][0] , \CACHE_mem[8][1] , \CACHE_mem[8][0] ,
         \CACHE_mem[9][1] , \CACHE_mem[9][0] , \CACHE_mem[10][1] ,
         \CACHE_mem[10][0] , \CACHE_mem[11][1] , \CACHE_mem[11][0] ,
         \CACHE_mem[12][1] , \CACHE_mem[12][0] , \CACHE_mem[13][1] ,
         \CACHE_mem[13][0] , \CACHE_mem[14][1] , \CACHE_mem[14][0] ,
         \CACHE_mem[15][1] , \CACHE_mem[15][0] , \CACHE_mem[16][1] ,
         \CACHE_mem[16][0] , \CACHE_mem[17][1] , \CACHE_mem[17][0] ,
         \CACHE_mem[18][1] , \CACHE_mem[18][0] , \CACHE_mem[19][1] ,
         \CACHE_mem[19][0] , \CACHE_mem[20][1] , \CACHE_mem[20][0] ,
         \CACHE_mem[21][1] , \CACHE_mem[21][0] , \CACHE_mem[22][1] ,
         \CACHE_mem[22][0] , \CACHE_mem[23][1] , \CACHE_mem[23][0] ,
         \CACHE_mem[24][1] , \CACHE_mem[24][0] , \CACHE_mem[25][1] ,
         \CACHE_mem[25][0] , \CACHE_mem[26][1] , \CACHE_mem[26][0] ,
         \CACHE_mem[27][1] , \CACHE_mem[27][0] , \CACHE_mem[28][1] ,
         \CACHE_mem[28][0] , \CACHE_mem[29][1] , \CACHE_mem[29][0] ,
         \CACHE_mem[30][1] , \CACHE_mem[30][0] , \CACHE_mem[31][1] ,
         \CACHE_mem[31][0] , N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N216, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N323, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N479, N480, N612, N613, N614, N615, N616, N617, N618, N619,
         N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630,
         N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641,
         N642, N643, N644, N645, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239;

  DLH_X1 \NPC_OUT_reg[31]  ( .G(n188), .D(n199), .Q(NPC_OUT[31]) );
  DLH_X1 \NPC_OUT_reg[30]  ( .G(n188), .D(n200), .Q(NPC_OUT[30]) );
  DLH_X1 \NPC_OUT_reg[29]  ( .G(n188), .D(n201), .Q(NPC_OUT[29]) );
  DLH_X1 \NPC_OUT_reg[28]  ( .G(n188), .D(n202), .Q(NPC_OUT[28]) );
  DLH_X1 \NPC_OUT_reg[27]  ( .G(n188), .D(n203), .Q(NPC_OUT[27]) );
  DLH_X1 \NPC_OUT_reg[26]  ( .G(n188), .D(n204), .Q(NPC_OUT[26]) );
  DLH_X1 \NPC_OUT_reg[25]  ( .G(n188), .D(n205), .Q(NPC_OUT[25]) );
  DLH_X1 \NPC_OUT_reg[24]  ( .G(n188), .D(n206), .Q(NPC_OUT[24]) );
  DLH_X1 \NPC_OUT_reg[23]  ( .G(n188), .D(n207), .Q(NPC_OUT[23]) );
  DLH_X1 \NPC_OUT_reg[22]  ( .G(n188), .D(n208), .Q(NPC_OUT[22]) );
  DLH_X1 \NPC_OUT_reg[21]  ( .G(n188), .D(n209), .Q(NPC_OUT[21]) );
  DLH_X1 \NPC_OUT_reg[20]  ( .G(n189), .D(n210), .Q(NPC_OUT[20]) );
  DLH_X1 \NPC_OUT_reg[19]  ( .G(n189), .D(n211), .Q(NPC_OUT[19]) );
  DLH_X1 \NPC_OUT_reg[18]  ( .G(n189), .D(n212), .Q(NPC_OUT[18]) );
  DLH_X1 \NPC_OUT_reg[17]  ( .G(n189), .D(n213), .Q(NPC_OUT[17]) );
  DLH_X1 \NPC_OUT_reg[16]  ( .G(n189), .D(n214), .Q(NPC_OUT[16]) );
  DLH_X1 \NPC_OUT_reg[15]  ( .G(n189), .D(n215), .Q(NPC_OUT[15]) );
  DLH_X1 \NPC_OUT_reg[14]  ( .G(n189), .D(n216), .Q(NPC_OUT[14]) );
  DLH_X1 \NPC_OUT_reg[13]  ( .G(n189), .D(n217), .Q(NPC_OUT[13]) );
  DLH_X1 \NPC_OUT_reg[12]  ( .G(n189), .D(n218), .Q(NPC_OUT[12]) );
  DLH_X1 \NPC_OUT_reg[11]  ( .G(n189), .D(n219), .Q(NPC_OUT[11]) );
  DLH_X1 \NPC_OUT_reg[10]  ( .G(n189), .D(n220), .Q(NPC_OUT[10]) );
  DLH_X1 \NPC_OUT_reg[9]  ( .G(n190), .D(n221), .Q(NPC_OUT[9]) );
  DLH_X1 \NPC_OUT_reg[8]  ( .G(n190), .D(n222), .Q(NPC_OUT[8]) );
  DLH_X1 \NPC_OUT_reg[7]  ( .G(n190), .D(n223), .Q(NPC_OUT[7]) );
  DLH_X1 \NPC_OUT_reg[6]  ( .G(n190), .D(n224), .Q(NPC_OUT[6]) );
  DLH_X1 \NPC_OUT_reg[5]  ( .G(n190), .D(n225), .Q(NPC_OUT[5]) );
  DLH_X1 \NPC_OUT_reg[4]  ( .G(n190), .D(n226), .Q(NPC_OUT[4]) );
  DLH_X1 \NPC_OUT_reg[3]  ( .G(n190), .D(n227), .Q(NPC_OUT[3]) );
  DLH_X1 \NPC_OUT_reg[2]  ( .G(n190), .D(n228), .Q(NPC_OUT[2]) );
  DLH_X1 \NPC_OUT_reg[1]  ( .G(n190), .D(n229), .Q(NPC_OUT[1]) );
  DLH_X1 \NPC_OUT_reg[0]  ( .G(n190), .D(n230), .Q(NPC_OUT[0]) );
  DLH_X1 \LINK_ADD_reg[31]  ( .G(n186), .D(N388), .Q(LINK_ADD[31]) );
  DLH_X1 \LINK_ADD_reg[30]  ( .G(n186), .D(N387), .Q(LINK_ADD[30]) );
  DLH_X1 \LINK_ADD_reg[29]  ( .G(n186), .D(N386), .Q(LINK_ADD[29]) );
  DLH_X1 \LINK_ADD_reg[28]  ( .G(n186), .D(N385), .Q(LINK_ADD[28]) );
  DLH_X1 \LINK_ADD_reg[27]  ( .G(n186), .D(N384), .Q(LINK_ADD[27]) );
  DLH_X1 \LINK_ADD_reg[26]  ( .G(n186), .D(N383), .Q(LINK_ADD[26]) );
  DLH_X1 \LINK_ADD_reg[25]  ( .G(n186), .D(N382), .Q(LINK_ADD[25]) );
  DLH_X1 \LINK_ADD_reg[24]  ( .G(n186), .D(N381), .Q(LINK_ADD[24]) );
  DLH_X1 \LINK_ADD_reg[23]  ( .G(n186), .D(N380), .Q(LINK_ADD[23]) );
  DLH_X1 \LINK_ADD_reg[22]  ( .G(n186), .D(N379), .Q(LINK_ADD[22]) );
  DLH_X1 \LINK_ADD_reg[21]  ( .G(n186), .D(N378), .Q(LINK_ADD[21]) );
  DLH_X1 \LINK_ADD_reg[20]  ( .G(n186), .D(N377), .Q(LINK_ADD[20]) );
  DLH_X1 \LINK_ADD_reg[19]  ( .G(n186), .D(N376), .Q(LINK_ADD[19]) );
  DLH_X1 \LINK_ADD_reg[18]  ( .G(n186), .D(N375), .Q(LINK_ADD[18]) );
  DLH_X1 \LINK_ADD_reg[17]  ( .G(n186), .D(N374), .Q(LINK_ADD[17]) );
  DLH_X1 \LINK_ADD_reg[16]  ( .G(n186), .D(N373), .Q(LINK_ADD[16]) );
  DLH_X1 \LINK_ADD_reg[15]  ( .G(n186), .D(N372), .Q(LINK_ADD[15]) );
  DLH_X1 \LINK_ADD_reg[14]  ( .G(n186), .D(N371), .Q(LINK_ADD[14]) );
  DLH_X1 \LINK_ADD_reg[13]  ( .G(n186), .D(N370), .Q(LINK_ADD[13]) );
  DLH_X1 \LINK_ADD_reg[12]  ( .G(n186), .D(N369), .Q(LINK_ADD[12]) );
  DLH_X1 \LINK_ADD_reg[11]  ( .G(n186), .D(N368), .Q(LINK_ADD[11]) );
  DLH_X1 \LINK_ADD_reg[10]  ( .G(n186), .D(N367), .Q(LINK_ADD[10]) );
  DLH_X1 \LINK_ADD_reg[9]  ( .G(n186), .D(N366), .Q(LINK_ADD[9]) );
  DLH_X1 \LINK_ADD_reg[8]  ( .G(n186), .D(N365), .Q(LINK_ADD[8]) );
  DLH_X1 \LINK_ADD_reg[7]  ( .G(n187), .D(N364), .Q(LINK_ADD[7]) );
  DLH_X1 \LINK_ADD_reg[6]  ( .G(n187), .D(N363), .Q(LINK_ADD[6]) );
  DLH_X1 \LINK_ADD_reg[5]  ( .G(n187), .D(N362), .Q(LINK_ADD[5]) );
  DLH_X1 \LINK_ADD_reg[4]  ( .G(n187), .D(N361), .Q(LINK_ADD[4]) );
  DLH_X1 \LINK_ADD_reg[3]  ( .G(n187), .D(N360), .Q(LINK_ADD[3]) );
  DLH_X1 \LINK_ADD_reg[2]  ( .G(n187), .D(N359), .Q(LINK_ADD[2]) );
  DLH_X1 \LINK_ADD_reg[1]  ( .G(n187), .D(N358), .Q(LINK_ADD[1]) );
  DLH_X1 \LINK_ADD_reg[0]  ( .G(n187), .D(N357), .Q(LINK_ADD[0]) );
  DLH_X1 \CACHE_mem_reg[0][1]  ( .G(N643), .D(n180), .Q(\CACHE_mem[0][1] ) );
  DLH_X1 \CACHE_mem_reg[0][0]  ( .G(N643), .D(n183), .Q(\CACHE_mem[0][0] ) );
  DLH_X1 \CACHE_mem_reg[1][1]  ( .G(N642), .D(n180), .Q(\CACHE_mem[1][1] ) );
  DLH_X1 \CACHE_mem_reg[1][0]  ( .G(N642), .D(n183), .Q(\CACHE_mem[1][0] ) );
  DLH_X1 \CACHE_mem_reg[2][1]  ( .G(N641), .D(n180), .Q(\CACHE_mem[2][1] ) );
  DLH_X1 \CACHE_mem_reg[2][0]  ( .G(N641), .D(n183), .Q(\CACHE_mem[2][0] ) );
  DLH_X1 \CACHE_mem_reg[3][1]  ( .G(N640), .D(n180), .Q(\CACHE_mem[3][1] ) );
  DLH_X1 \CACHE_mem_reg[3][0]  ( .G(N640), .D(n183), .Q(\CACHE_mem[3][0] ) );
  DLH_X1 \CACHE_mem_reg[4][1]  ( .G(N639), .D(n180), .Q(\CACHE_mem[4][1] ) );
  DLH_X1 \CACHE_mem_reg[4][0]  ( .G(N639), .D(n183), .Q(\CACHE_mem[4][0] ) );
  DLH_X1 \CACHE_mem_reg[5][1]  ( .G(N638), .D(n180), .Q(\CACHE_mem[5][1] ) );
  DLH_X1 \CACHE_mem_reg[5][0]  ( .G(N638), .D(n183), .Q(\CACHE_mem[5][0] ) );
  DLH_X1 \CACHE_mem_reg[6][1]  ( .G(N637), .D(n180), .Q(\CACHE_mem[6][1] ) );
  DLH_X1 \CACHE_mem_reg[6][0]  ( .G(N637), .D(n183), .Q(\CACHE_mem[6][0] ) );
  DLH_X1 \CACHE_mem_reg[7][1]  ( .G(N636), .D(n180), .Q(\CACHE_mem[7][1] ) );
  DLH_X1 \CACHE_mem_reg[7][0]  ( .G(N636), .D(n183), .Q(\CACHE_mem[7][0] ) );
  DLH_X1 \CACHE_mem_reg[8][1]  ( .G(N635), .D(n180), .Q(\CACHE_mem[8][1] ) );
  DLH_X1 \CACHE_mem_reg[8][0]  ( .G(N635), .D(n183), .Q(\CACHE_mem[8][0] ) );
  DLH_X1 \CACHE_mem_reg[9][1]  ( .G(N634), .D(n180), .Q(\CACHE_mem[9][1] ) );
  DLH_X1 \CACHE_mem_reg[9][0]  ( .G(N634), .D(n183), .Q(\CACHE_mem[9][0] ) );
  DLH_X1 \CACHE_mem_reg[10][1]  ( .G(N633), .D(n180), .Q(\CACHE_mem[10][1] )
         );
  DLH_X1 \CACHE_mem_reg[10][0]  ( .G(N633), .D(n183), .Q(\CACHE_mem[10][0] )
         );
  DLH_X1 \CACHE_mem_reg[11][1]  ( .G(N632), .D(n181), .Q(\CACHE_mem[11][1] )
         );
  DLH_X1 \CACHE_mem_reg[11][0]  ( .G(N632), .D(n184), .Q(\CACHE_mem[11][0] )
         );
  DLH_X1 \CACHE_mem_reg[12][1]  ( .G(N631), .D(n181), .Q(\CACHE_mem[12][1] )
         );
  DLH_X1 \CACHE_mem_reg[12][0]  ( .G(N631), .D(n184), .Q(\CACHE_mem[12][0] )
         );
  DLH_X1 \CACHE_mem_reg[13][1]  ( .G(N630), .D(n181), .Q(\CACHE_mem[13][1] )
         );
  DLH_X1 \CACHE_mem_reg[13][0]  ( .G(N630), .D(n184), .Q(\CACHE_mem[13][0] )
         );
  DLH_X1 \CACHE_mem_reg[14][1]  ( .G(N629), .D(n181), .Q(\CACHE_mem[14][1] )
         );
  DLH_X1 \CACHE_mem_reg[14][0]  ( .G(N629), .D(n184), .Q(\CACHE_mem[14][0] )
         );
  DLH_X1 \CACHE_mem_reg[15][1]  ( .G(N628), .D(n181), .Q(\CACHE_mem[15][1] )
         );
  DLH_X1 \CACHE_mem_reg[15][0]  ( .G(N628), .D(n184), .Q(\CACHE_mem[15][0] )
         );
  DLH_X1 \CACHE_mem_reg[16][1]  ( .G(N627), .D(n181), .Q(\CACHE_mem[16][1] )
         );
  DLH_X1 \CACHE_mem_reg[16][0]  ( .G(N627), .D(n184), .Q(\CACHE_mem[16][0] )
         );
  DLH_X1 \CACHE_mem_reg[17][1]  ( .G(N626), .D(n181), .Q(\CACHE_mem[17][1] )
         );
  DLH_X1 \CACHE_mem_reg[17][0]  ( .G(N626), .D(n184), .Q(\CACHE_mem[17][0] )
         );
  DLH_X1 \CACHE_mem_reg[18][1]  ( .G(N625), .D(n181), .Q(\CACHE_mem[18][1] )
         );
  DLH_X1 \CACHE_mem_reg[18][0]  ( .G(N625), .D(n184), .Q(\CACHE_mem[18][0] )
         );
  DLH_X1 \CACHE_mem_reg[19][1]  ( .G(N624), .D(n181), .Q(\CACHE_mem[19][1] )
         );
  DLH_X1 \CACHE_mem_reg[19][0]  ( .G(N624), .D(n184), .Q(\CACHE_mem[19][0] )
         );
  DLH_X1 \CACHE_mem_reg[20][1]  ( .G(N623), .D(n181), .Q(\CACHE_mem[20][1] )
         );
  DLH_X1 \CACHE_mem_reg[20][0]  ( .G(N623), .D(n184), .Q(\CACHE_mem[20][0] )
         );
  DLH_X1 \CACHE_mem_reg[21][1]  ( .G(N622), .D(n181), .Q(\CACHE_mem[21][1] )
         );
  DLH_X1 \CACHE_mem_reg[21][0]  ( .G(N622), .D(n184), .Q(\CACHE_mem[21][0] )
         );
  DLH_X1 \CACHE_mem_reg[22][1]  ( .G(N621), .D(n182), .Q(\CACHE_mem[22][1] )
         );
  DLH_X1 \CACHE_mem_reg[22][0]  ( .G(N621), .D(n185), .Q(\CACHE_mem[22][0] )
         );
  DLH_X1 \CACHE_mem_reg[23][1]  ( .G(N620), .D(n182), .Q(\CACHE_mem[23][1] )
         );
  DLH_X1 \CACHE_mem_reg[23][0]  ( .G(N620), .D(n185), .Q(\CACHE_mem[23][0] )
         );
  DLH_X1 \CACHE_mem_reg[24][1]  ( .G(N619), .D(n182), .Q(\CACHE_mem[24][1] )
         );
  DLH_X1 \CACHE_mem_reg[24][0]  ( .G(N619), .D(n185), .Q(\CACHE_mem[24][0] )
         );
  DLH_X1 \CACHE_mem_reg[25][1]  ( .G(N618), .D(n182), .Q(\CACHE_mem[25][1] )
         );
  DLH_X1 \CACHE_mem_reg[25][0]  ( .G(N618), .D(n185), .Q(\CACHE_mem[25][0] )
         );
  DLH_X1 \CACHE_mem_reg[26][1]  ( .G(N617), .D(n182), .Q(\CACHE_mem[26][1] )
         );
  DLH_X1 \CACHE_mem_reg[26][0]  ( .G(N617), .D(n185), .Q(\CACHE_mem[26][0] )
         );
  DLH_X1 \CACHE_mem_reg[27][1]  ( .G(N616), .D(n182), .Q(\CACHE_mem[27][1] )
         );
  DLH_X1 \CACHE_mem_reg[27][0]  ( .G(N616), .D(n185), .Q(\CACHE_mem[27][0] )
         );
  DLH_X1 \CACHE_mem_reg[28][1]  ( .G(N615), .D(n182), .Q(\CACHE_mem[28][1] )
         );
  DLH_X1 \CACHE_mem_reg[28][0]  ( .G(N615), .D(n185), .Q(\CACHE_mem[28][0] )
         );
  DLH_X1 \CACHE_mem_reg[29][1]  ( .G(N614), .D(n182), .Q(\CACHE_mem[29][1] )
         );
  DLH_X1 \CACHE_mem_reg[29][0]  ( .G(N614), .D(n185), .Q(\CACHE_mem[29][0] )
         );
  DLH_X1 \CACHE_mem_reg[30][1]  ( .G(N613), .D(n182), .Q(\CACHE_mem[30][1] )
         );
  DLH_X1 \CACHE_mem_reg[30][0]  ( .G(N613), .D(n185), .Q(\CACHE_mem[30][0] )
         );
  DLH_X1 \CACHE_mem_reg[31][1]  ( .G(N612), .D(n182), .Q(\CACHE_mem[31][1] )
         );
  DLH_X1 \CACHE_mem_reg[31][0]  ( .G(N612), .D(n185), .Q(\CACHE_mem[31][0] )
         );
  NAND3_X1 U166 ( .A1(n233), .A2(n191), .A3(n69), .ZN(n60) );
  NAND3_X1 U167 ( .A1(n69), .A2(n191), .A3(PC_FAIL[5]), .ZN(n70) );
  NAND3_X1 U168 ( .A1(n69), .A2(n233), .A3(PC_FAIL[6]), .ZN(n71) );
  NAND3_X1 U169 ( .A1(n235), .A2(n234), .A3(n236), .ZN(n61) );
  NAND3_X1 U170 ( .A1(n235), .A2(n234), .A3(PC_FAIL[2]), .ZN(n62) );
  NAND3_X1 U171 ( .A1(n236), .A2(n234), .A3(PC_FAIL[3]), .ZN(n63) );
  NAND3_X1 U172 ( .A1(PC_FAIL[2]), .A2(n234), .A3(PC_FAIL[3]), .ZN(n64) );
  NAND3_X1 U173 ( .A1(n236), .A2(n235), .A3(PC_FAIL[4]), .ZN(n65) );
  NAND3_X1 U174 ( .A1(PC_FAIL[2]), .A2(n235), .A3(PC_FAIL[4]), .ZN(n66) );
  NAND3_X1 U175 ( .A1(PC_FAIL[3]), .A2(n236), .A3(PC_FAIL[4]), .ZN(n67) );
  NAND3_X1 U176 ( .A1(PC_FAIL[5]), .A2(n69), .A3(PC_FAIL[6]), .ZN(n72) );
  NAND3_X1 U177 ( .A1(PC_FAIL[3]), .A2(PC_FAIL[2]), .A3(PC_FAIL[4]), .ZN(n68)
         );
  NAND3_X1 U178 ( .A1(n109), .A2(n239), .A3(IR_IN[27]), .ZN(n108) );
  branch_predictor_DW01_add_0 add_65 ( .A(PC_IN), .B({IR_IN[15], IR_IN[15], 
        IR_IN[15], IR_IN[15], IR_IN[15], IR_IN[15], IR_IN[15], IR_IN[15], 
        IR_IN[15], IR_IN[15], IR_IN[15], IR_IN[15], IR_IN[15], IR_IN[15], 
        IR_IN[15], IR_IN[15], IR_IN[15:0]}), .CI(1'b0), .SUM({N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219}) );
  branch_predictor_DW01_add_1 add_60 ( .A(PC_IN), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N144, N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, 
        N116, N115, N114, N113}) );
  branch_predictor_DW01_add_2 add_59 ( .A(PC_IN), .B({IR_IN[25], IR_IN[25], 
        IR_IN[25], IR_IN[25], IR_IN[25], IR_IN[25], IR_IN[25:0]}), .CI(1'b0), 
        .SUM({N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81}) );
  branch_predictor_DW01_add_3 add_53_aco ( .A(PC_FAIL), .B({n5, n5, n5, n5, n5, 
        n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, n19, n18, n17, n16, 
        n15, n14, n13, n12, n11, n7, n10, n9, n8, n6, n20}), .CI(1'b0), .SUM({
        N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46}) );
  AND2_X1 U3 ( .A1(N116), .A2(n192), .ZN(N360) );
  AND2_X1 U4 ( .A1(N117), .A2(n193), .ZN(N361) );
  AND2_X1 U5 ( .A1(N118), .A2(n192), .ZN(N362) );
  AND2_X1 U6 ( .A1(N119), .A2(n195), .ZN(N363) );
  AND2_X1 U7 ( .A1(N120), .A2(n195), .ZN(N364) );
  AND2_X1 U8 ( .A1(N121), .A2(n195), .ZN(N365) );
  AND2_X1 U9 ( .A1(N122), .A2(n195), .ZN(N366) );
  AND2_X1 U14 ( .A1(N123), .A2(n195), .ZN(N367) );
  AND2_X1 U15 ( .A1(N124), .A2(n195), .ZN(N368) );
  AND2_X1 U16 ( .A1(N125), .A2(n195), .ZN(N369) );
  AND2_X1 U17 ( .A1(N126), .A2(n195), .ZN(N370) );
  AND2_X1 U18 ( .A1(N127), .A2(n194), .ZN(N371) );
  AND2_X1 U19 ( .A1(N128), .A2(n195), .ZN(N372) );
  AND2_X1 U20 ( .A1(N129), .A2(n195), .ZN(N373) );
  AND2_X1 U21 ( .A1(N130), .A2(n195), .ZN(N374) );
  AND2_X1 U22 ( .A1(N131), .A2(n195), .ZN(N375) );
  AND2_X1 U23 ( .A1(N132), .A2(n195), .ZN(N376) );
  AND2_X1 U24 ( .A1(N133), .A2(n195), .ZN(N377) );
  AND2_X1 U25 ( .A1(N134), .A2(n195), .ZN(N378) );
  AND2_X1 U26 ( .A1(N135), .A2(n195), .ZN(N379) );
  AND2_X1 U27 ( .A1(N136), .A2(n195), .ZN(N380) );
  AND2_X1 U28 ( .A1(N137), .A2(n195), .ZN(N381) );
  AND2_X1 U29 ( .A1(N138), .A2(n195), .ZN(N382) );
  AND2_X1 U30 ( .A1(N139), .A2(n195), .ZN(N383) );
  AND2_X1 U31 ( .A1(N140), .A2(n194), .ZN(N384) );
  AND2_X1 U32 ( .A1(N141), .A2(n194), .ZN(N385) );
  AND2_X1 U33 ( .A1(N142), .A2(n194), .ZN(N386) );
  AND2_X1 U34 ( .A1(N143), .A2(n194), .ZN(N387) );
  AND2_X1 U35 ( .A1(N144), .A2(n194), .ZN(N388) );
  AND2_X2 U36 ( .A1(IR_FAIL[15]), .A2(N479), .ZN(n5) );
  AND2_X1 U37 ( .A1(IR_FAIL[1]), .A2(N479), .ZN(n6) );
  BUF_X1 U38 ( .A(n231), .Z(n173) );
  BUF_X1 U39 ( .A(n231), .Z(n171) );
  BUF_X1 U40 ( .A(n231), .Z(n172) );
  BUF_X1 U41 ( .A(n75), .Z(n174) );
  BUF_X1 U42 ( .A(n75), .Z(n175) );
  BUF_X1 U43 ( .A(n75), .Z(n176) );
  INV_X1 U44 ( .A(n56), .ZN(n231) );
  BUF_X1 U45 ( .A(n53), .Z(n179) );
  NOR2_X1 U46 ( .A1(n197), .A2(WRONG_PRE), .ZN(n107) );
  INV_X1 U47 ( .A(n198), .ZN(n192) );
  INV_X1 U48 ( .A(n198), .ZN(n193) );
  INV_X1 U49 ( .A(n197), .ZN(n195) );
  INV_X1 U50 ( .A(n198), .ZN(n194) );
  BUF_X1 U51 ( .A(n53), .Z(n177) );
  BUF_X1 U52 ( .A(n53), .Z(n178) );
  OAI21_X1 U53 ( .B1(n60), .B2(n61), .A(n193), .ZN(N643) );
  BUF_X1 U54 ( .A(N356), .Z(n186) );
  NAND2_X1 U55 ( .A1(WRONG_PRE), .A2(n192), .ZN(n56) );
  BUF_X1 U56 ( .A(PC_FAIL[6]), .Z(n140) );
  BUF_X1 U57 ( .A(PC_FAIL[6]), .Z(n139) );
  OAI21_X1 U58 ( .B1(n61), .B2(n71), .A(n193), .ZN(N627) );
  BUF_X1 U59 ( .A(PC_FAIL[6]), .Z(n138) );
  BUF_X1 U60 ( .A(N323), .Z(n189) );
  BUF_X1 U61 ( .A(N323), .Z(n188) );
  BUF_X1 U62 ( .A(N644), .Z(n184) );
  BUF_X1 U63 ( .A(N644), .Z(n183) );
  BUF_X1 U64 ( .A(N645), .Z(n181) );
  BUF_X1 U65 ( .A(N645), .Z(n180) );
  BUF_X1 U66 ( .A(N323), .Z(n190) );
  AND2_X1 U67 ( .A1(n238), .A2(n107), .ZN(n75) );
  BUF_X1 U68 ( .A(N644), .Z(n185) );
  BUF_X1 U69 ( .A(N645), .Z(n182) );
  BUF_X1 U70 ( .A(N356), .Z(n187) );
  AND2_X1 U71 ( .A1(n107), .A2(n108), .ZN(n53) );
  AND2_X1 U72 ( .A1(n179), .A2(n54), .ZN(TAKEN) );
  OAI21_X1 U73 ( .B1(n60), .B2(n68), .A(n192), .ZN(N636) );
  OAI21_X1 U74 ( .B1(n60), .B2(n67), .A(n192), .ZN(N637) );
  OAI21_X1 U75 ( .B1(n60), .B2(n66), .A(n192), .ZN(N638) );
  OAI21_X1 U76 ( .B1(n60), .B2(n65), .A(n192), .ZN(N639) );
  OAI21_X1 U77 ( .B1(n60), .B2(n64), .A(n192), .ZN(N640) );
  OAI21_X1 U78 ( .B1(n60), .B2(n63), .A(n192), .ZN(N641) );
  OAI21_X1 U79 ( .B1(n60), .B2(n62), .A(n192), .ZN(N642) );
  OAI21_X1 U80 ( .B1(n68), .B2(n72), .A(n194), .ZN(N612) );
  OAI21_X1 U81 ( .B1(n67), .B2(n72), .A(n194), .ZN(N613) );
  OAI21_X1 U82 ( .B1(n66), .B2(n72), .A(n194), .ZN(N614) );
  OAI21_X1 U83 ( .B1(n65), .B2(n72), .A(n194), .ZN(N615) );
  OAI21_X1 U84 ( .B1(n64), .B2(n72), .A(n194), .ZN(N616) );
  OAI21_X1 U85 ( .B1(n63), .B2(n72), .A(n194), .ZN(N617) );
  OAI21_X1 U86 ( .B1(n62), .B2(n72), .A(n194), .ZN(N618) );
  OAI21_X1 U87 ( .B1(n61), .B2(n72), .A(n194), .ZN(N619) );
  OAI21_X1 U88 ( .B1(n68), .B2(n70), .A(n193), .ZN(N628) );
  OAI21_X1 U89 ( .B1(n67), .B2(n70), .A(n193), .ZN(N629) );
  OAI21_X1 U90 ( .B1(n66), .B2(n70), .A(n193), .ZN(N630) );
  OAI21_X1 U91 ( .B1(n65), .B2(n70), .A(n192), .ZN(N631) );
  OAI21_X1 U92 ( .B1(n64), .B2(n70), .A(n193), .ZN(N632) );
  OAI21_X1 U93 ( .B1(n63), .B2(n70), .A(n192), .ZN(N633) );
  OAI21_X1 U94 ( .B1(n62), .B2(n70), .A(n192), .ZN(N634) );
  OAI21_X1 U95 ( .B1(n61), .B2(n70), .A(n192), .ZN(N635) );
  OAI21_X1 U96 ( .B1(n68), .B2(n71), .A(n193), .ZN(N620) );
  OAI21_X1 U97 ( .B1(n67), .B2(n71), .A(n193), .ZN(N621) );
  OAI21_X1 U98 ( .B1(n66), .B2(n71), .A(n193), .ZN(N622) );
  OAI21_X1 U99 ( .B1(n65), .B2(n71), .A(n193), .ZN(N623) );
  OAI21_X1 U100 ( .B1(n64), .B2(n71), .A(n193), .ZN(N624) );
  OAI21_X1 U101 ( .B1(n63), .B2(n71), .A(n193), .ZN(N625) );
  OAI21_X1 U102 ( .B1(n62), .B2(n71), .A(n193), .ZN(N626) );
  OAI21_X1 U103 ( .B1(WRONG_PRE), .B2(n108), .A(n192), .ZN(N356) );
  INV_X1 U104 ( .A(N479), .ZN(n232) );
  NOR2_X1 U105 ( .A1(N480), .A2(n56), .ZN(N644) );
  NOR2_X1 U106 ( .A1(n57), .A2(n196), .ZN(N645) );
  AOI22_X1 U107 ( .A1(n173), .A2(n58), .B1(n59), .B2(n56), .ZN(n57) );
  OAI21_X1 U108 ( .B1(N480), .B2(n232), .A(n59), .ZN(n58) );
  NAND2_X1 U109 ( .A1(N480), .A2(n232), .ZN(n59) );
  NAND2_X1 U110 ( .A1(n56), .A2(n73), .ZN(n69) );
  NAND2_X1 U111 ( .A1(RIGHT_PRE), .A2(N480), .ZN(n73) );
  OAI21_X1 U112 ( .B1(n55), .B2(n196), .A(n56), .ZN(SEL) );
  NOR2_X1 U113 ( .A1(n238), .A2(n54), .ZN(n55) );
  INV_X1 U114 ( .A(n108), .ZN(n238) );
  OR3_X1 U115 ( .A1(n186), .A2(WRONG_PRE), .A3(n54), .ZN(N323) );
  INV_X1 U116 ( .A(n82), .ZN(n206) );
  AOI222_X1 U117 ( .A1(N70), .A2(n173), .B1(N105), .B2(n176), .C1(N243), .C2(
        n179), .ZN(n82) );
  INV_X1 U118 ( .A(n81), .ZN(n205) );
  AOI222_X1 U119 ( .A1(N71), .A2(n173), .B1(N106), .B2(n176), .C1(N244), .C2(
        n179), .ZN(n81) );
  INV_X1 U120 ( .A(n80), .ZN(n204) );
  AOI222_X1 U121 ( .A1(N72), .A2(n173), .B1(N107), .B2(n176), .C1(N245), .C2(
        n179), .ZN(n80) );
  INV_X1 U122 ( .A(n79), .ZN(n203) );
  AOI222_X1 U123 ( .A1(N73), .A2(n173), .B1(N108), .B2(n176), .C1(N246), .C2(
        n179), .ZN(n79) );
  INV_X1 U124 ( .A(n78), .ZN(n202) );
  AOI222_X1 U125 ( .A1(N74), .A2(n173), .B1(N109), .B2(n176), .C1(N247), .C2(
        n179), .ZN(n78) );
  INV_X1 U126 ( .A(n77), .ZN(n201) );
  AOI222_X1 U127 ( .A1(N75), .A2(n173), .B1(N110), .B2(n176), .C1(N248), .C2(
        n179), .ZN(n77) );
  INV_X1 U128 ( .A(n76), .ZN(n200) );
  AOI222_X1 U129 ( .A1(N76), .A2(n173), .B1(N111), .B2(n176), .C1(N249), .C2(
        n179), .ZN(n76) );
  INV_X1 U130 ( .A(n106), .ZN(n230) );
  AOI222_X1 U131 ( .A1(N46), .A2(n171), .B1(N81), .B2(n174), .C1(N219), .C2(
        n177), .ZN(n106) );
  INV_X1 U132 ( .A(n105), .ZN(n229) );
  AOI222_X1 U133 ( .A1(N47), .A2(n171), .B1(N82), .B2(n174), .C1(N220), .C2(
        n177), .ZN(n105) );
  INV_X1 U134 ( .A(n104), .ZN(n228) );
  AOI222_X1 U135 ( .A1(N48), .A2(n171), .B1(N83), .B2(n174), .C1(N221), .C2(
        n177), .ZN(n104) );
  INV_X1 U136 ( .A(n103), .ZN(n227) );
  AOI222_X1 U137 ( .A1(N49), .A2(n171), .B1(N84), .B2(n174), .C1(N222), .C2(
        n177), .ZN(n103) );
  INV_X1 U138 ( .A(n102), .ZN(n226) );
  AOI222_X1 U139 ( .A1(N50), .A2(n171), .B1(N85), .B2(n174), .C1(N223), .C2(
        n177), .ZN(n102) );
  INV_X1 U140 ( .A(n101), .ZN(n225) );
  AOI222_X1 U141 ( .A1(N51), .A2(n171), .B1(N86), .B2(n174), .C1(N224), .C2(
        n177), .ZN(n101) );
  INV_X1 U142 ( .A(n100), .ZN(n224) );
  AOI222_X1 U143 ( .A1(N52), .A2(n171), .B1(N87), .B2(n174), .C1(N225), .C2(
        n177), .ZN(n100) );
  INV_X1 U144 ( .A(n99), .ZN(n223) );
  AOI222_X1 U145 ( .A1(N53), .A2(n171), .B1(N88), .B2(n174), .C1(N226), .C2(
        n177), .ZN(n99) );
  INV_X1 U146 ( .A(n98), .ZN(n222) );
  AOI222_X1 U147 ( .A1(N54), .A2(n171), .B1(N89), .B2(n174), .C1(N227), .C2(
        n177), .ZN(n98) );
  INV_X1 U148 ( .A(n97), .ZN(n221) );
  AOI222_X1 U149 ( .A1(N55), .A2(n171), .B1(N90), .B2(n174), .C1(N228), .C2(
        n177), .ZN(n97) );
  INV_X1 U150 ( .A(n96), .ZN(n220) );
  AOI222_X1 U151 ( .A1(N56), .A2(n171), .B1(N91), .B2(n174), .C1(N229), .C2(
        n177), .ZN(n96) );
  INV_X1 U152 ( .A(n95), .ZN(n219) );
  AOI222_X1 U153 ( .A1(N57), .A2(n171), .B1(N92), .B2(n174), .C1(N230), .C2(
        n177), .ZN(n95) );
  INV_X1 U154 ( .A(n94), .ZN(n218) );
  AOI222_X1 U155 ( .A1(N58), .A2(n172), .B1(N93), .B2(n175), .C1(N231), .C2(
        n178), .ZN(n94) );
  INV_X1 U156 ( .A(n93), .ZN(n217) );
  AOI222_X1 U157 ( .A1(N59), .A2(n172), .B1(N94), .B2(n175), .C1(N232), .C2(
        n178), .ZN(n93) );
  INV_X1 U158 ( .A(n92), .ZN(n216) );
  AOI222_X1 U159 ( .A1(N60), .A2(n172), .B1(N95), .B2(n175), .C1(N233), .C2(
        n178), .ZN(n92) );
  INV_X1 U160 ( .A(n91), .ZN(n215) );
  AOI222_X1 U161 ( .A1(N61), .A2(n172), .B1(N96), .B2(n175), .C1(N234), .C2(
        n178), .ZN(n91) );
  INV_X1 U162 ( .A(n90), .ZN(n214) );
  AOI222_X1 U163 ( .A1(N62), .A2(n172), .B1(N97), .B2(n175), .C1(N235), .C2(
        n178), .ZN(n90) );
  INV_X1 U164 ( .A(n89), .ZN(n213) );
  AOI222_X1 U165 ( .A1(N63), .A2(n172), .B1(N98), .B2(n175), .C1(N236), .C2(
        n178), .ZN(n89) );
  INV_X1 U179 ( .A(n88), .ZN(n212) );
  AOI222_X1 U180 ( .A1(N64), .A2(n172), .B1(N99), .B2(n175), .C1(N237), .C2(
        n178), .ZN(n88) );
  INV_X1 U181 ( .A(n87), .ZN(n211) );
  AOI222_X1 U182 ( .A1(N65), .A2(n172), .B1(N100), .B2(n175), .C1(N238), .C2(
        n178), .ZN(n87) );
  INV_X1 U183 ( .A(n86), .ZN(n210) );
  AOI222_X1 U184 ( .A1(N66), .A2(n172), .B1(N101), .B2(n175), .C1(N239), .C2(
        n178), .ZN(n86) );
  INV_X1 U185 ( .A(n85), .ZN(n209) );
  AOI222_X1 U186 ( .A1(N67), .A2(n172), .B1(N102), .B2(n175), .C1(N240), .C2(
        n178), .ZN(n85) );
  INV_X1 U187 ( .A(n84), .ZN(n208) );
  AOI222_X1 U188 ( .A1(N68), .A2(n172), .B1(N103), .B2(n175), .C1(N241), .C2(
        n178), .ZN(n84) );
  INV_X1 U189 ( .A(n83), .ZN(n207) );
  AOI222_X1 U190 ( .A1(N69), .A2(n172), .B1(N104), .B2(n175), .C1(N242), .C2(
        n178), .ZN(n83) );
  NOR4_X1 U191 ( .A1(n237), .A2(n239), .A3(N216), .A4(IR_IN[27]), .ZN(n54) );
  INV_X1 U192 ( .A(n109), .ZN(n237) );
  NOR3_X1 U193 ( .A1(IR_IN[31]), .A2(IR_IN[30]), .A3(IR_IN[29]), .ZN(n109) );
  INV_X1 U194 ( .A(PC_FAIL[5]), .ZN(n233) );
  INV_X1 U195 ( .A(PC_FAIL[4]), .ZN(n234) );
  INV_X1 U196 ( .A(PC_FAIL[2]), .ZN(n236) );
  AND2_X1 U197 ( .A1(IR_FAIL[5]), .A2(N479), .ZN(n7) );
  AND2_X1 U198 ( .A1(IR_FAIL[2]), .A2(N479), .ZN(n8) );
  AND2_X1 U199 ( .A1(IR_FAIL[3]), .A2(N479), .ZN(n9) );
  AND2_X1 U200 ( .A1(IR_FAIL[4]), .A2(N479), .ZN(n10) );
  AND2_X1 U201 ( .A1(IR_FAIL[6]), .A2(N479), .ZN(n11) );
  AND2_X1 U202 ( .A1(IR_FAIL[7]), .A2(N479), .ZN(n12) );
  AND2_X1 U203 ( .A1(IR_FAIL[8]), .A2(N479), .ZN(n13) );
  AND2_X1 U204 ( .A1(N479), .A2(IR_FAIL[9]), .ZN(n14) );
  AND2_X1 U205 ( .A1(IR_FAIL[10]), .A2(N479), .ZN(n15) );
  AND2_X1 U206 ( .A1(IR_FAIL[11]), .A2(N479), .ZN(n16) );
  AND2_X1 U207 ( .A1(IR_FAIL[12]), .A2(N479), .ZN(n17) );
  AND2_X1 U208 ( .A1(IR_FAIL[13]), .A2(N479), .ZN(n18) );
  AND2_X1 U209 ( .A1(IR_FAIL[14]), .A2(N479), .ZN(n19) );
  INV_X1 U210 ( .A(PC_FAIL[3]), .ZN(n235) );
  AND2_X1 U211 ( .A1(IR_FAIL[0]), .A2(N479), .ZN(n20) );
  INV_X1 U212 ( .A(n74), .ZN(n199) );
  AOI222_X1 U213 ( .A1(N77), .A2(n173), .B1(N112), .B2(n176), .C1(N250), .C2(
        n179), .ZN(n74) );
  INV_X1 U214 ( .A(IR_IN[28]), .ZN(n239) );
  AND2_X1 U215 ( .A1(N114), .A2(n193), .ZN(N358) );
  AND2_X1 U216 ( .A1(N115), .A2(n193), .ZN(N359) );
  MUX2_X1 U217 ( .A(\CACHE_mem[15][0] ), .B(\CACHE_mem[31][0] ), .S(n138), .Z(
        n21) );
  MUX2_X1 U218 ( .A(\CACHE_mem[7][0] ), .B(\CACHE_mem[23][0] ), .S(n138), .Z(
        n22) );
  MUX2_X1 U219 ( .A(n22), .B(n21), .S(PC_FAIL[5]), .Z(n23) );
  MUX2_X1 U220 ( .A(\CACHE_mem[11][0] ), .B(\CACHE_mem[27][0] ), .S(n138), .Z(
        n24) );
  MUX2_X1 U221 ( .A(\CACHE_mem[3][0] ), .B(\CACHE_mem[19][0] ), .S(n138), .Z(
        n25) );
  MUX2_X1 U222 ( .A(n25), .B(n24), .S(PC_FAIL[5]), .Z(n26) );
  MUX2_X1 U223 ( .A(n26), .B(n23), .S(PC_FAIL[4]), .Z(n27) );
  MUX2_X1 U224 ( .A(\CACHE_mem[14][0] ), .B(\CACHE_mem[30][0] ), .S(n138), .Z(
        n28) );
  MUX2_X1 U225 ( .A(\CACHE_mem[6][0] ), .B(\CACHE_mem[22][0] ), .S(n138), .Z(
        n29) );
  MUX2_X1 U226 ( .A(n29), .B(n28), .S(PC_FAIL[5]), .Z(n30) );
  MUX2_X1 U227 ( .A(\CACHE_mem[10][0] ), .B(\CACHE_mem[26][0] ), .S(n138), .Z(
        n31) );
  MUX2_X1 U228 ( .A(\CACHE_mem[2][0] ), .B(\CACHE_mem[18][0] ), .S(n138), .Z(
        n32) );
  MUX2_X1 U229 ( .A(n32), .B(n31), .S(PC_FAIL[5]), .Z(n33) );
  MUX2_X1 U230 ( .A(n33), .B(n30), .S(PC_FAIL[4]), .Z(n34) );
  MUX2_X1 U231 ( .A(n34), .B(n27), .S(PC_FAIL[2]), .Z(n35) );
  MUX2_X1 U232 ( .A(\CACHE_mem[13][0] ), .B(\CACHE_mem[29][0] ), .S(n139), .Z(
        n36) );
  MUX2_X1 U233 ( .A(\CACHE_mem[5][0] ), .B(\CACHE_mem[21][0] ), .S(n139), .Z(
        n37) );
  MUX2_X1 U234 ( .A(n37), .B(n36), .S(PC_FAIL[5]), .Z(n38) );
  MUX2_X1 U235 ( .A(\CACHE_mem[9][0] ), .B(\CACHE_mem[25][0] ), .S(n139), .Z(
        n39) );
  MUX2_X1 U236 ( .A(\CACHE_mem[1][0] ), .B(\CACHE_mem[17][0] ), .S(n139), .Z(
        n40) );
  MUX2_X1 U237 ( .A(n40), .B(n39), .S(PC_FAIL[5]), .Z(n41) );
  MUX2_X1 U238 ( .A(n41), .B(n38), .S(PC_FAIL[4]), .Z(n42) );
  MUX2_X1 U239 ( .A(\CACHE_mem[12][0] ), .B(\CACHE_mem[28][0] ), .S(n139), .Z(
        n43) );
  MUX2_X1 U240 ( .A(\CACHE_mem[4][0] ), .B(\CACHE_mem[20][0] ), .S(n139), .Z(
        n44) );
  MUX2_X1 U241 ( .A(n44), .B(n43), .S(PC_FAIL[5]), .Z(n45) );
  MUX2_X1 U242 ( .A(\CACHE_mem[8][0] ), .B(\CACHE_mem[24][0] ), .S(n139), .Z(
        n46) );
  MUX2_X1 U243 ( .A(\CACHE_mem[0][0] ), .B(\CACHE_mem[16][0] ), .S(n139), .Z(
        n47) );
  MUX2_X1 U244 ( .A(n47), .B(n46), .S(PC_FAIL[5]), .Z(n48) );
  MUX2_X1 U245 ( .A(n48), .B(n45), .S(PC_FAIL[4]), .Z(n49) );
  MUX2_X1 U246 ( .A(n49), .B(n42), .S(PC_FAIL[2]), .Z(n50) );
  MUX2_X1 U247 ( .A(n50), .B(n35), .S(PC_FAIL[3]), .Z(N480) );
  MUX2_X1 U248 ( .A(\CACHE_mem[15][1] ), .B(\CACHE_mem[31][1] ), .S(n139), .Z(
        n51) );
  MUX2_X1 U249 ( .A(\CACHE_mem[7][1] ), .B(\CACHE_mem[23][1] ), .S(n139), .Z(
        n52) );
  MUX2_X1 U250 ( .A(n52), .B(n51), .S(PC_FAIL[5]), .Z(n110) );
  MUX2_X1 U251 ( .A(\CACHE_mem[11][1] ), .B(\CACHE_mem[27][1] ), .S(n139), .Z(
        n111) );
  MUX2_X1 U252 ( .A(\CACHE_mem[3][1] ), .B(\CACHE_mem[19][1] ), .S(n139), .Z(
        n112) );
  MUX2_X1 U253 ( .A(n112), .B(n111), .S(PC_FAIL[5]), .Z(n113) );
  MUX2_X1 U254 ( .A(n113), .B(n110), .S(PC_FAIL[4]), .Z(n114) );
  MUX2_X1 U255 ( .A(\CACHE_mem[14][1] ), .B(\CACHE_mem[30][1] ), .S(n140), .Z(
        n115) );
  MUX2_X1 U256 ( .A(\CACHE_mem[6][1] ), .B(\CACHE_mem[22][1] ), .S(n140), .Z(
        n116) );
  MUX2_X1 U257 ( .A(n116), .B(n115), .S(PC_FAIL[5]), .Z(n117) );
  MUX2_X1 U258 ( .A(\CACHE_mem[10][1] ), .B(\CACHE_mem[26][1] ), .S(n140), .Z(
        n118) );
  MUX2_X1 U259 ( .A(\CACHE_mem[2][1] ), .B(\CACHE_mem[18][1] ), .S(n140), .Z(
        n119) );
  MUX2_X1 U260 ( .A(n119), .B(n118), .S(PC_FAIL[5]), .Z(n120) );
  MUX2_X1 U261 ( .A(n120), .B(n117), .S(PC_FAIL[4]), .Z(n121) );
  MUX2_X1 U262 ( .A(n121), .B(n114), .S(PC_FAIL[2]), .Z(n122) );
  MUX2_X1 U263 ( .A(\CACHE_mem[13][1] ), .B(\CACHE_mem[29][1] ), .S(n140), .Z(
        n123) );
  MUX2_X1 U264 ( .A(\CACHE_mem[5][1] ), .B(\CACHE_mem[21][1] ), .S(n140), .Z(
        n124) );
  MUX2_X1 U265 ( .A(n124), .B(n123), .S(PC_FAIL[5]), .Z(n125) );
  MUX2_X1 U266 ( .A(\CACHE_mem[9][1] ), .B(\CACHE_mem[25][1] ), .S(n140), .Z(
        n126) );
  MUX2_X1 U267 ( .A(\CACHE_mem[1][1] ), .B(\CACHE_mem[17][1] ), .S(n140), .Z(
        n127) );
  MUX2_X1 U268 ( .A(n127), .B(n126), .S(PC_FAIL[5]), .Z(n128) );
  MUX2_X1 U269 ( .A(n128), .B(n125), .S(PC_FAIL[4]), .Z(n129) );
  MUX2_X1 U270 ( .A(\CACHE_mem[12][1] ), .B(\CACHE_mem[28][1] ), .S(n140), .Z(
        n130) );
  MUX2_X1 U271 ( .A(\CACHE_mem[4][1] ), .B(\CACHE_mem[20][1] ), .S(n140), .Z(
        n131) );
  MUX2_X1 U272 ( .A(n131), .B(n130), .S(PC_FAIL[5]), .Z(n132) );
  MUX2_X1 U273 ( .A(\CACHE_mem[8][1] ), .B(\CACHE_mem[24][1] ), .S(n140), .Z(
        n133) );
  MUX2_X1 U274 ( .A(\CACHE_mem[0][1] ), .B(\CACHE_mem[16][1] ), .S(n140), .Z(
        n134) );
  MUX2_X1 U275 ( .A(n134), .B(n133), .S(PC_FAIL[5]), .Z(n135) );
  MUX2_X1 U276 ( .A(n135), .B(n132), .S(PC_FAIL[4]), .Z(n136) );
  MUX2_X1 U277 ( .A(n136), .B(n129), .S(PC_FAIL[2]), .Z(n137) );
  MUX2_X1 U278 ( .A(n137), .B(n122), .S(PC_FAIL[3]), .Z(N479) );
  MUX2_X1 U279 ( .A(\CACHE_mem[15][1] ), .B(\CACHE_mem[31][1] ), .S(PC_IN[6]), 
        .Z(n141) );
  MUX2_X1 U280 ( .A(\CACHE_mem[7][1] ), .B(\CACHE_mem[23][1] ), .S(PC_IN[6]), 
        .Z(n142) );
  MUX2_X1 U281 ( .A(n142), .B(n141), .S(PC_IN[5]), .Z(n143) );
  MUX2_X1 U282 ( .A(\CACHE_mem[11][1] ), .B(\CACHE_mem[27][1] ), .S(PC_IN[6]), 
        .Z(n144) );
  MUX2_X1 U283 ( .A(\CACHE_mem[3][1] ), .B(\CACHE_mem[19][1] ), .S(PC_IN[6]), 
        .Z(n145) );
  MUX2_X1 U284 ( .A(n145), .B(n144), .S(PC_IN[5]), .Z(n146) );
  MUX2_X1 U285 ( .A(n146), .B(n143), .S(PC_IN[4]), .Z(n147) );
  MUX2_X1 U286 ( .A(\CACHE_mem[14][1] ), .B(\CACHE_mem[30][1] ), .S(PC_IN[6]), 
        .Z(n148) );
  MUX2_X1 U287 ( .A(\CACHE_mem[6][1] ), .B(\CACHE_mem[22][1] ), .S(PC_IN[6]), 
        .Z(n149) );
  MUX2_X1 U288 ( .A(n149), .B(n148), .S(PC_IN[5]), .Z(n150) );
  MUX2_X1 U289 ( .A(\CACHE_mem[10][1] ), .B(\CACHE_mem[26][1] ), .S(PC_IN[6]), 
        .Z(n151) );
  MUX2_X1 U290 ( .A(\CACHE_mem[2][1] ), .B(\CACHE_mem[18][1] ), .S(PC_IN[6]), 
        .Z(n152) );
  MUX2_X1 U291 ( .A(n152), .B(n151), .S(PC_IN[5]), .Z(n153) );
  MUX2_X1 U292 ( .A(n153), .B(n150), .S(PC_IN[4]), .Z(n154) );
  MUX2_X1 U293 ( .A(n154), .B(n147), .S(PC_IN[2]), .Z(n155) );
  MUX2_X1 U294 ( .A(\CACHE_mem[13][1] ), .B(\CACHE_mem[29][1] ), .S(PC_IN[6]), 
        .Z(n156) );
  MUX2_X1 U295 ( .A(\CACHE_mem[5][1] ), .B(\CACHE_mem[21][1] ), .S(PC_IN[6]), 
        .Z(n157) );
  MUX2_X1 U296 ( .A(n157), .B(n156), .S(PC_IN[5]), .Z(n158) );
  MUX2_X1 U297 ( .A(\CACHE_mem[9][1] ), .B(\CACHE_mem[25][1] ), .S(PC_IN[6]), 
        .Z(n159) );
  MUX2_X1 U298 ( .A(\CACHE_mem[1][1] ), .B(\CACHE_mem[17][1] ), .S(PC_IN[6]), 
        .Z(n160) );
  MUX2_X1 U299 ( .A(n160), .B(n159), .S(PC_IN[5]), .Z(n161) );
  MUX2_X1 U300 ( .A(n161), .B(n158), .S(PC_IN[4]), .Z(n162) );
  MUX2_X1 U301 ( .A(\CACHE_mem[12][1] ), .B(\CACHE_mem[28][1] ), .S(PC_IN[6]), 
        .Z(n163) );
  MUX2_X1 U302 ( .A(\CACHE_mem[4][1] ), .B(\CACHE_mem[20][1] ), .S(PC_IN[6]), 
        .Z(n164) );
  MUX2_X1 U303 ( .A(n164), .B(n163), .S(PC_IN[5]), .Z(n165) );
  MUX2_X1 U304 ( .A(\CACHE_mem[8][1] ), .B(\CACHE_mem[24][1] ), .S(PC_IN[6]), 
        .Z(n166) );
  MUX2_X1 U305 ( .A(\CACHE_mem[0][1] ), .B(\CACHE_mem[16][1] ), .S(PC_IN[6]), 
        .Z(n167) );
  MUX2_X1 U306 ( .A(n167), .B(n166), .S(PC_IN[5]), .Z(n168) );
  MUX2_X1 U307 ( .A(n168), .B(n165), .S(PC_IN[4]), .Z(n169) );
  MUX2_X1 U308 ( .A(n169), .B(n162), .S(PC_IN[2]), .Z(n170) );
  MUX2_X1 U309 ( .A(n170), .B(n155), .S(PC_IN[3]), .Z(N216) );
  AND2_X1 U310 ( .A1(N113), .A2(n194), .ZN(N357) );
  INV_X1 U311 ( .A(PC_FAIL[6]), .ZN(n191) );
  INV_X1 U312 ( .A(RST), .ZN(n196) );
  INV_X1 U313 ( .A(RST), .ZN(n197) );
  INV_X1 U314 ( .A(RST), .ZN(n198) );
endmodule


module MUX21_GENERIC_N32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106;

  BUF_X1 U1 ( .A(n10), .Z(n3) );
  BUF_X1 U2 ( .A(n10), .Z(n2) );
  BUF_X1 U3 ( .A(n10), .Z(n8) );
  BUF_X1 U4 ( .A(n8), .Z(n7) );
  BUF_X1 U5 ( .A(n9), .Z(n6) );
  BUF_X1 U6 ( .A(n3), .Z(n5) );
  BUF_X1 U7 ( .A(n10), .Z(n4) );
  BUF_X1 U8 ( .A(n10), .Z(n9) );
  INV_X1 U9 ( .A(n1), .ZN(n10) );
  BUF_X1 U10 ( .A(SEL), .Z(n1) );
  INV_X1 U11 ( .A(n97), .ZN(Y[2]) );
  AOI22_X1 U12 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n4), .ZN(n97) );
  INV_X1 U13 ( .A(n103), .ZN(Y[6]) );
  AOI22_X1 U14 ( .A1(A[6]), .A2(SEL), .B1(B[6]), .B2(n2), .ZN(n103) );
  INV_X1 U15 ( .A(n102), .ZN(Y[5]) );
  AOI22_X1 U16 ( .A1(A[5]), .A2(n1), .B1(B[5]), .B2(n3), .ZN(n102) );
  INV_X1 U17 ( .A(n101), .ZN(Y[4]) );
  AOI22_X1 U18 ( .A1(A[4]), .A2(SEL), .B1(B[4]), .B2(n3), .ZN(n101) );
  INV_X1 U19 ( .A(n106), .ZN(Y[9]) );
  AOI22_X1 U20 ( .A1(n1), .A2(A[9]), .B1(B[9]), .B2(n2), .ZN(n106) );
  INV_X1 U21 ( .A(n77), .ZN(Y[11]) );
  AOI22_X1 U22 ( .A1(A[11]), .A2(SEL), .B1(B[11]), .B2(n9), .ZN(n77) );
  INV_X1 U23 ( .A(n80), .ZN(Y[14]) );
  AOI22_X1 U24 ( .A1(A[14]), .A2(n1), .B1(B[14]), .B2(n8), .ZN(n80) );
  INV_X1 U25 ( .A(n83), .ZN(Y[17]) );
  AOI22_X1 U26 ( .A1(A[17]), .A2(SEL), .B1(B[17]), .B2(n7), .ZN(n83) );
  INV_X1 U27 ( .A(n89), .ZN(Y[22]) );
  AOI22_X1 U28 ( .A1(A[22]), .A2(n1), .B1(B[22]), .B2(n6), .ZN(n89) );
  INV_X1 U29 ( .A(n92), .ZN(Y[25]) );
  AOI22_X1 U30 ( .A1(A[25]), .A2(n1), .B1(B[25]), .B2(n5), .ZN(n92) );
  INV_X1 U31 ( .A(n95), .ZN(Y[28]) );
  AOI22_X1 U32 ( .A1(A[28]), .A2(n1), .B1(B[28]), .B2(n4), .ZN(n95) );
  INV_X1 U33 ( .A(n88), .ZN(Y[21]) );
  AOI22_X1 U34 ( .A1(A[21]), .A2(n1), .B1(B[21]), .B2(n6), .ZN(n88) );
  INV_X1 U35 ( .A(n79), .ZN(Y[13]) );
  AOI22_X1 U36 ( .A1(A[13]), .A2(n1), .B1(B[13]), .B2(n8), .ZN(n79) );
  INV_X1 U37 ( .A(n82), .ZN(Y[16]) );
  AOI22_X1 U38 ( .A1(A[16]), .A2(SEL), .B1(B[16]), .B2(n8), .ZN(n82) );
  INV_X1 U39 ( .A(n85), .ZN(Y[19]) );
  AOI22_X1 U40 ( .A1(A[19]), .A2(n1), .B1(B[19]), .B2(n7), .ZN(n85) );
  INV_X1 U41 ( .A(n91), .ZN(Y[24]) );
  AOI22_X1 U42 ( .A1(A[24]), .A2(n1), .B1(B[24]), .B2(n5), .ZN(n91) );
  INV_X1 U43 ( .A(n94), .ZN(Y[27]) );
  AOI22_X1 U44 ( .A1(A[27]), .A2(n1), .B1(B[27]), .B2(n5), .ZN(n94) );
  INV_X1 U45 ( .A(n98), .ZN(Y[30]) );
  AOI22_X1 U46 ( .A1(A[30]), .A2(n1), .B1(B[30]), .B2(n4), .ZN(n98) );
  INV_X1 U47 ( .A(n87), .ZN(Y[20]) );
  AOI22_X1 U48 ( .A1(A[20]), .A2(n1), .B1(B[20]), .B2(n6), .ZN(n87) );
  INV_X1 U49 ( .A(n76), .ZN(Y[10]) );
  AOI22_X1 U50 ( .A1(A[10]), .A2(SEL), .B1(B[10]), .B2(n9), .ZN(n76) );
  INV_X1 U51 ( .A(n78), .ZN(Y[12]) );
  AOI22_X1 U52 ( .A1(A[12]), .A2(n1), .B1(B[12]), .B2(n9), .ZN(n78) );
  INV_X1 U53 ( .A(n81), .ZN(Y[15]) );
  AOI22_X1 U54 ( .A1(A[15]), .A2(SEL), .B1(B[15]), .B2(n8), .ZN(n81) );
  INV_X1 U55 ( .A(n84), .ZN(Y[18]) );
  AOI22_X1 U56 ( .A1(A[18]), .A2(n1), .B1(B[18]), .B2(n7), .ZN(n84) );
  INV_X1 U57 ( .A(n90), .ZN(Y[23]) );
  AOI22_X1 U58 ( .A1(A[23]), .A2(n1), .B1(B[23]), .B2(n6), .ZN(n90) );
  INV_X1 U59 ( .A(n93), .ZN(Y[26]) );
  AOI22_X1 U60 ( .A1(A[26]), .A2(n1), .B1(B[26]), .B2(n5), .ZN(n93) );
  INV_X1 U61 ( .A(n96), .ZN(Y[29]) );
  AOI22_X1 U62 ( .A1(A[29]), .A2(n1), .B1(B[29]), .B2(n4), .ZN(n96) );
  INV_X1 U63 ( .A(n100), .ZN(Y[3]) );
  AOI22_X1 U64 ( .A1(A[3]), .A2(n1), .B1(B[3]), .B2(n3), .ZN(n100) );
  INV_X1 U65 ( .A(n104), .ZN(Y[7]) );
  AOI22_X1 U66 ( .A1(A[7]), .A2(SEL), .B1(B[7]), .B2(n2), .ZN(n104) );
  INV_X1 U67 ( .A(n105), .ZN(Y[8]) );
  AOI22_X1 U68 ( .A1(A[8]), .A2(n1), .B1(B[8]), .B2(n2), .ZN(n105) );
  INV_X1 U69 ( .A(n99), .ZN(Y[31]) );
  AOI22_X1 U70 ( .A1(A[31]), .A2(SEL), .B1(B[31]), .B2(n3), .ZN(n99) );
  INV_X1 U71 ( .A(n75), .ZN(Y[0]) );
  INV_X1 U72 ( .A(n86), .ZN(Y[1]) );
  AOI22_X1 U73 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n86) );
  AOI22_X1 U74 ( .A1(A[0]), .A2(n1), .B1(B[0]), .B2(n9), .ZN(n75) );
endmodule


module NPC_adder_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X1 U1 ( .A1(A[6]), .A2(n2), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[5]), .A2(n3), .ZN(n2) );
  AND2_X1 U3 ( .A1(A[4]), .A2(n25), .ZN(n3) );
  AND2_X1 U4 ( .A1(A[9]), .A2(n27), .ZN(n4) );
  AND2_X1 U5 ( .A1(A[11]), .A2(n15), .ZN(n5) );
  AND2_X1 U6 ( .A1(A[14]), .A2(n12), .ZN(n6) );
  AND2_X1 U7 ( .A1(A[17]), .A2(n13), .ZN(n7) );
  AND2_X1 U8 ( .A1(A[22]), .A2(n11), .ZN(n8) );
  AND2_X1 U9 ( .A1(A[25]), .A2(n17), .ZN(n9) );
  AND2_X1 U10 ( .A1(A[28]), .A2(n18), .ZN(n10) );
  AND2_X1 U11 ( .A1(A[21]), .A2(n16), .ZN(n11) );
  AND2_X1 U12 ( .A1(A[13]), .A2(n19), .ZN(n12) );
  AND2_X1 U13 ( .A1(A[16]), .A2(n20), .ZN(n13) );
  AND2_X1 U14 ( .A1(A[19]), .A2(n21), .ZN(n14) );
  AND2_X1 U15 ( .A1(A[10]), .A2(n4), .ZN(n15) );
  AND2_X1 U16 ( .A1(A[20]), .A2(n14), .ZN(n16) );
  AND2_X1 U17 ( .A1(A[24]), .A2(n22), .ZN(n17) );
  AND2_X1 U18 ( .A1(A[27]), .A2(n23), .ZN(n18) );
  AND2_X1 U19 ( .A1(A[12]), .A2(n5), .ZN(n19) );
  AND2_X1 U20 ( .A1(A[15]), .A2(n6), .ZN(n20) );
  AND2_X1 U21 ( .A1(A[18]), .A2(n7), .ZN(n21) );
  AND2_X1 U22 ( .A1(A[23]), .A2(n8), .ZN(n22) );
  AND2_X1 U23 ( .A1(A[26]), .A2(n9), .ZN(n23) );
  AND2_X1 U24 ( .A1(A[29]), .A2(n10), .ZN(n24) );
  AND2_X1 U25 ( .A1(A[3]), .A2(A[2]), .ZN(n25) );
  AND2_X1 U26 ( .A1(A[7]), .A2(n1), .ZN(n26) );
  AND2_X1 U27 ( .A1(A[8]), .A2(n26), .ZN(n27) );
  INV_X1 U28 ( .A(A[2]), .ZN(SUM[2]) );
  XOR2_X1 U29 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U30 ( .A(A[7]), .B(n1), .Z(SUM[7]) );
  XOR2_X1 U31 ( .A(A[6]), .B(n2), .Z(SUM[6]) );
  XOR2_X1 U32 ( .A(A[5]), .B(n3), .Z(SUM[5]) );
  XOR2_X1 U33 ( .A(A[4]), .B(n25), .Z(SUM[4]) );
  XOR2_X1 U34 ( .A(A[10]), .B(n4), .Z(SUM[10]) );
  XOR2_X1 U35 ( .A(A[11]), .B(n15), .Z(SUM[11]) );
  XOR2_X1 U36 ( .A(A[12]), .B(n5), .Z(SUM[12]) );
  XOR2_X1 U37 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  XOR2_X1 U38 ( .A(A[14]), .B(n12), .Z(SUM[14]) );
  XOR2_X1 U39 ( .A(A[15]), .B(n6), .Z(SUM[15]) );
  XOR2_X1 U40 ( .A(A[16]), .B(n20), .Z(SUM[16]) );
  XOR2_X1 U41 ( .A(A[17]), .B(n13), .Z(SUM[17]) );
  XOR2_X1 U42 ( .A(A[18]), .B(n7), .Z(SUM[18]) );
  XOR2_X1 U43 ( .A(A[19]), .B(n21), .Z(SUM[19]) );
  XOR2_X1 U44 ( .A(A[20]), .B(n14), .Z(SUM[20]) );
  XOR2_X1 U45 ( .A(A[21]), .B(n16), .Z(SUM[21]) );
  XOR2_X1 U46 ( .A(A[22]), .B(n11), .Z(SUM[22]) );
  XOR2_X1 U47 ( .A(A[23]), .B(n8), .Z(SUM[23]) );
  XOR2_X1 U48 ( .A(A[24]), .B(n22), .Z(SUM[24]) );
  XOR2_X1 U49 ( .A(A[25]), .B(n17), .Z(SUM[25]) );
  XOR2_X1 U50 ( .A(A[26]), .B(n9), .Z(SUM[26]) );
  XOR2_X1 U51 ( .A(A[27]), .B(n23), .Z(SUM[27]) );
  XOR2_X1 U52 ( .A(A[28]), .B(n18), .Z(SUM[28]) );
  XOR2_X1 U53 ( .A(A[29]), .B(n10), .Z(SUM[29]) );
  XOR2_X1 U54 ( .A(A[30]), .B(n24), .Z(SUM[30]) );
  XOR2_X1 U55 ( .A(A[8]), .B(n26), .Z(SUM[8]) );
  XOR2_X1 U56 ( .A(A[9]), .B(n27), .Z(SUM[9]) );
  XNOR2_X1 U57 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  NAND2_X1 U58 ( .A1(A[30]), .A2(n24), .ZN(n57) );
endmodule


module NPC_adder ( inPC, outPC );
  input [31:0] inPC;
  output [31:0] outPC;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17;

  DLH_X1 \outPC_reg[31]  ( .G(n4), .D(N32), .Q(outPC[31]) );
  DLH_X1 \outPC_reg[30]  ( .G(n4), .D(N31), .Q(outPC[30]) );
  DLH_X1 \outPC_reg[29]  ( .G(n4), .D(N30), .Q(outPC[29]) );
  DLH_X1 \outPC_reg[28]  ( .G(n4), .D(N29), .Q(outPC[28]) );
  DLH_X1 \outPC_reg[27]  ( .G(n4), .D(N28), .Q(outPC[27]) );
  DLH_X1 \outPC_reg[26]  ( .G(n4), .D(N27), .Q(outPC[26]) );
  DLH_X1 \outPC_reg[25]  ( .G(n4), .D(N26), .Q(outPC[25]) );
  DLH_X1 \outPC_reg[24]  ( .G(n4), .D(N25), .Q(outPC[24]) );
  DLH_X1 \outPC_reg[23]  ( .G(n4), .D(N24), .Q(outPC[23]) );
  DLH_X1 \outPC_reg[22]  ( .G(n4), .D(N23), .Q(outPC[22]) );
  DLH_X1 \outPC_reg[21]  ( .G(n3), .D(N22), .Q(outPC[21]) );
  DLH_X1 \outPC_reg[20]  ( .G(n3), .D(N21), .Q(outPC[20]) );
  DLH_X1 \outPC_reg[19]  ( .G(n3), .D(N20), .Q(outPC[19]) );
  DLH_X1 \outPC_reg[18]  ( .G(n3), .D(N19), .Q(outPC[18]) );
  DLH_X1 \outPC_reg[17]  ( .G(n3), .D(N18), .Q(outPC[17]) );
  DLH_X1 \outPC_reg[16]  ( .G(n3), .D(N17), .Q(outPC[16]) );
  DLH_X1 \outPC_reg[15]  ( .G(n3), .D(N16), .Q(outPC[15]) );
  DLH_X1 \outPC_reg[14]  ( .G(n3), .D(N15), .Q(outPC[14]) );
  DLH_X1 \outPC_reg[13]  ( .G(n3), .D(N14), .Q(outPC[13]) );
  DLH_X1 \outPC_reg[12]  ( .G(n3), .D(N13), .Q(outPC[12]) );
  DLH_X1 \outPC_reg[11]  ( .G(n3), .D(N12), .Q(outPC[11]) );
  DLH_X1 \outPC_reg[10]  ( .G(n2), .D(N11), .Q(outPC[10]) );
  DLH_X1 \outPC_reg[9]  ( .G(n2), .D(N10), .Q(outPC[9]) );
  DLH_X1 \outPC_reg[8]  ( .G(n2), .D(N9), .Q(outPC[8]) );
  DLH_X1 \outPC_reg[7]  ( .G(n2), .D(N8), .Q(outPC[7]) );
  DLH_X1 \outPC_reg[6]  ( .G(n2), .D(N7), .Q(outPC[6]) );
  DLH_X1 \outPC_reg[5]  ( .G(n2), .D(N6), .Q(outPC[5]) );
  DLH_X1 \outPC_reg[4]  ( .G(n2), .D(N5), .Q(outPC[4]) );
  DLH_X1 \outPC_reg[3]  ( .G(n2), .D(N4), .Q(outPC[3]) );
  DLH_X1 \outPC_reg[2]  ( .G(n2), .D(N3), .Q(outPC[2]) );
  DLH_X1 \outPC_reg[1]  ( .G(n2), .D(N2), .Q(outPC[1]) );
  DLH_X1 \outPC_reg[0]  ( .G(n2), .D(N1), .Q(outPC[0]) );
  NPC_adder_DW01_add_0 add_40 ( .A(inPC), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  BUF_X1 U4 ( .A(N0), .Z(n2) );
  BUF_X1 U5 ( .A(N0), .Z(n3) );
  BUF_X1 U6 ( .A(N0), .Z(n4) );
  INV_X1 U7 ( .A(inPC[31]), .ZN(n17) );
  NOR2_X1 U8 ( .A1(inPC[21]), .A2(inPC[20]), .ZN(n8) );
  NOR3_X1 U9 ( .A1(inPC[22]), .A2(inPC[24]), .A3(inPC[23]), .ZN(n7) );
  NOR3_X1 U10 ( .A1(inPC[25]), .A2(inPC[27]), .A3(inPC[26]), .ZN(n6) );
  NOR3_X1 U11 ( .A1(inPC[28]), .A2(inPC[30]), .A3(inPC[29]), .ZN(n5) );
  NAND4_X1 U12 ( .A1(n8), .A2(n7), .A3(n6), .A4(n5), .ZN(n16) );
  AND4_X1 U13 ( .A1(inPC[9]), .A2(inPC[8]), .A3(inPC[7]), .A4(inPC[6]), .ZN(
        n10) );
  AND4_X1 U14 ( .A1(inPC[5]), .A2(inPC[4]), .A3(inPC[3]), .A4(inPC[2]), .ZN(n9) );
  AOI21_X1 U15 ( .B1(n10), .B2(n9), .A(inPC[10]), .ZN(n14) );
  NOR3_X1 U16 ( .A1(inPC[11]), .A2(inPC[13]), .A3(inPC[12]), .ZN(n13) );
  NOR3_X1 U17 ( .A1(inPC[14]), .A2(inPC[16]), .A3(inPC[15]), .ZN(n12) );
  NOR3_X1 U18 ( .A1(inPC[17]), .A2(inPC[19]), .A3(inPC[18]), .ZN(n11) );
  NAND4_X1 U19 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(n15) );
  OAI21_X1 U20 ( .B1(n16), .B2(n15), .A(n17), .ZN(N0) );
endmodule


module SNPS_CLOCK_GATE_HIGH_IF_ID ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module IF_ID ( CLK, RST, DISCARD, NPC_IN, NPC_L_IN, IR_IN, PR_IN, NPC_OUT, 
        NPC_L_OUT, IR_OUT, PR_OUT );
  input [31:0] NPC_IN;
  input [31:0] NPC_L_IN;
  input [31:0] IR_IN;
  output [31:0] NPC_OUT;
  output [31:0] NPC_L_OUT;
  output [31:0] IR_OUT;
  input CLK, RST, DISCARD, PR_IN;
  output PR_OUT;
  wire   net1013, n99, n101, n103, n105, n107, n109, n111, n113, n115, n117,
         n119, n121, n123, n125, n127, n129, n131, n133, n135, n137, n139,
         n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, n161,
         n163, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n100, n102, n104, n106, n108, n110, n112, n114, n116, n118, n120,
         n122, n124, n126, n128, n130;

  DFFR_X1 PR_OUT_reg ( .D(PR_IN), .CK(net1013), .RN(n47), .Q(PR_OUT) );
  DFFR_X1 \IR_OUT_reg[31]  ( .D(IR_IN[31]), .CK(CLK), .RN(n35), .Q(IR_OUT[31])
         );
  DFFS_X1 \IR_OUT_reg[30]  ( .D(IR_IN[30]), .CK(CLK), .SN(n36), .Q(IR_OUT[30])
         );
  DFFR_X1 \IR_OUT_reg[29]  ( .D(IR_IN[29]), .CK(CLK), .RN(n34), .Q(IR_OUT[29])
         );
  DFFS_X1 \IR_OUT_reg[28]  ( .D(IR_IN[28]), .CK(CLK), .SN(n36), .Q(IR_OUT[28])
         );
  DFFR_X1 \IR_OUT_reg[27]  ( .D(IR_IN[27]), .CK(CLK), .RN(n34), .Q(IR_OUT[27])
         );
  DFFS_X1 \IR_OUT_reg[26]  ( .D(IR_IN[26]), .CK(CLK), .SN(n36), .Q(IR_OUT[26])
         );
  DFFR_X1 \IR_OUT_reg[25]  ( .D(IR_IN[25]), .CK(CLK), .RN(n34), .Q(IR_OUT[25])
         );
  DFFR_X1 \IR_OUT_reg[24]  ( .D(IR_IN[24]), .CK(CLK), .RN(n34), .Q(IR_OUT[24])
         );
  DFFR_X1 \IR_OUT_reg[23]  ( .D(IR_IN[23]), .CK(CLK), .RN(n34), .Q(IR_OUT[23])
         );
  DFFR_X1 \IR_OUT_reg[22]  ( .D(IR_IN[22]), .CK(CLK), .RN(n34), .Q(IR_OUT[22])
         );
  DFFR_X1 \IR_OUT_reg[21]  ( .D(IR_IN[21]), .CK(CLK), .RN(n34), .Q(IR_OUT[21])
         );
  DFFR_X1 \IR_OUT_reg[20]  ( .D(IR_IN[20]), .CK(CLK), .RN(n34), .Q(IR_OUT[20])
         );
  DFFR_X1 \IR_OUT_reg[19]  ( .D(IR_IN[19]), .CK(CLK), .RN(n34), .Q(IR_OUT[19])
         );
  DFFR_X1 \IR_OUT_reg[18]  ( .D(IR_IN[18]), .CK(CLK), .RN(n34), .Q(IR_OUT[18])
         );
  DFFR_X1 \IR_OUT_reg[17]  ( .D(IR_IN[17]), .CK(CLK), .RN(n34), .Q(IR_OUT[17])
         );
  DFFR_X1 \IR_OUT_reg[16]  ( .D(IR_IN[16]), .CK(CLK), .RN(n35), .Q(IR_OUT[16])
         );
  DFFR_X1 \IR_OUT_reg[15]  ( .D(IR_IN[15]), .CK(CLK), .RN(n35), .Q(IR_OUT[15])
         );
  DFFR_X1 \IR_OUT_reg[14]  ( .D(IR_IN[14]), .CK(CLK), .RN(n35), .Q(IR_OUT[14])
         );
  DFFR_X1 \IR_OUT_reg[13]  ( .D(IR_IN[13]), .CK(CLK), .RN(n35), .Q(IR_OUT[13])
         );
  DFFR_X1 \IR_OUT_reg[12]  ( .D(IR_IN[12]), .CK(CLK), .RN(n35), .Q(IR_OUT[12])
         );
  DFFR_X1 \IR_OUT_reg[11]  ( .D(IR_IN[11]), .CK(CLK), .RN(n35), .Q(IR_OUT[11])
         );
  DFFR_X1 \IR_OUT_reg[10]  ( .D(IR_IN[10]), .CK(CLK), .RN(n35), .Q(IR_OUT[10])
         );
  DFFR_X1 \IR_OUT_reg[9]  ( .D(IR_IN[9]), .CK(CLK), .RN(n35), .Q(IR_OUT[9]) );
  DFFR_X1 \IR_OUT_reg[8]  ( .D(IR_IN[8]), .CK(CLK), .RN(n35), .Q(IR_OUT[8]) );
  DFFR_X1 \IR_OUT_reg[7]  ( .D(IR_IN[7]), .CK(CLK), .RN(n35), .Q(IR_OUT[7]) );
  DFFR_X1 \IR_OUT_reg[6]  ( .D(IR_IN[6]), .CK(CLK), .RN(n35), .Q(IR_OUT[6]) );
  DFFR_X1 \IR_OUT_reg[5]  ( .D(IR_IN[5]), .CK(CLK), .RN(n36), .Q(IR_OUT[5]) );
  DFFR_X1 \IR_OUT_reg[4]  ( .D(IR_IN[4]), .CK(CLK), .RN(n36), .Q(IR_OUT[4]) );
  DFFR_X1 \IR_OUT_reg[3]  ( .D(IR_IN[3]), .CK(CLK), .RN(n36), .Q(IR_OUT[3]) );
  DFFR_X1 \IR_OUT_reg[2]  ( .D(IR_IN[2]), .CK(CLK), .RN(n36), .Q(IR_OUT[2]) );
  DFFR_X1 \IR_OUT_reg[1]  ( .D(IR_IN[1]), .CK(CLK), .RN(n36), .Q(IR_OUT[1]) );
  DFFR_X1 \IR_OUT_reg[0]  ( .D(IR_IN[0]), .CK(CLK), .RN(n34), .Q(IR_OUT[0]) );
  DFFR_X1 \NPC_L_OUT_reg[31]  ( .D(NPC_L_IN[31]), .CK(net1013), .RN(n47), .Q(
        NPC_L_OUT[31]) );
  DFFR_X1 \NPC_L_OUT_reg[30]  ( .D(NPC_L_IN[30]), .CK(net1013), .RN(n47), .Q(
        NPC_L_OUT[30]) );
  DFFR_X1 \NPC_L_OUT_reg[29]  ( .D(NPC_L_IN[29]), .CK(net1013), .RN(n47), .Q(
        NPC_L_OUT[29]) );
  DFFR_X1 \NPC_L_OUT_reg[28]  ( .D(NPC_L_IN[28]), .CK(net1013), .RN(n47), .Q(
        NPC_L_OUT[28]) );
  DFFR_X1 \NPC_L_OUT_reg[27]  ( .D(NPC_L_IN[27]), .CK(net1013), .RN(n47), .Q(
        NPC_L_OUT[27]) );
  DFFR_X1 \NPC_L_OUT_reg[26]  ( .D(NPC_L_IN[26]), .CK(net1013), .RN(n47), .Q(
        NPC_L_OUT[26]) );
  DFFR_X1 \NPC_L_OUT_reg[25]  ( .D(NPC_L_IN[25]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[25]) );
  DFFR_X1 \NPC_L_OUT_reg[24]  ( .D(NPC_L_IN[24]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[24]) );
  DFFR_X1 \NPC_L_OUT_reg[23]  ( .D(NPC_L_IN[23]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[23]) );
  DFFR_X1 \NPC_L_OUT_reg[22]  ( .D(NPC_L_IN[22]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[22]) );
  DFFR_X1 \NPC_L_OUT_reg[21]  ( .D(NPC_L_IN[21]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[21]) );
  DFFR_X1 \NPC_L_OUT_reg[20]  ( .D(NPC_L_IN[20]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[20]) );
  DFFR_X1 \NPC_L_OUT_reg[19]  ( .D(NPC_L_IN[19]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[19]) );
  DFFR_X1 \NPC_L_OUT_reg[18]  ( .D(NPC_L_IN[18]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[18]) );
  DFFR_X1 \NPC_L_OUT_reg[17]  ( .D(NPC_L_IN[17]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[17]) );
  DFFR_X1 \NPC_L_OUT_reg[16]  ( .D(NPC_L_IN[16]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[16]) );
  DFFR_X1 \NPC_L_OUT_reg[15]  ( .D(NPC_L_IN[15]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[15]) );
  DFFR_X1 \NPC_L_OUT_reg[14]  ( .D(NPC_L_IN[14]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[14]) );
  DFFR_X1 \NPC_L_OUT_reg[13]  ( .D(NPC_L_IN[13]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[13]) );
  DFFR_X1 \NPC_L_OUT_reg[12]  ( .D(NPC_L_IN[12]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[12]) );
  DFFR_X1 \NPC_L_OUT_reg[11]  ( .D(NPC_L_IN[11]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[11]) );
  DFFR_X1 \NPC_L_OUT_reg[10]  ( .D(NPC_L_IN[10]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[10]) );
  DFFR_X1 \NPC_L_OUT_reg[9]  ( .D(NPC_L_IN[9]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[9]) );
  DFFR_X1 \NPC_L_OUT_reg[8]  ( .D(NPC_L_IN[8]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[8]) );
  DFFR_X1 \NPC_L_OUT_reg[7]  ( .D(NPC_L_IN[7]), .CK(net1013), .RN(n48), .Q(
        NPC_L_OUT[7]) );
  DFFR_X1 \NPC_L_OUT_reg[6]  ( .D(NPC_L_IN[6]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[6]) );
  DFFR_X1 \NPC_L_OUT_reg[5]  ( .D(NPC_L_IN[5]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[5]) );
  DFFR_X1 \NPC_L_OUT_reg[4]  ( .D(NPC_L_IN[4]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[4]) );
  DFFR_X1 \NPC_L_OUT_reg[3]  ( .D(NPC_L_IN[3]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[3]) );
  DFFR_X1 \NPC_L_OUT_reg[2]  ( .D(NPC_L_IN[2]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[2]) );
  DFFR_X1 \NPC_L_OUT_reg[1]  ( .D(NPC_L_IN[1]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[1]) );
  DFFR_X1 \NPC_L_OUT_reg[0]  ( .D(NPC_L_IN[0]), .CK(net1013), .RN(n49), .Q(
        NPC_L_OUT[0]) );
  SNPS_CLOCK_GATE_HIGH_IF_ID clk_gate_PR_OUT_reg ( .CLK(CLK), .EN(n39), 
        .ENCLK(net1013), .TE(1'b0) );
  DFFRS_X1 \NPC_OUT_reg[31]  ( .D(NPC_IN[31]), .CK(CLK), .RN(n73), .SN(n25), 
        .Q(NPC_OUT[31]) );
  DFFRS_X1 \NPC_OUT_reg[30]  ( .D(NPC_IN[30]), .CK(CLK), .RN(n72), .SN(n24), 
        .Q(NPC_OUT[30]) );
  DFFRS_X1 \NPC_OUT_reg[29]  ( .D(NPC_IN[29]), .CK(CLK), .RN(n71), .SN(n23), 
        .Q(NPC_OUT[29]) );
  DFFRS_X1 \NPC_OUT_reg[28]  ( .D(NPC_IN[28]), .CK(CLK), .RN(n70), .SN(n22), 
        .Q(NPC_OUT[28]) );
  DFFRS_X1 \NPC_OUT_reg[27]  ( .D(NPC_IN[27]), .CK(CLK), .RN(n69), .SN(n21), 
        .Q(NPC_OUT[27]) );
  DFFRS_X1 \NPC_OUT_reg[26]  ( .D(NPC_IN[26]), .CK(CLK), .RN(n68), .SN(n20), 
        .Q(NPC_OUT[26]) );
  DFFRS_X1 \NPC_OUT_reg[25]  ( .D(NPC_IN[25]), .CK(CLK), .RN(n67), .SN(n19), 
        .Q(NPC_OUT[25]) );
  DFFRS_X1 \NPC_OUT_reg[24]  ( .D(NPC_IN[24]), .CK(CLK), .RN(n66), .SN(n18), 
        .Q(NPC_OUT[24]) );
  DFFRS_X1 \NPC_OUT_reg[23]  ( .D(NPC_IN[23]), .CK(CLK), .RN(n65), .SN(n17), 
        .Q(NPC_OUT[23]) );
  DFFRS_X1 \NPC_OUT_reg[22]  ( .D(NPC_IN[22]), .CK(CLK), .RN(n64), .SN(n16), 
        .Q(NPC_OUT[22]) );
  DFFRS_X1 \NPC_OUT_reg[21]  ( .D(NPC_IN[21]), .CK(CLK), .RN(n63), .SN(n15), 
        .Q(NPC_OUT[21]) );
  DFFRS_X1 \NPC_OUT_reg[20]  ( .D(NPC_IN[20]), .CK(CLK), .RN(n62), .SN(n14), 
        .Q(NPC_OUT[20]) );
  DFFRS_X1 \NPC_OUT_reg[19]  ( .D(NPC_IN[19]), .CK(CLK), .RN(n61), .SN(n13), 
        .Q(NPC_OUT[19]) );
  DFFRS_X1 \NPC_OUT_reg[18]  ( .D(NPC_IN[18]), .CK(CLK), .RN(n60), .SN(n12), 
        .Q(NPC_OUT[18]) );
  DFFRS_X1 \NPC_OUT_reg[17]  ( .D(NPC_IN[17]), .CK(CLK), .RN(n59), .SN(n11), 
        .Q(NPC_OUT[17]) );
  DFFRS_X1 \NPC_OUT_reg[16]  ( .D(NPC_IN[16]), .CK(CLK), .RN(n58), .SN(n33), 
        .Q(NPC_OUT[16]) );
  DFFRS_X1 \NPC_OUT_reg[15]  ( .D(NPC_IN[15]), .CK(CLK), .RN(n57), .SN(n32), 
        .Q(NPC_OUT[15]) );
  DFFRS_X1 \NPC_OUT_reg[14]  ( .D(NPC_IN[14]), .CK(CLK), .RN(n56), .SN(n31), 
        .Q(NPC_OUT[14]) );
  DFFRS_X1 \NPC_OUT_reg[13]  ( .D(NPC_IN[13]), .CK(CLK), .RN(n55), .SN(n30), 
        .Q(NPC_OUT[13]) );
  DFFRS_X1 \NPC_OUT_reg[12]  ( .D(NPC_IN[12]), .CK(CLK), .RN(n54), .SN(n29), 
        .Q(NPC_OUT[12]) );
  DFFRS_X1 \NPC_OUT_reg[11]  ( .D(NPC_IN[11]), .CK(CLK), .RN(n53), .SN(n28), 
        .Q(NPC_OUT[11]) );
  DFFRS_X1 \NPC_OUT_reg[10]  ( .D(NPC_IN[10]), .CK(CLK), .RN(n52), .SN(n27), 
        .Q(NPC_OUT[10]) );
  DFFRS_X1 \NPC_OUT_reg[9]  ( .D(NPC_IN[9]), .CK(CLK), .RN(n51), .SN(n26), .Q(
        NPC_OUT[9]) );
  DFFRS_X1 \NPC_OUT_reg[8]  ( .D(NPC_IN[8]), .CK(CLK), .RN(n50), .SN(n10), .Q(
        NPC_OUT[8]) );
  DFFRS_X1 \NPC_OUT_reg[7]  ( .D(NPC_IN[7]), .CK(CLK), .RN(n81), .SN(n9), .Q(
        NPC_OUT[7]) );
  DFFRS_X1 \NPC_OUT_reg[6]  ( .D(NPC_IN[6]), .CK(CLK), .RN(n80), .SN(n8), .Q(
        NPC_OUT[6]) );
  DFFRS_X1 \NPC_OUT_reg[5]  ( .D(NPC_IN[5]), .CK(CLK), .RN(n79), .SN(n7), .Q(
        NPC_OUT[5]) );
  DFFRS_X1 \NPC_OUT_reg[4]  ( .D(NPC_IN[4]), .CK(CLK), .RN(n78), .SN(n6), .Q(
        NPC_OUT[4]) );
  DFFRS_X1 \NPC_OUT_reg[3]  ( .D(NPC_IN[3]), .CK(CLK), .RN(n77), .SN(n5), .Q(
        NPC_OUT[3]) );
  DFFRS_X1 \NPC_OUT_reg[2]  ( .D(NPC_IN[2]), .CK(CLK), .RN(n76), .SN(n4), .Q(
        NPC_OUT[2]) );
  DFFRS_X1 \NPC_OUT_reg[1]  ( .D(NPC_IN[1]), .CK(CLK), .RN(n75), .SN(n3), .Q(
        NPC_OUT[1]) );
  DFFRS_X1 \NPC_OUT_reg[0]  ( .D(NPC_IN[0]), .CK(CLK), .RN(n74), .SN(n2), .Q(
        NPC_OUT[0]) );
  INV_X1 U3 ( .A(NPC_IN[0]), .ZN(n130) );
  INV_X1 U4 ( .A(NPC_IN[1]), .ZN(n128) );
  INV_X1 U5 ( .A(NPC_IN[2]), .ZN(n126) );
  INV_X1 U6 ( .A(NPC_IN[3]), .ZN(n124) );
  INV_X1 U7 ( .A(NPC_IN[4]), .ZN(n122) );
  INV_X1 U8 ( .A(NPC_IN[5]), .ZN(n120) );
  INV_X1 U9 ( .A(NPC_IN[6]), .ZN(n118) );
  INV_X1 U10 ( .A(NPC_IN[7]), .ZN(n116) );
  INV_X1 U11 ( .A(NPC_IN[8]), .ZN(n114) );
  INV_X1 U12 ( .A(NPC_IN[9]), .ZN(n112) );
  INV_X1 U13 ( .A(NPC_IN[10]), .ZN(n110) );
  INV_X1 U14 ( .A(NPC_IN[11]), .ZN(n108) );
  INV_X1 U15 ( .A(NPC_IN[12]), .ZN(n106) );
  INV_X1 U16 ( .A(NPC_IN[13]), .ZN(n104) );
  INV_X1 U17 ( .A(NPC_IN[14]), .ZN(n102) );
  INV_X1 U18 ( .A(NPC_IN[15]), .ZN(n100) );
  INV_X1 U19 ( .A(NPC_IN[16]), .ZN(n98) );
  INV_X1 U20 ( .A(NPC_IN[17]), .ZN(n97) );
  INV_X1 U21 ( .A(NPC_IN[18]), .ZN(n96) );
  INV_X1 U22 ( .A(NPC_IN[19]), .ZN(n95) );
  INV_X1 U23 ( .A(NPC_IN[20]), .ZN(n94) );
  INV_X1 U24 ( .A(NPC_IN[21]), .ZN(n93) );
  INV_X1 U25 ( .A(NPC_IN[22]), .ZN(n92) );
  INV_X1 U26 ( .A(NPC_IN[23]), .ZN(n91) );
  INV_X1 U27 ( .A(NPC_IN[24]), .ZN(n90) );
  INV_X1 U28 ( .A(NPC_IN[25]), .ZN(n89) );
  INV_X1 U29 ( .A(NPC_IN[26]), .ZN(n88) );
  INV_X1 U30 ( .A(NPC_IN[27]), .ZN(n87) );
  INV_X1 U31 ( .A(NPC_IN[28]), .ZN(n86) );
  INV_X1 U32 ( .A(NPC_IN[29]), .ZN(n85) );
  INV_X1 U33 ( .A(NPC_IN[30]), .ZN(n84) );
  INV_X1 U34 ( .A(NPC_IN[31]), .ZN(n83) );
  BUF_X1 U35 ( .A(n1), .Z(n34) );
  BUF_X1 U36 ( .A(n1), .Z(n35) );
  BUF_X1 U37 ( .A(n1), .Z(n36) );
  BUF_X1 U38 ( .A(n82), .Z(n39) );
  BUF_X1 U39 ( .A(n82), .Z(n37) );
  BUF_X1 U40 ( .A(n82), .Z(n38) );
  BUF_X1 U41 ( .A(n99), .Z(n41) );
  BUF_X1 U42 ( .A(n99), .Z(n40) );
  BUF_X1 U43 ( .A(n99), .Z(n42) );
  AND2_X1 U44 ( .A1(n47), .A2(n37), .ZN(n1) );
  INV_X1 U45 ( .A(DISCARD), .ZN(n82) );
  BUF_X1 U46 ( .A(n44), .Z(n48) );
  BUF_X1 U47 ( .A(n43), .Z(n45) );
  BUF_X1 U48 ( .A(n43), .Z(n46) );
  BUF_X1 U49 ( .A(n43), .Z(n47) );
  NAND2_X1 U50 ( .A1(DISCARD), .A2(n45), .ZN(n99) );
  BUF_X1 U51 ( .A(n44), .Z(n49) );
  BUF_X1 U52 ( .A(RST), .Z(n43) );
  BUF_X1 U53 ( .A(RST), .Z(n44) );
  INV_X1 U54 ( .A(n101), .ZN(n74) );
  OAI21_X1 U55 ( .B1(NPC_IN[0]), .B2(n39), .A(n46), .ZN(n101) );
  INV_X1 U56 ( .A(n103), .ZN(n75) );
  OAI21_X1 U57 ( .B1(NPC_IN[1]), .B2(n39), .A(n46), .ZN(n103) );
  INV_X1 U58 ( .A(n105), .ZN(n76) );
  OAI21_X1 U59 ( .B1(NPC_IN[2]), .B2(n39), .A(n47), .ZN(n105) );
  INV_X1 U60 ( .A(n107), .ZN(n77) );
  OAI21_X1 U61 ( .B1(NPC_IN[3]), .B2(n39), .A(n47), .ZN(n107) );
  INV_X1 U62 ( .A(n109), .ZN(n78) );
  OAI21_X1 U63 ( .B1(NPC_IN[4]), .B2(n39), .A(n47), .ZN(n109) );
  INV_X1 U64 ( .A(n111), .ZN(n79) );
  OAI21_X1 U65 ( .B1(NPC_IN[5]), .B2(n39), .A(n47), .ZN(n111) );
  INV_X1 U66 ( .A(n113), .ZN(n80) );
  OAI21_X1 U67 ( .B1(NPC_IN[6]), .B2(n39), .A(n47), .ZN(n113) );
  INV_X1 U68 ( .A(n115), .ZN(n81) );
  OAI21_X1 U69 ( .B1(NPC_IN[7]), .B2(n39), .A(n47), .ZN(n115) );
  INV_X1 U70 ( .A(n163), .ZN(n73) );
  OAI21_X1 U71 ( .B1(NPC_IN[31]), .B2(n39), .A(n46), .ZN(n163) );
  INV_X1 U72 ( .A(n119), .ZN(n51) );
  OAI21_X1 U73 ( .B1(NPC_IN[9]), .B2(n37), .A(n45), .ZN(n119) );
  INV_X1 U74 ( .A(n121), .ZN(n52) );
  OAI21_X1 U75 ( .B1(NPC_IN[10]), .B2(n37), .A(n45), .ZN(n121) );
  INV_X1 U76 ( .A(n123), .ZN(n53) );
  OAI21_X1 U77 ( .B1(NPC_IN[11]), .B2(n37), .A(n45), .ZN(n123) );
  INV_X1 U78 ( .A(n125), .ZN(n54) );
  OAI21_X1 U79 ( .B1(NPC_IN[12]), .B2(n37), .A(n45), .ZN(n125) );
  INV_X1 U80 ( .A(n127), .ZN(n55) );
  OAI21_X1 U81 ( .B1(NPC_IN[13]), .B2(n37), .A(n45), .ZN(n127) );
  INV_X1 U82 ( .A(n129), .ZN(n56) );
  OAI21_X1 U83 ( .B1(NPC_IN[14]), .B2(n37), .A(n45), .ZN(n129) );
  INV_X1 U84 ( .A(n131), .ZN(n57) );
  OAI21_X1 U85 ( .B1(NPC_IN[15]), .B2(n37), .A(n45), .ZN(n131) );
  INV_X1 U86 ( .A(n133), .ZN(n58) );
  OAI21_X1 U87 ( .B1(NPC_IN[16]), .B2(n37), .A(n45), .ZN(n133) );
  INV_X1 U88 ( .A(n135), .ZN(n59) );
  OAI21_X1 U89 ( .B1(NPC_IN[17]), .B2(n37), .A(n45), .ZN(n135) );
  INV_X1 U90 ( .A(n137), .ZN(n60) );
  OAI21_X1 U91 ( .B1(NPC_IN[18]), .B2(n37), .A(n45), .ZN(n137) );
  INV_X1 U92 ( .A(n139), .ZN(n61) );
  OAI21_X1 U93 ( .B1(NPC_IN[19]), .B2(n37), .A(n45), .ZN(n139) );
  INV_X1 U94 ( .A(n117), .ZN(n50) );
  OAI21_X1 U95 ( .B1(NPC_IN[8]), .B2(n38), .A(n47), .ZN(n117) );
  INV_X1 U96 ( .A(n141), .ZN(n62) );
  OAI21_X1 U97 ( .B1(NPC_IN[20]), .B2(n38), .A(n45), .ZN(n141) );
  INV_X1 U98 ( .A(n143), .ZN(n63) );
  OAI21_X1 U99 ( .B1(NPC_IN[21]), .B2(n38), .A(n46), .ZN(n143) );
  INV_X1 U100 ( .A(n145), .ZN(n64) );
  OAI21_X1 U101 ( .B1(NPC_IN[22]), .B2(n38), .A(n46), .ZN(n145) );
  INV_X1 U102 ( .A(n147), .ZN(n65) );
  OAI21_X1 U103 ( .B1(NPC_IN[23]), .B2(n38), .A(n46), .ZN(n147) );
  INV_X1 U104 ( .A(n149), .ZN(n66) );
  OAI21_X1 U105 ( .B1(NPC_IN[24]), .B2(n38), .A(n46), .ZN(n149) );
  INV_X1 U106 ( .A(n151), .ZN(n67) );
  OAI21_X1 U107 ( .B1(NPC_IN[25]), .B2(n38), .A(n46), .ZN(n151) );
  INV_X1 U108 ( .A(n153), .ZN(n68) );
  OAI21_X1 U109 ( .B1(NPC_IN[26]), .B2(n38), .A(n46), .ZN(n153) );
  INV_X1 U110 ( .A(n155), .ZN(n69) );
  OAI21_X1 U111 ( .B1(NPC_IN[27]), .B2(n38), .A(n46), .ZN(n155) );
  INV_X1 U112 ( .A(n157), .ZN(n70) );
  OAI21_X1 U113 ( .B1(NPC_IN[28]), .B2(n38), .A(n46), .ZN(n157) );
  INV_X1 U114 ( .A(n159), .ZN(n71) );
  OAI21_X1 U115 ( .B1(NPC_IN[29]), .B2(n38), .A(n46), .ZN(n159) );
  INV_X1 U116 ( .A(n161), .ZN(n72) );
  OAI21_X1 U117 ( .B1(NPC_IN[30]), .B2(n38), .A(n46), .ZN(n161) );
  OR2_X1 U118 ( .A1(n40), .A2(n130), .ZN(n2) );
  OR2_X1 U119 ( .A1(n40), .A2(n128), .ZN(n3) );
  OR2_X1 U120 ( .A1(n40), .A2(n126), .ZN(n4) );
  OR2_X1 U121 ( .A1(n40), .A2(n124), .ZN(n5) );
  OR2_X1 U122 ( .A1(n40), .A2(n122), .ZN(n6) );
  OR2_X1 U123 ( .A1(n40), .A2(n120), .ZN(n7) );
  OR2_X1 U124 ( .A1(n40), .A2(n118), .ZN(n8) );
  OR2_X1 U125 ( .A1(n40), .A2(n116), .ZN(n9) );
  OR2_X1 U126 ( .A1(n40), .A2(n114), .ZN(n10) );
  OR2_X1 U127 ( .A1(n41), .A2(n97), .ZN(n11) );
  OR2_X1 U128 ( .A1(n41), .A2(n96), .ZN(n12) );
  OR2_X1 U129 ( .A1(n41), .A2(n95), .ZN(n13) );
  OR2_X1 U130 ( .A1(n41), .A2(n94), .ZN(n14) );
  OR2_X1 U131 ( .A1(n41), .A2(n93), .ZN(n15) );
  OR2_X1 U132 ( .A1(n41), .A2(n92), .ZN(n16) );
  OR2_X1 U133 ( .A1(n41), .A2(n91), .ZN(n17) );
  OR2_X1 U134 ( .A1(n41), .A2(n90), .ZN(n18) );
  OR2_X1 U135 ( .A1(n41), .A2(n89), .ZN(n19) );
  OR2_X1 U136 ( .A1(n41), .A2(n88), .ZN(n20) );
  OR2_X1 U137 ( .A1(n41), .A2(n87), .ZN(n21) );
  OR2_X1 U138 ( .A1(n41), .A2(n86), .ZN(n22) );
  OR2_X1 U139 ( .A1(n40), .A2(n85), .ZN(n23) );
  OR2_X1 U140 ( .A1(n40), .A2(n84), .ZN(n24) );
  OR2_X1 U141 ( .A1(n40), .A2(n83), .ZN(n25) );
  OR2_X1 U142 ( .A1(n42), .A2(n112), .ZN(n26) );
  OR2_X1 U143 ( .A1(n42), .A2(n110), .ZN(n27) );
  OR2_X1 U144 ( .A1(n42), .A2(n108), .ZN(n28) );
  OR2_X1 U145 ( .A1(n42), .A2(n106), .ZN(n29) );
  OR2_X1 U146 ( .A1(n42), .A2(n104), .ZN(n30) );
  OR2_X1 U147 ( .A1(n42), .A2(n102), .ZN(n31) );
  OR2_X1 U148 ( .A1(n42), .A2(n100), .ZN(n32) );
  OR2_X1 U149 ( .A1(n42), .A2(n98), .ZN(n33) );
endmodule


module IR_decoder ( rst, IR_OUT, ADDS1, ADDS2, ADDD );
  input [20:0] IR_OUT;
  output [4:0] ADDS1;
  output [4:0] ADDS2;
  output [4:0] ADDD;
  input rst;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n34;

  NAND3_X1 U50 ( .A1(n5), .A2(n4), .A3(n6), .ZN(n28) );
  AOI211_X1 U3 ( .C1(n13), .C2(n14), .A(n9), .B(n2), .ZN(ADDS2[4]) );
  AND2_X1 U4 ( .A1(n15), .A2(n16), .ZN(n13) );
  NOR2_X1 U5 ( .A1(n17), .A2(n34), .ZN(ADDS2[0]) );
  NOR2_X1 U6 ( .A1(n17), .A2(n11), .ZN(ADDS2[2]) );
  NOR2_X1 U7 ( .A1(n17), .A2(n12), .ZN(ADDS2[1]) );
  NOR2_X1 U8 ( .A1(n17), .A2(n10), .ZN(ADDS2[3]) );
  OAI21_X1 U9 ( .B1(n3), .B2(n18), .A(n1), .ZN(n17) );
  NAND2_X1 U10 ( .A1(n16), .A2(n15), .ZN(n18) );
  INV_X1 U11 ( .A(n14), .ZN(n3) );
  NOR2_X1 U12 ( .A1(n16), .A2(n2), .ZN(n23) );
  NAND2_X1 U13 ( .A1(n1), .A2(n19), .ZN(n22) );
  INV_X1 U14 ( .A(rst), .ZN(n2) );
  NAND4_X1 U15 ( .A1(IR_OUT[20]), .A2(IR_OUT[18]), .A3(n30), .A4(n31), .ZN(n15) );
  NOR2_X1 U16 ( .A1(IR_OUT[19]), .A2(IR_OUT[17]), .ZN(n30) );
  NOR3_X1 U17 ( .A1(n28), .A2(n7), .A3(n8), .ZN(n19) );
  INV_X1 U18 ( .A(IR_OUT[16]), .ZN(n7) );
  NAND2_X1 U19 ( .A1(IR_OUT[16]), .A2(n8), .ZN(n31) );
  NAND2_X1 U20 ( .A1(IR_OUT[19]), .A2(n19), .ZN(n14) );
  INV_X1 U21 ( .A(IR_OUT[17]), .ZN(n6) );
  INV_X1 U22 ( .A(IR_OUT[18]), .ZN(n5) );
  OR4_X1 U23 ( .A1(n28), .A2(IR_OUT[15]), .A3(IR_OUT[16]), .A4(IR_OUT[19]), 
        .ZN(n16) );
  INV_X1 U24 ( .A(IR_OUT[20]), .ZN(n4) );
  AND2_X1 U25 ( .A1(IR_OUT[10]), .A2(n1), .ZN(ADDS1[0]) );
  AND2_X1 U26 ( .A1(IR_OUT[14]), .A2(n1), .ZN(ADDS1[4]) );
  AND2_X1 U27 ( .A1(IR_OUT[12]), .A2(n1), .ZN(ADDS1[2]) );
  AND2_X1 U28 ( .A1(IR_OUT[11]), .A2(n1), .ZN(ADDS1[1]) );
  INV_X1 U29 ( .A(IR_OUT[15]), .ZN(n8) );
  AND2_X1 U30 ( .A1(IR_OUT[13]), .A2(n1), .ZN(ADDS1[3]) );
  INV_X1 U31 ( .A(IR_OUT[5]), .ZN(n34) );
  INV_X1 U32 ( .A(IR_OUT[6]), .ZN(n12) );
  INV_X1 U33 ( .A(IR_OUT[7]), .ZN(n11) );
  INV_X1 U34 ( .A(IR_OUT[8]), .ZN(n10) );
  INV_X1 U35 ( .A(IR_OUT[9]), .ZN(n9) );
  NAND4_X1 U36 ( .A1(n1), .A2(n16), .A3(n29), .A4(n15), .ZN(n20) );
  OAI211_X1 U37 ( .C1(n32), .C2(n33), .A(n5), .B(n4), .ZN(n29) );
  NOR2_X1 U38 ( .A1(IR_OUT[17]), .A2(n31), .ZN(n33) );
  NOR3_X1 U39 ( .A1(n6), .A2(IR_OUT[19]), .A3(IR_OUT[16]), .ZN(n32) );
  OAI211_X1 U40 ( .C1(n34), .C2(n20), .A(n27), .B(n22), .ZN(ADDD[0]) );
  NAND2_X1 U41 ( .A1(IR_OUT[0]), .A2(n23), .ZN(n27) );
  OAI211_X1 U42 ( .C1(n12), .C2(n20), .A(n26), .B(n22), .ZN(ADDD[1]) );
  NAND2_X1 U43 ( .A1(IR_OUT[1]), .A2(n23), .ZN(n26) );
  OAI211_X1 U44 ( .C1(n11), .C2(n20), .A(n25), .B(n22), .ZN(ADDD[2]) );
  NAND2_X1 U45 ( .A1(IR_OUT[2]), .A2(n23), .ZN(n25) );
  OAI211_X1 U46 ( .C1(n10), .C2(n20), .A(n24), .B(n22), .ZN(ADDD[3]) );
  NAND2_X1 U47 ( .A1(IR_OUT[3]), .A2(n23), .ZN(n24) );
  OAI211_X1 U48 ( .C1(n9), .C2(n20), .A(n21), .B(n22), .ZN(ADDD[4]) );
  NAND2_X1 U49 ( .A1(IR_OUT[4]), .A2(n23), .ZN(n21) );
  INV_X1 U51 ( .A(n2), .ZN(n1) );
endmodule


module register_file_N32_addBit5 ( RESET, RE, WE, ADD_WR, ADD_RDA, ADD_RDB, 
        DATAIN, OUTA, OUTB );
  input [4:0] ADD_WR;
  input [4:0] ADD_RDA;
  input [4:0] ADD_RDB;
  input [31:0] DATAIN;
  output [31:0] OUTA;
  output [31:0] OUTB;
  input RESET, RE, WE;
  wire   \REGISTERS[1][31] , \REGISTERS[1][30] , \REGISTERS[1][29] ,
         \REGISTERS[1][28] , \REGISTERS[1][27] , \REGISTERS[1][26] ,
         \REGISTERS[1][25] , \REGISTERS[1][24] , \REGISTERS[1][23] ,
         \REGISTERS[1][22] , \REGISTERS[1][21] , \REGISTERS[1][20] ,
         \REGISTERS[1][19] , \REGISTERS[1][18] , \REGISTERS[1][17] ,
         \REGISTERS[1][16] , \REGISTERS[1][15] , \REGISTERS[1][14] ,
         \REGISTERS[1][13] , \REGISTERS[1][12] , \REGISTERS[1][11] ,
         \REGISTERS[1][10] , \REGISTERS[1][9] , \REGISTERS[1][8] ,
         \REGISTERS[1][7] , \REGISTERS[1][6] , \REGISTERS[1][5] ,
         \REGISTERS[1][4] , \REGISTERS[1][3] , \REGISTERS[1][2] ,
         \REGISTERS[1][1] , \REGISTERS[1][0] , \REGISTERS[2][31] ,
         \REGISTERS[2][30] , \REGISTERS[2][29] , \REGISTERS[2][28] ,
         \REGISTERS[2][27] , \REGISTERS[2][26] , \REGISTERS[2][25] ,
         \REGISTERS[2][24] , \REGISTERS[2][23] , \REGISTERS[2][22] ,
         \REGISTERS[2][21] , \REGISTERS[2][20] , \REGISTERS[2][19] ,
         \REGISTERS[2][18] , \REGISTERS[2][17] , \REGISTERS[2][16] ,
         \REGISTERS[2][15] , \REGISTERS[2][14] , \REGISTERS[2][13] ,
         \REGISTERS[2][12] , \REGISTERS[2][11] , \REGISTERS[2][10] ,
         \REGISTERS[2][9] , \REGISTERS[2][8] , \REGISTERS[2][7] ,
         \REGISTERS[2][6] , \REGISTERS[2][5] , \REGISTERS[2][4] ,
         \REGISTERS[2][3] , \REGISTERS[2][2] , \REGISTERS[2][1] ,
         \REGISTERS[2][0] , \REGISTERS[3][31] , \REGISTERS[3][30] ,
         \REGISTERS[3][29] , \REGISTERS[3][28] , \REGISTERS[3][27] ,
         \REGISTERS[3][26] , \REGISTERS[3][25] , \REGISTERS[3][24] ,
         \REGISTERS[3][23] , \REGISTERS[3][22] , \REGISTERS[3][21] ,
         \REGISTERS[3][20] , \REGISTERS[3][19] , \REGISTERS[3][18] ,
         \REGISTERS[3][17] , \REGISTERS[3][16] , \REGISTERS[3][15] ,
         \REGISTERS[3][14] , \REGISTERS[3][13] , \REGISTERS[3][12] ,
         \REGISTERS[3][11] , \REGISTERS[3][10] , \REGISTERS[3][9] ,
         \REGISTERS[3][8] , \REGISTERS[3][7] , \REGISTERS[3][6] ,
         \REGISTERS[3][5] , \REGISTERS[3][4] , \REGISTERS[3][3] ,
         \REGISTERS[3][2] , \REGISTERS[3][1] , \REGISTERS[3][0] ,
         \REGISTERS[4][31] , \REGISTERS[4][30] , \REGISTERS[4][29] ,
         \REGISTERS[4][28] , \REGISTERS[4][27] , \REGISTERS[4][26] ,
         \REGISTERS[4][25] , \REGISTERS[4][24] , \REGISTERS[4][23] ,
         \REGISTERS[4][22] , \REGISTERS[4][21] , \REGISTERS[4][20] ,
         \REGISTERS[4][19] , \REGISTERS[4][18] , \REGISTERS[4][17] ,
         \REGISTERS[4][16] , \REGISTERS[4][15] , \REGISTERS[4][14] ,
         \REGISTERS[4][13] , \REGISTERS[4][12] , \REGISTERS[4][11] ,
         \REGISTERS[4][10] , \REGISTERS[4][9] , \REGISTERS[4][8] ,
         \REGISTERS[4][7] , \REGISTERS[4][6] , \REGISTERS[4][5] ,
         \REGISTERS[4][4] , \REGISTERS[4][3] , \REGISTERS[4][2] ,
         \REGISTERS[4][1] , \REGISTERS[4][0] , \REGISTERS[5][31] ,
         \REGISTERS[5][30] , \REGISTERS[5][29] , \REGISTERS[5][28] ,
         \REGISTERS[5][27] , \REGISTERS[5][26] , \REGISTERS[5][25] ,
         \REGISTERS[5][24] , \REGISTERS[5][23] , \REGISTERS[5][22] ,
         \REGISTERS[5][21] , \REGISTERS[5][20] , \REGISTERS[5][19] ,
         \REGISTERS[5][18] , \REGISTERS[5][17] , \REGISTERS[5][16] ,
         \REGISTERS[5][15] , \REGISTERS[5][14] , \REGISTERS[5][13] ,
         \REGISTERS[5][12] , \REGISTERS[5][11] , \REGISTERS[5][10] ,
         \REGISTERS[5][9] , \REGISTERS[5][8] , \REGISTERS[5][7] ,
         \REGISTERS[5][6] , \REGISTERS[5][5] , \REGISTERS[5][4] ,
         \REGISTERS[5][3] , \REGISTERS[5][2] , \REGISTERS[5][1] ,
         \REGISTERS[5][0] , \REGISTERS[6][31] , \REGISTERS[6][30] ,
         \REGISTERS[6][29] , \REGISTERS[6][28] , \REGISTERS[6][27] ,
         \REGISTERS[6][26] , \REGISTERS[6][25] , \REGISTERS[6][24] ,
         \REGISTERS[6][23] , \REGISTERS[6][22] , \REGISTERS[6][21] ,
         \REGISTERS[6][20] , \REGISTERS[6][19] , \REGISTERS[6][18] ,
         \REGISTERS[6][17] , \REGISTERS[6][16] , \REGISTERS[6][15] ,
         \REGISTERS[6][14] , \REGISTERS[6][13] , \REGISTERS[6][12] ,
         \REGISTERS[6][11] , \REGISTERS[6][10] , \REGISTERS[6][9] ,
         \REGISTERS[6][8] , \REGISTERS[6][7] , \REGISTERS[6][6] ,
         \REGISTERS[6][5] , \REGISTERS[6][4] , \REGISTERS[6][3] ,
         \REGISTERS[6][2] , \REGISTERS[6][1] , \REGISTERS[6][0] ,
         \REGISTERS[7][31] , \REGISTERS[7][30] , \REGISTERS[7][29] ,
         \REGISTERS[7][28] , \REGISTERS[7][27] , \REGISTERS[7][26] ,
         \REGISTERS[7][25] , \REGISTERS[7][24] , \REGISTERS[7][23] ,
         \REGISTERS[7][22] , \REGISTERS[7][21] , \REGISTERS[7][20] ,
         \REGISTERS[7][19] , \REGISTERS[7][18] , \REGISTERS[7][17] ,
         \REGISTERS[7][16] , \REGISTERS[7][15] , \REGISTERS[7][14] ,
         \REGISTERS[7][13] , \REGISTERS[7][12] , \REGISTERS[7][11] ,
         \REGISTERS[7][10] , \REGISTERS[7][9] , \REGISTERS[7][8] ,
         \REGISTERS[7][7] , \REGISTERS[7][6] , \REGISTERS[7][5] ,
         \REGISTERS[7][4] , \REGISTERS[7][3] , \REGISTERS[7][2] ,
         \REGISTERS[7][1] , \REGISTERS[7][0] , \REGISTERS[8][31] ,
         \REGISTERS[8][30] , \REGISTERS[8][29] , \REGISTERS[8][28] ,
         \REGISTERS[8][27] , \REGISTERS[8][26] , \REGISTERS[8][25] ,
         \REGISTERS[8][24] , \REGISTERS[8][23] , \REGISTERS[8][22] ,
         \REGISTERS[8][21] , \REGISTERS[8][20] , \REGISTERS[8][19] ,
         \REGISTERS[8][18] , \REGISTERS[8][17] , \REGISTERS[8][16] ,
         \REGISTERS[8][15] , \REGISTERS[8][14] , \REGISTERS[8][13] ,
         \REGISTERS[8][12] , \REGISTERS[8][11] , \REGISTERS[8][10] ,
         \REGISTERS[8][9] , \REGISTERS[8][8] , \REGISTERS[8][7] ,
         \REGISTERS[8][6] , \REGISTERS[8][5] , \REGISTERS[8][4] ,
         \REGISTERS[8][3] , \REGISTERS[8][2] , \REGISTERS[8][1] ,
         \REGISTERS[8][0] , \REGISTERS[9][31] , \REGISTERS[9][30] ,
         \REGISTERS[9][29] , \REGISTERS[9][28] , \REGISTERS[9][27] ,
         \REGISTERS[9][26] , \REGISTERS[9][25] , \REGISTERS[9][24] ,
         \REGISTERS[9][23] , \REGISTERS[9][22] , \REGISTERS[9][21] ,
         \REGISTERS[9][20] , \REGISTERS[9][19] , \REGISTERS[9][18] ,
         \REGISTERS[9][17] , \REGISTERS[9][16] , \REGISTERS[9][15] ,
         \REGISTERS[9][14] , \REGISTERS[9][13] , \REGISTERS[9][12] ,
         \REGISTERS[9][11] , \REGISTERS[9][10] , \REGISTERS[9][9] ,
         \REGISTERS[9][8] , \REGISTERS[9][7] , \REGISTERS[9][6] ,
         \REGISTERS[9][5] , \REGISTERS[9][4] , \REGISTERS[9][3] ,
         \REGISTERS[9][2] , \REGISTERS[9][1] , \REGISTERS[9][0] ,
         \REGISTERS[10][31] , \REGISTERS[10][30] , \REGISTERS[10][29] ,
         \REGISTERS[10][28] , \REGISTERS[10][27] , \REGISTERS[10][26] ,
         \REGISTERS[10][25] , \REGISTERS[10][24] , \REGISTERS[10][23] ,
         \REGISTERS[10][22] , \REGISTERS[10][21] , \REGISTERS[10][20] ,
         \REGISTERS[10][19] , \REGISTERS[10][18] , \REGISTERS[10][17] ,
         \REGISTERS[10][16] , \REGISTERS[10][15] , \REGISTERS[10][14] ,
         \REGISTERS[10][13] , \REGISTERS[10][12] , \REGISTERS[10][11] ,
         \REGISTERS[10][10] , \REGISTERS[10][9] , \REGISTERS[10][8] ,
         \REGISTERS[10][7] , \REGISTERS[10][6] , \REGISTERS[10][5] ,
         \REGISTERS[10][4] , \REGISTERS[10][3] , \REGISTERS[10][2] ,
         \REGISTERS[10][1] , \REGISTERS[10][0] , \REGISTERS[11][31] ,
         \REGISTERS[11][30] , \REGISTERS[11][29] , \REGISTERS[11][28] ,
         \REGISTERS[11][27] , \REGISTERS[11][26] , \REGISTERS[11][25] ,
         \REGISTERS[11][24] , \REGISTERS[11][23] , \REGISTERS[11][22] ,
         \REGISTERS[11][21] , \REGISTERS[11][20] , \REGISTERS[11][19] ,
         \REGISTERS[11][18] , \REGISTERS[11][17] , \REGISTERS[11][16] ,
         \REGISTERS[11][15] , \REGISTERS[11][14] , \REGISTERS[11][13] ,
         \REGISTERS[11][12] , \REGISTERS[11][11] , \REGISTERS[11][10] ,
         \REGISTERS[11][9] , \REGISTERS[11][8] , \REGISTERS[11][7] ,
         \REGISTERS[11][6] , \REGISTERS[11][5] , \REGISTERS[11][4] ,
         \REGISTERS[11][3] , \REGISTERS[11][2] , \REGISTERS[11][1] ,
         \REGISTERS[11][0] , \REGISTERS[12][31] , \REGISTERS[12][30] ,
         \REGISTERS[12][29] , \REGISTERS[12][28] , \REGISTERS[12][27] ,
         \REGISTERS[12][26] , \REGISTERS[12][25] , \REGISTERS[12][24] ,
         \REGISTERS[12][23] , \REGISTERS[12][22] , \REGISTERS[12][21] ,
         \REGISTERS[12][20] , \REGISTERS[12][19] , \REGISTERS[12][18] ,
         \REGISTERS[12][17] , \REGISTERS[12][16] , \REGISTERS[12][15] ,
         \REGISTERS[12][14] , \REGISTERS[12][13] , \REGISTERS[12][12] ,
         \REGISTERS[12][11] , \REGISTERS[12][10] , \REGISTERS[12][9] ,
         \REGISTERS[12][8] , \REGISTERS[12][7] , \REGISTERS[12][6] ,
         \REGISTERS[12][5] , \REGISTERS[12][4] , \REGISTERS[12][3] ,
         \REGISTERS[12][2] , \REGISTERS[12][1] , \REGISTERS[12][0] ,
         \REGISTERS[13][31] , \REGISTERS[13][30] , \REGISTERS[13][29] ,
         \REGISTERS[13][28] , \REGISTERS[13][27] , \REGISTERS[13][26] ,
         \REGISTERS[13][25] , \REGISTERS[13][24] , \REGISTERS[13][23] ,
         \REGISTERS[13][22] , \REGISTERS[13][21] , \REGISTERS[13][20] ,
         \REGISTERS[13][19] , \REGISTERS[13][18] , \REGISTERS[13][17] ,
         \REGISTERS[13][16] , \REGISTERS[13][15] , \REGISTERS[13][14] ,
         \REGISTERS[13][13] , \REGISTERS[13][12] , \REGISTERS[13][11] ,
         \REGISTERS[13][10] , \REGISTERS[13][9] , \REGISTERS[13][8] ,
         \REGISTERS[13][7] , \REGISTERS[13][6] , \REGISTERS[13][5] ,
         \REGISTERS[13][4] , \REGISTERS[13][3] , \REGISTERS[13][2] ,
         \REGISTERS[13][1] , \REGISTERS[13][0] , \REGISTERS[14][31] ,
         \REGISTERS[14][30] , \REGISTERS[14][29] , \REGISTERS[14][28] ,
         \REGISTERS[14][27] , \REGISTERS[14][26] , \REGISTERS[14][25] ,
         \REGISTERS[14][24] , \REGISTERS[14][23] , \REGISTERS[14][22] ,
         \REGISTERS[14][21] , \REGISTERS[14][20] , \REGISTERS[14][19] ,
         \REGISTERS[14][18] , \REGISTERS[14][17] , \REGISTERS[14][16] ,
         \REGISTERS[14][15] , \REGISTERS[14][14] , \REGISTERS[14][13] ,
         \REGISTERS[14][12] , \REGISTERS[14][11] , \REGISTERS[14][10] ,
         \REGISTERS[14][9] , \REGISTERS[14][8] , \REGISTERS[14][7] ,
         \REGISTERS[14][6] , \REGISTERS[14][5] , \REGISTERS[14][4] ,
         \REGISTERS[14][3] , \REGISTERS[14][2] , \REGISTERS[14][1] ,
         \REGISTERS[14][0] , \REGISTERS[15][31] , \REGISTERS[15][30] ,
         \REGISTERS[15][29] , \REGISTERS[15][28] , \REGISTERS[15][27] ,
         \REGISTERS[15][26] , \REGISTERS[15][25] , \REGISTERS[15][24] ,
         \REGISTERS[15][23] , \REGISTERS[15][22] , \REGISTERS[15][21] ,
         \REGISTERS[15][20] , \REGISTERS[15][19] , \REGISTERS[15][18] ,
         \REGISTERS[15][17] , \REGISTERS[15][16] , \REGISTERS[15][15] ,
         \REGISTERS[15][14] , \REGISTERS[15][13] , \REGISTERS[15][12] ,
         \REGISTERS[15][11] , \REGISTERS[15][10] , \REGISTERS[15][9] ,
         \REGISTERS[15][8] , \REGISTERS[15][7] , \REGISTERS[15][6] ,
         \REGISTERS[15][5] , \REGISTERS[15][4] , \REGISTERS[15][3] ,
         \REGISTERS[15][2] , \REGISTERS[15][1] , \REGISTERS[15][0] ,
         \REGISTERS[16][31] , \REGISTERS[16][30] , \REGISTERS[16][29] ,
         \REGISTERS[16][28] , \REGISTERS[16][27] , \REGISTERS[16][26] ,
         \REGISTERS[16][25] , \REGISTERS[16][24] , \REGISTERS[16][23] ,
         \REGISTERS[16][22] , \REGISTERS[16][21] , \REGISTERS[16][20] ,
         \REGISTERS[16][19] , \REGISTERS[16][18] , \REGISTERS[16][17] ,
         \REGISTERS[16][16] , \REGISTERS[16][15] , \REGISTERS[16][14] ,
         \REGISTERS[16][13] , \REGISTERS[16][12] , \REGISTERS[16][11] ,
         \REGISTERS[16][10] , \REGISTERS[16][9] , \REGISTERS[16][8] ,
         \REGISTERS[16][7] , \REGISTERS[16][6] , \REGISTERS[16][5] ,
         \REGISTERS[16][4] , \REGISTERS[16][3] , \REGISTERS[16][2] ,
         \REGISTERS[16][1] , \REGISTERS[16][0] , \REGISTERS[17][31] ,
         \REGISTERS[17][30] , \REGISTERS[17][29] , \REGISTERS[17][28] ,
         \REGISTERS[17][27] , \REGISTERS[17][26] , \REGISTERS[17][25] ,
         \REGISTERS[17][24] , \REGISTERS[17][23] , \REGISTERS[17][22] ,
         \REGISTERS[17][21] , \REGISTERS[17][20] , \REGISTERS[17][19] ,
         \REGISTERS[17][18] , \REGISTERS[17][17] , \REGISTERS[17][16] ,
         \REGISTERS[17][15] , \REGISTERS[17][14] , \REGISTERS[17][13] ,
         \REGISTERS[17][12] , \REGISTERS[17][11] , \REGISTERS[17][10] ,
         \REGISTERS[17][9] , \REGISTERS[17][8] , \REGISTERS[17][7] ,
         \REGISTERS[17][6] , \REGISTERS[17][5] , \REGISTERS[17][4] ,
         \REGISTERS[17][3] , \REGISTERS[17][2] , \REGISTERS[17][1] ,
         \REGISTERS[17][0] , \REGISTERS[18][31] , \REGISTERS[18][30] ,
         \REGISTERS[18][29] , \REGISTERS[18][28] , \REGISTERS[18][27] ,
         \REGISTERS[18][26] , \REGISTERS[18][25] , \REGISTERS[18][24] ,
         \REGISTERS[18][23] , \REGISTERS[18][22] , \REGISTERS[18][21] ,
         \REGISTERS[18][20] , \REGISTERS[18][19] , \REGISTERS[18][18] ,
         \REGISTERS[18][17] , \REGISTERS[18][16] , \REGISTERS[18][15] ,
         \REGISTERS[18][14] , \REGISTERS[18][13] , \REGISTERS[18][12] ,
         \REGISTERS[18][11] , \REGISTERS[18][10] , \REGISTERS[18][9] ,
         \REGISTERS[18][8] , \REGISTERS[18][7] , \REGISTERS[18][6] ,
         \REGISTERS[18][5] , \REGISTERS[18][4] , \REGISTERS[18][3] ,
         \REGISTERS[18][2] , \REGISTERS[18][1] , \REGISTERS[18][0] ,
         \REGISTERS[19][31] , \REGISTERS[19][30] , \REGISTERS[19][29] ,
         \REGISTERS[19][28] , \REGISTERS[19][27] , \REGISTERS[19][26] ,
         \REGISTERS[19][25] , \REGISTERS[19][24] , \REGISTERS[19][23] ,
         \REGISTERS[19][22] , \REGISTERS[19][21] , \REGISTERS[19][20] ,
         \REGISTERS[19][19] , \REGISTERS[19][18] , \REGISTERS[19][17] ,
         \REGISTERS[19][16] , \REGISTERS[19][15] , \REGISTERS[19][14] ,
         \REGISTERS[19][13] , \REGISTERS[19][12] , \REGISTERS[19][11] ,
         \REGISTERS[19][10] , \REGISTERS[19][9] , \REGISTERS[19][8] ,
         \REGISTERS[19][7] , \REGISTERS[19][6] , \REGISTERS[19][5] ,
         \REGISTERS[19][4] , \REGISTERS[19][3] , \REGISTERS[19][2] ,
         \REGISTERS[19][1] , \REGISTERS[19][0] , \REGISTERS[20][31] ,
         \REGISTERS[20][30] , \REGISTERS[20][29] , \REGISTERS[20][28] ,
         \REGISTERS[20][27] , \REGISTERS[20][26] , \REGISTERS[20][25] ,
         \REGISTERS[20][24] , \REGISTERS[20][23] , \REGISTERS[20][22] ,
         \REGISTERS[20][21] , \REGISTERS[20][20] , \REGISTERS[20][19] ,
         \REGISTERS[20][18] , \REGISTERS[20][17] , \REGISTERS[20][16] ,
         \REGISTERS[20][15] , \REGISTERS[20][14] , \REGISTERS[20][13] ,
         \REGISTERS[20][12] , \REGISTERS[20][11] , \REGISTERS[20][10] ,
         \REGISTERS[20][9] , \REGISTERS[20][8] , \REGISTERS[20][7] ,
         \REGISTERS[20][6] , \REGISTERS[20][5] , \REGISTERS[20][4] ,
         \REGISTERS[20][3] , \REGISTERS[20][2] , \REGISTERS[20][1] ,
         \REGISTERS[20][0] , \REGISTERS[21][31] , \REGISTERS[21][30] ,
         \REGISTERS[21][29] , \REGISTERS[21][28] , \REGISTERS[21][27] ,
         \REGISTERS[21][26] , \REGISTERS[21][25] , \REGISTERS[21][24] ,
         \REGISTERS[21][23] , \REGISTERS[21][22] , \REGISTERS[21][21] ,
         \REGISTERS[21][20] , \REGISTERS[21][19] , \REGISTERS[21][18] ,
         \REGISTERS[21][17] , \REGISTERS[21][16] , \REGISTERS[21][15] ,
         \REGISTERS[21][14] , \REGISTERS[21][13] , \REGISTERS[21][12] ,
         \REGISTERS[21][11] , \REGISTERS[21][10] , \REGISTERS[21][9] ,
         \REGISTERS[21][8] , \REGISTERS[21][7] , \REGISTERS[21][6] ,
         \REGISTERS[21][5] , \REGISTERS[21][4] , \REGISTERS[21][3] ,
         \REGISTERS[21][2] , \REGISTERS[21][1] , \REGISTERS[21][0] ,
         \REGISTERS[22][31] , \REGISTERS[22][30] , \REGISTERS[22][29] ,
         \REGISTERS[22][28] , \REGISTERS[22][27] , \REGISTERS[22][26] ,
         \REGISTERS[22][25] , \REGISTERS[22][24] , \REGISTERS[22][23] ,
         \REGISTERS[22][22] , \REGISTERS[22][21] , \REGISTERS[22][20] ,
         \REGISTERS[22][19] , \REGISTERS[22][18] , \REGISTERS[22][17] ,
         \REGISTERS[22][16] , \REGISTERS[22][15] , \REGISTERS[22][14] ,
         \REGISTERS[22][13] , \REGISTERS[22][12] , \REGISTERS[22][11] ,
         \REGISTERS[22][10] , \REGISTERS[22][9] , \REGISTERS[22][8] ,
         \REGISTERS[22][7] , \REGISTERS[22][6] , \REGISTERS[22][5] ,
         \REGISTERS[22][4] , \REGISTERS[22][3] , \REGISTERS[22][2] ,
         \REGISTERS[22][1] , \REGISTERS[22][0] , \REGISTERS[23][31] ,
         \REGISTERS[23][30] , \REGISTERS[23][29] , \REGISTERS[23][28] ,
         \REGISTERS[23][27] , \REGISTERS[23][26] , \REGISTERS[23][25] ,
         \REGISTERS[23][24] , \REGISTERS[23][23] , \REGISTERS[23][22] ,
         \REGISTERS[23][21] , \REGISTERS[23][20] , \REGISTERS[23][19] ,
         \REGISTERS[23][18] , \REGISTERS[23][17] , \REGISTERS[23][16] ,
         \REGISTERS[23][15] , \REGISTERS[23][14] , \REGISTERS[23][13] ,
         \REGISTERS[23][12] , \REGISTERS[23][11] , \REGISTERS[23][10] ,
         \REGISTERS[23][9] , \REGISTERS[23][8] , \REGISTERS[23][7] ,
         \REGISTERS[23][6] , \REGISTERS[23][5] , \REGISTERS[23][4] ,
         \REGISTERS[23][3] , \REGISTERS[23][2] , \REGISTERS[23][1] ,
         \REGISTERS[23][0] , \REGISTERS[24][31] , \REGISTERS[24][30] ,
         \REGISTERS[24][29] , \REGISTERS[24][28] , \REGISTERS[24][27] ,
         \REGISTERS[24][26] , \REGISTERS[24][25] , \REGISTERS[24][24] ,
         \REGISTERS[24][23] , \REGISTERS[24][22] , \REGISTERS[24][21] ,
         \REGISTERS[24][20] , \REGISTERS[24][19] , \REGISTERS[24][18] ,
         \REGISTERS[24][17] , \REGISTERS[24][16] , \REGISTERS[24][15] ,
         \REGISTERS[24][14] , \REGISTERS[24][13] , \REGISTERS[24][12] ,
         \REGISTERS[24][11] , \REGISTERS[24][10] , \REGISTERS[24][9] ,
         \REGISTERS[24][8] , \REGISTERS[24][7] , \REGISTERS[24][6] ,
         \REGISTERS[24][5] , \REGISTERS[24][4] , \REGISTERS[24][3] ,
         \REGISTERS[24][2] , \REGISTERS[24][1] , \REGISTERS[24][0] ,
         \REGISTERS[25][31] , \REGISTERS[25][30] , \REGISTERS[25][29] ,
         \REGISTERS[25][28] , \REGISTERS[25][27] , \REGISTERS[25][26] ,
         \REGISTERS[25][25] , \REGISTERS[25][24] , \REGISTERS[25][23] ,
         \REGISTERS[25][22] , \REGISTERS[25][21] , \REGISTERS[25][20] ,
         \REGISTERS[25][19] , \REGISTERS[25][18] , \REGISTERS[25][17] ,
         \REGISTERS[25][16] , \REGISTERS[25][15] , \REGISTERS[25][14] ,
         \REGISTERS[25][13] , \REGISTERS[25][12] , \REGISTERS[25][11] ,
         \REGISTERS[25][10] , \REGISTERS[25][9] , \REGISTERS[25][8] ,
         \REGISTERS[25][7] , \REGISTERS[25][6] , \REGISTERS[25][5] ,
         \REGISTERS[25][4] , \REGISTERS[25][3] , \REGISTERS[25][2] ,
         \REGISTERS[25][1] , \REGISTERS[25][0] , \REGISTERS[26][31] ,
         \REGISTERS[26][30] , \REGISTERS[26][29] , \REGISTERS[26][28] ,
         \REGISTERS[26][27] , \REGISTERS[26][26] , \REGISTERS[26][25] ,
         \REGISTERS[26][24] , \REGISTERS[26][23] , \REGISTERS[26][22] ,
         \REGISTERS[26][21] , \REGISTERS[26][20] , \REGISTERS[26][19] ,
         \REGISTERS[26][18] , \REGISTERS[26][17] , \REGISTERS[26][16] ,
         \REGISTERS[26][15] , \REGISTERS[26][14] , \REGISTERS[26][13] ,
         \REGISTERS[26][12] , \REGISTERS[26][11] , \REGISTERS[26][10] ,
         \REGISTERS[26][9] , \REGISTERS[26][8] , \REGISTERS[26][7] ,
         \REGISTERS[26][6] , \REGISTERS[26][5] , \REGISTERS[26][4] ,
         \REGISTERS[26][3] , \REGISTERS[26][2] , \REGISTERS[26][1] ,
         \REGISTERS[26][0] , \REGISTERS[27][31] , \REGISTERS[27][30] ,
         \REGISTERS[27][29] , \REGISTERS[27][28] , \REGISTERS[27][27] ,
         \REGISTERS[27][26] , \REGISTERS[27][25] , \REGISTERS[27][24] ,
         \REGISTERS[27][23] , \REGISTERS[27][22] , \REGISTERS[27][21] ,
         \REGISTERS[27][20] , \REGISTERS[27][19] , \REGISTERS[27][18] ,
         \REGISTERS[27][17] , \REGISTERS[27][16] , \REGISTERS[27][15] ,
         \REGISTERS[27][14] , \REGISTERS[27][13] , \REGISTERS[27][12] ,
         \REGISTERS[27][11] , \REGISTERS[27][10] , \REGISTERS[27][9] ,
         \REGISTERS[27][8] , \REGISTERS[27][7] , \REGISTERS[27][6] ,
         \REGISTERS[27][5] , \REGISTERS[27][4] , \REGISTERS[27][3] ,
         \REGISTERS[27][2] , \REGISTERS[27][1] , \REGISTERS[27][0] ,
         \REGISTERS[28][31] , \REGISTERS[28][30] , \REGISTERS[28][29] ,
         \REGISTERS[28][28] , \REGISTERS[28][27] , \REGISTERS[28][26] ,
         \REGISTERS[28][25] , \REGISTERS[28][24] , \REGISTERS[28][23] ,
         \REGISTERS[28][22] , \REGISTERS[28][21] , \REGISTERS[28][20] ,
         \REGISTERS[28][19] , \REGISTERS[28][18] , \REGISTERS[28][17] ,
         \REGISTERS[28][16] , \REGISTERS[28][15] , \REGISTERS[28][14] ,
         \REGISTERS[28][13] , \REGISTERS[28][12] , \REGISTERS[28][11] ,
         \REGISTERS[28][10] , \REGISTERS[28][9] , \REGISTERS[28][8] ,
         \REGISTERS[28][7] , \REGISTERS[28][6] , \REGISTERS[28][5] ,
         \REGISTERS[28][4] , \REGISTERS[28][3] , \REGISTERS[28][2] ,
         \REGISTERS[28][1] , \REGISTERS[28][0] , \REGISTERS[29][31] ,
         \REGISTERS[29][30] , \REGISTERS[29][29] , \REGISTERS[29][28] ,
         \REGISTERS[29][27] , \REGISTERS[29][26] , \REGISTERS[29][25] ,
         \REGISTERS[29][24] , \REGISTERS[29][23] , \REGISTERS[29][22] ,
         \REGISTERS[29][21] , \REGISTERS[29][20] , \REGISTERS[29][19] ,
         \REGISTERS[29][18] , \REGISTERS[29][17] , \REGISTERS[29][16] ,
         \REGISTERS[29][15] , \REGISTERS[29][14] , \REGISTERS[29][13] ,
         \REGISTERS[29][12] , \REGISTERS[29][11] , \REGISTERS[29][10] ,
         \REGISTERS[29][9] , \REGISTERS[29][8] , \REGISTERS[29][7] ,
         \REGISTERS[29][6] , \REGISTERS[29][5] , \REGISTERS[29][4] ,
         \REGISTERS[29][3] , \REGISTERS[29][2] , \REGISTERS[29][1] ,
         \REGISTERS[29][0] , \REGISTERS[30][31] , \REGISTERS[30][30] ,
         \REGISTERS[30][29] , \REGISTERS[30][28] , \REGISTERS[30][27] ,
         \REGISTERS[30][26] , \REGISTERS[30][25] , \REGISTERS[30][24] ,
         \REGISTERS[30][23] , \REGISTERS[30][22] , \REGISTERS[30][21] ,
         \REGISTERS[30][20] , \REGISTERS[30][19] , \REGISTERS[30][18] ,
         \REGISTERS[30][17] , \REGISTERS[30][16] , \REGISTERS[30][15] ,
         \REGISTERS[30][14] , \REGISTERS[30][13] , \REGISTERS[30][12] ,
         \REGISTERS[30][11] , \REGISTERS[30][10] , \REGISTERS[30][9] ,
         \REGISTERS[30][8] , \REGISTERS[30][7] , \REGISTERS[30][6] ,
         \REGISTERS[30][5] , \REGISTERS[30][4] , \REGISTERS[30][3] ,
         \REGISTERS[30][2] , \REGISTERS[30][1] , \REGISTERS[30][0] ,
         \REGISTERS[31][31] , \REGISTERS[31][30] , \REGISTERS[31][29] ,
         \REGISTERS[31][28] , \REGISTERS[31][27] , \REGISTERS[31][26] ,
         \REGISTERS[31][25] , \REGISTERS[31][24] , \REGISTERS[31][23] ,
         \REGISTERS[31][22] , \REGISTERS[31][21] , \REGISTERS[31][20] ,
         \REGISTERS[31][19] , \REGISTERS[31][18] , \REGISTERS[31][17] ,
         \REGISTERS[31][16] , \REGISTERS[31][15] , \REGISTERS[31][14] ,
         \REGISTERS[31][13] , \REGISTERS[31][12] , \REGISTERS[31][11] ,
         \REGISTERS[31][10] , \REGISTERS[31][9] , \REGISTERS[31][8] ,
         \REGISTERS[31][7] , \REGISTERS[31][6] , \REGISTERS[31][5] ,
         \REGISTERS[31][4] , \REGISTERS[31][3] , \REGISTERS[31][2] ,
         \REGISTERS[31][1] , \REGISTERS[31][0] , N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n558, n1182, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157;

  DLH_X1 \REGISTERS_reg[1][31]  ( .G(n195), .D(n283), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(n195), .D(n286), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(n195), .D(n289), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(n195), .D(n292), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(n195), .D(n295), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(n195), .D(n298), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(n195), .D(n301), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(n195), .D(n304), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(n195), .D(n307), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(n195), .D(n310), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(n194), .D(n313), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n194), .D(n316), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n194), .D(n319), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(n194), .D(n322), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(n194), .D(n325), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(n194), .D(n328), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(n194), .D(n331), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(n194), .D(n334), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(n194), .D(n337), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(n194), .D(n340), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n194), .D(n343), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(n193), .D(n346), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(n193), .D(n349), .Q(\REGISTERS[1][9] ) );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(n193), .D(n352), .Q(\REGISTERS[1][8] ) );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n193), .D(n355), .Q(\REGISTERS[1][7] ) );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(n193), .D(n358), .Q(\REGISTERS[1][6] ) );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n193), .D(n361), .Q(\REGISTERS[1][5] ) );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(n193), .D(n364), .Q(\REGISTERS[1][4] ) );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(n193), .D(n367), .Q(\REGISTERS[1][3] ) );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(n193), .D(n370), .Q(\REGISTERS[1][2] ) );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(n193), .D(n373), .Q(\REGISTERS[1][1] ) );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n193), .D(n376), .Q(\REGISTERS[1][0] ) );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(n198), .D(n283), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(n198), .D(n286), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(n198), .D(n289), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(n198), .D(n292), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(n198), .D(n295), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(n198), .D(n298), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(n198), .D(n301), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(n198), .D(n304), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n198), .D(n307), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n198), .D(n310), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(n197), .D(n313), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(n197), .D(n316), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n197), .D(n319), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(n197), .D(n322), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n197), .D(n325), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(n197), .D(n328), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(n197), .D(n331), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(n197), .D(n334), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(n197), .D(n337), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(n197), .D(n340), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(n197), .D(n343), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n196), .D(n346), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(n196), .D(n349), .Q(\REGISTERS[2][9] ) );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(n196), .D(n352), .Q(\REGISTERS[2][8] ) );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n196), .D(n355), .Q(\REGISTERS[2][7] ) );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(n196), .D(n358), .Q(\REGISTERS[2][6] ) );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(n196), .D(n361), .Q(\REGISTERS[2][5] ) );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(n196), .D(n364), .Q(\REGISTERS[2][4] ) );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(n196), .D(n367), .Q(\REGISTERS[2][3] ) );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(n196), .D(n370), .Q(\REGISTERS[2][2] ) );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(n196), .D(n373), .Q(\REGISTERS[2][1] ) );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(n196), .D(n376), .Q(\REGISTERS[2][0] ) );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(n201), .D(n283), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(n201), .D(n286), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(n201), .D(n289), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(n201), .D(n292), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(n201), .D(n295), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(n201), .D(n298), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(n201), .D(n301), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(n201), .D(n304), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n201), .D(n307), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n201), .D(n310), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(n200), .D(n313), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(n200), .D(n316), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n200), .D(n319), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(n200), .D(n322), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n200), .D(n325), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(n200), .D(n328), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(n200), .D(n331), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(n200), .D(n334), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(n200), .D(n337), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(n200), .D(n340), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(n200), .D(n343), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n199), .D(n346), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(n199), .D(n349), .Q(\REGISTERS[3][9] ) );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(n199), .D(n352), .Q(\REGISTERS[3][8] ) );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n199), .D(n355), .Q(\REGISTERS[3][7] ) );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(n199), .D(n358), .Q(\REGISTERS[3][6] ) );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(n199), .D(n361), .Q(\REGISTERS[3][5] ) );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(n199), .D(n364), .Q(\REGISTERS[3][4] ) );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(n199), .D(n367), .Q(\REGISTERS[3][3] ) );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(n199), .D(n370), .Q(\REGISTERS[3][2] ) );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(n199), .D(n373), .Q(\REGISTERS[3][1] ) );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(n199), .D(n376), .Q(\REGISTERS[3][0] ) );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(n204), .D(n283), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(n204), .D(n286), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(n204), .D(n289), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(n204), .D(n292), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(n204), .D(n295), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(n204), .D(n298), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(n204), .D(n301), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(n204), .D(n304), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n204), .D(n307), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n204), .D(n310), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(n203), .D(n313), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(n203), .D(n316), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n203), .D(n319), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(n203), .D(n322), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n203), .D(n325), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(n203), .D(n328), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(n203), .D(n331), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(n203), .D(n334), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(n203), .D(n337), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(n203), .D(n340), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(n203), .D(n343), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n202), .D(n346), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(n202), .D(n349), .Q(\REGISTERS[4][9] ) );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(n202), .D(n352), .Q(\REGISTERS[4][8] ) );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(n202), .D(n355), .Q(\REGISTERS[4][7] ) );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(n202), .D(n358), .Q(\REGISTERS[4][6] ) );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(n202), .D(n361), .Q(\REGISTERS[4][5] ) );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(n202), .D(n364), .Q(\REGISTERS[4][4] ) );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(n202), .D(n367), .Q(\REGISTERS[4][3] ) );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(n202), .D(n370), .Q(\REGISTERS[4][2] ) );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(n202), .D(n373), .Q(\REGISTERS[4][1] ) );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n202), .D(n376), .Q(\REGISTERS[4][0] ) );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(n207), .D(n283), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(n207), .D(n286), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(n207), .D(n289), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(n207), .D(n292), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(n207), .D(n295), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(n207), .D(n298), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(n207), .D(n301), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(n207), .D(n304), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n207), .D(n307), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n207), .D(n310), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(n206), .D(n313), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(n206), .D(n316), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n206), .D(n319), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(n206), .D(n322), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n206), .D(n325), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(n206), .D(n328), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(n206), .D(n331), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(n206), .D(n334), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(n206), .D(n337), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(n206), .D(n340), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(n206), .D(n343), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n205), .D(n346), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(n205), .D(n349), .Q(\REGISTERS[5][9] ) );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(n205), .D(n352), .Q(\REGISTERS[5][8] ) );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n205), .D(n355), .Q(\REGISTERS[5][7] ) );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(n205), .D(n358), .Q(\REGISTERS[5][6] ) );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(n205), .D(n361), .Q(\REGISTERS[5][5] ) );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(n205), .D(n364), .Q(\REGISTERS[5][4] ) );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(n205), .D(n367), .Q(\REGISTERS[5][3] ) );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(n205), .D(n370), .Q(\REGISTERS[5][2] ) );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(n205), .D(n373), .Q(\REGISTERS[5][1] ) );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(n205), .D(n376), .Q(\REGISTERS[5][0] ) );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(n210), .D(n283), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(n210), .D(n286), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(n210), .D(n289), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(n210), .D(n292), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(n210), .D(n295), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(n210), .D(n298), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(n210), .D(n301), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(n210), .D(n304), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n210), .D(n307), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n210), .D(n310), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(n209), .D(n313), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(n209), .D(n316), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n209), .D(n319), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(n209), .D(n322), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n209), .D(n325), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(n209), .D(n328), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(n209), .D(n331), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(n209), .D(n334), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(n209), .D(n337), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(n209), .D(n340), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(n209), .D(n343), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n208), .D(n346), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(n208), .D(n349), .Q(\REGISTERS[6][9] ) );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(n208), .D(n352), .Q(\REGISTERS[6][8] ) );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(n208), .D(n355), .Q(\REGISTERS[6][7] ) );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(n208), .D(n358), .Q(\REGISTERS[6][6] ) );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(n208), .D(n361), .Q(\REGISTERS[6][5] ) );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(n208), .D(n364), .Q(\REGISTERS[6][4] ) );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(n208), .D(n367), .Q(\REGISTERS[6][3] ) );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(n208), .D(n370), .Q(\REGISTERS[6][2] ) );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(n208), .D(n373), .Q(\REGISTERS[6][1] ) );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n208), .D(n376), .Q(\REGISTERS[6][0] ) );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(n213), .D(n283), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(n213), .D(n286), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(n213), .D(n289), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(n213), .D(n292), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(n213), .D(n295), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(n213), .D(n298), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(n213), .D(n301), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(n213), .D(n304), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n213), .D(n307), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n213), .D(n310), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(n212), .D(n313), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(n212), .D(n316), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n212), .D(n319), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(n212), .D(n322), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n212), .D(n325), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(n212), .D(n328), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(n212), .D(n331), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(n212), .D(n334), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(n212), .D(n337), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(n212), .D(n340), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(n212), .D(n343), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n211), .D(n346), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(n211), .D(n349), .Q(\REGISTERS[7][9] ) );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(n211), .D(n352), .Q(\REGISTERS[7][8] ) );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n211), .D(n355), .Q(\REGISTERS[7][7] ) );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(n211), .D(n358), .Q(\REGISTERS[7][6] ) );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(n211), .D(n361), .Q(\REGISTERS[7][5] ) );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(n211), .D(n364), .Q(\REGISTERS[7][4] ) );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(n211), .D(n367), .Q(\REGISTERS[7][3] ) );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(n211), .D(n370), .Q(\REGISTERS[7][2] ) );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(n211), .D(n373), .Q(\REGISTERS[7][1] ) );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(n211), .D(n376), .Q(\REGISTERS[7][0] ) );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(n216), .D(n283), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(n216), .D(n286), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(n216), .D(n289), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(n216), .D(n292), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(n216), .D(n295), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(n216), .D(n298), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(n216), .D(n301), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(n216), .D(n304), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n216), .D(n307), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n216), .D(n310), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(n215), .D(n313), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(n215), .D(n316), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n215), .D(n319), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(n215), .D(n322), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n215), .D(n325), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(n215), .D(n328), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(n215), .D(n331), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(n215), .D(n334), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(n215), .D(n337), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(n215), .D(n340), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(n215), .D(n343), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n214), .D(n346), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(n214), .D(n349), .Q(\REGISTERS[8][9] ) );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(n214), .D(n352), .Q(\REGISTERS[8][8] ) );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n214), .D(n355), .Q(\REGISTERS[8][7] ) );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(n214), .D(n358), .Q(\REGISTERS[8][6] ) );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(n214), .D(n361), .Q(\REGISTERS[8][5] ) );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(n214), .D(n364), .Q(\REGISTERS[8][4] ) );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(n214), .D(n367), .Q(\REGISTERS[8][3] ) );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(n214), .D(n370), .Q(\REGISTERS[8][2] ) );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(n214), .D(n373), .Q(\REGISTERS[8][1] ) );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(n214), .D(n376), .Q(\REGISTERS[8][0] ) );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(n219), .D(n283), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(n219), .D(n286), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(n219), .D(n289), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(n219), .D(n292), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(n219), .D(n295), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(n219), .D(n298), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(n219), .D(n301), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(n219), .D(n304), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n219), .D(n307), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n219), .D(n310), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(n218), .D(n313), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(n218), .D(n316), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n218), .D(n319), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(n218), .D(n322), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n218), .D(n325), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(n218), .D(n328), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(n218), .D(n331), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(n218), .D(n334), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(n218), .D(n337), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(n218), .D(n340), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(n218), .D(n343), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n217), .D(n346), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(n217), .D(n349), .Q(\REGISTERS[9][9] ) );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(n217), .D(n352), .Q(\REGISTERS[9][8] ) );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n217), .D(n355), .Q(\REGISTERS[9][7] ) );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(n217), .D(n358), .Q(\REGISTERS[9][6] ) );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(n217), .D(n361), .Q(\REGISTERS[9][5] ) );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(n217), .D(n364), .Q(\REGISTERS[9][4] ) );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(n217), .D(n367), .Q(\REGISTERS[9][3] ) );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(n217), .D(n370), .Q(\REGISTERS[9][2] ) );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(n217), .D(n373), .Q(\REGISTERS[9][1] ) );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(n217), .D(n376), .Q(\REGISTERS[9][0] ) );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(n222), .D(n283), .Q(\REGISTERS[10][31] )
         );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(n222), .D(n286), .Q(\REGISTERS[10][30] )
         );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(n222), .D(n289), .Q(\REGISTERS[10][29] )
         );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(n222), .D(n292), .Q(\REGISTERS[10][28] )
         );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(n222), .D(n295), .Q(\REGISTERS[10][27] )
         );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(n222), .D(n298), .Q(\REGISTERS[10][26] )
         );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(n222), .D(n301), .Q(\REGISTERS[10][25] )
         );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(n222), .D(n304), .Q(\REGISTERS[10][24] )
         );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n222), .D(n307), .Q(\REGISTERS[10][23] )
         );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(n222), .D(n310), .Q(\REGISTERS[10][22] )
         );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(n221), .D(n313), .Q(\REGISTERS[10][21] )
         );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(n221), .D(n316), .Q(\REGISTERS[10][20] )
         );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n221), .D(n319), .Q(\REGISTERS[10][19] )
         );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(n221), .D(n322), .Q(\REGISTERS[10][18] )
         );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(n221), .D(n325), .Q(\REGISTERS[10][17] )
         );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n221), .D(n328), .Q(\REGISTERS[10][16] )
         );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(n221), .D(n331), .Q(\REGISTERS[10][15] )
         );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(n221), .D(n334), .Q(\REGISTERS[10][14] )
         );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n221), .D(n337), .Q(\REGISTERS[10][13] )
         );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(n221), .D(n340), .Q(\REGISTERS[10][12] )
         );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n221), .D(n343), .Q(\REGISTERS[10][11] )
         );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n220), .D(n346), .Q(\REGISTERS[10][10] )
         );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(n220), .D(n349), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(n220), .D(n352), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(n220), .D(n355), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(n220), .D(n358), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(n220), .D(n361), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(n220), .D(n364), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(n220), .D(n367), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(n220), .D(n370), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(n220), .D(n373), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(n220), .D(n376), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(n225), .D(n283), .Q(\REGISTERS[11][31] )
         );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(n225), .D(n286), .Q(\REGISTERS[11][30] )
         );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(n225), .D(n289), .Q(\REGISTERS[11][29] )
         );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(n225), .D(n292), .Q(\REGISTERS[11][28] )
         );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(n225), .D(n295), .Q(\REGISTERS[11][27] )
         );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(n225), .D(n298), .Q(\REGISTERS[11][26] )
         );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(n225), .D(n301), .Q(\REGISTERS[11][25] )
         );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(n225), .D(n304), .Q(\REGISTERS[11][24] )
         );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n225), .D(n307), .Q(\REGISTERS[11][23] )
         );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n225), .D(n310), .Q(\REGISTERS[11][22] )
         );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(n224), .D(n313), .Q(\REGISTERS[11][21] )
         );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(n224), .D(n316), .Q(\REGISTERS[11][20] )
         );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n224), .D(n319), .Q(\REGISTERS[11][19] )
         );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(n224), .D(n322), .Q(\REGISTERS[11][18] )
         );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n224), .D(n325), .Q(\REGISTERS[11][17] )
         );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(n224), .D(n328), .Q(\REGISTERS[11][16] )
         );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(n224), .D(n331), .Q(\REGISTERS[11][15] )
         );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(n224), .D(n334), .Q(\REGISTERS[11][14] )
         );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(n224), .D(n337), .Q(\REGISTERS[11][13] )
         );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(n224), .D(n340), .Q(\REGISTERS[11][12] )
         );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(n224), .D(n343), .Q(\REGISTERS[11][11] )
         );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n223), .D(n346), .Q(\REGISTERS[11][10] )
         );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(n223), .D(n349), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(n223), .D(n352), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n223), .D(n355), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(n223), .D(n358), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(n223), .D(n361), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(n223), .D(n364), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(n223), .D(n367), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(n223), .D(n370), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(n223), .D(n373), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(n223), .D(n376), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(n228), .D(n284), .Q(\REGISTERS[12][31] )
         );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(n228), .D(n287), .Q(\REGISTERS[12][30] )
         );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(n228), .D(n290), .Q(\REGISTERS[12][29] )
         );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(n228), .D(n293), .Q(\REGISTERS[12][28] )
         );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(n228), .D(n296), .Q(\REGISTERS[12][27] )
         );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(n228), .D(n299), .Q(\REGISTERS[12][26] )
         );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(n228), .D(n302), .Q(\REGISTERS[12][25] )
         );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(n228), .D(n305), .Q(\REGISTERS[12][24] )
         );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n228), .D(n308), .Q(\REGISTERS[12][23] )
         );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n228), .D(n311), .Q(\REGISTERS[12][22] )
         );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(n227), .D(n314), .Q(\REGISTERS[12][21] )
         );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(n227), .D(n317), .Q(\REGISTERS[12][20] )
         );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n227), .D(n320), .Q(\REGISTERS[12][19] )
         );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(n227), .D(n323), .Q(\REGISTERS[12][18] )
         );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n227), .D(n326), .Q(\REGISTERS[12][17] )
         );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(n227), .D(n329), .Q(\REGISTERS[12][16] )
         );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(n227), .D(n332), .Q(\REGISTERS[12][15] )
         );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(n227), .D(n335), .Q(\REGISTERS[12][14] )
         );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(n227), .D(n338), .Q(\REGISTERS[12][13] )
         );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(n227), .D(n341), .Q(\REGISTERS[12][12] )
         );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n227), .D(n344), .Q(\REGISTERS[12][11] )
         );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n226), .D(n347), .Q(\REGISTERS[12][10] )
         );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(n226), .D(n350), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(n226), .D(n353), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(n226), .D(n356), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(n226), .D(n359), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(n226), .D(n362), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(n226), .D(n365), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(n226), .D(n368), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(n226), .D(n371), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(n226), .D(n374), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(n226), .D(n377), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(n231), .D(n284), .Q(\REGISTERS[13][31] )
         );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(n231), .D(n287), .Q(\REGISTERS[13][30] )
         );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(n231), .D(n290), .Q(\REGISTERS[13][29] )
         );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(n231), .D(n293), .Q(\REGISTERS[13][28] )
         );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(n231), .D(n296), .Q(\REGISTERS[13][27] )
         );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(n231), .D(n299), .Q(\REGISTERS[13][26] )
         );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(n231), .D(n302), .Q(\REGISTERS[13][25] )
         );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(n231), .D(n305), .Q(\REGISTERS[13][24] )
         );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n231), .D(n308), .Q(\REGISTERS[13][23] )
         );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n231), .D(n311), .Q(\REGISTERS[13][22] )
         );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(n230), .D(n314), .Q(\REGISTERS[13][21] )
         );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(n230), .D(n317), .Q(\REGISTERS[13][20] )
         );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n230), .D(n320), .Q(\REGISTERS[13][19] )
         );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(n230), .D(n323), .Q(\REGISTERS[13][18] )
         );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n230), .D(n326), .Q(\REGISTERS[13][17] )
         );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(n230), .D(n329), .Q(\REGISTERS[13][16] )
         );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(n230), .D(n332), .Q(\REGISTERS[13][15] )
         );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(n230), .D(n335), .Q(\REGISTERS[13][14] )
         );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(n230), .D(n338), .Q(\REGISTERS[13][13] )
         );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(n230), .D(n341), .Q(\REGISTERS[13][12] )
         );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(n230), .D(n344), .Q(\REGISTERS[13][11] )
         );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n229), .D(n347), .Q(\REGISTERS[13][10] )
         );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(n229), .D(n350), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(n229), .D(n353), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n229), .D(n356), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(n229), .D(n359), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(n229), .D(n362), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(n229), .D(n365), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(n229), .D(n368), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(n229), .D(n371), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(n229), .D(n374), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(n229), .D(n377), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(n234), .D(n284), .Q(\REGISTERS[14][31] )
         );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(n234), .D(n287), .Q(\REGISTERS[14][30] )
         );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(n234), .D(n290), .Q(\REGISTERS[14][29] )
         );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(n234), .D(n293), .Q(\REGISTERS[14][28] )
         );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(n234), .D(n296), .Q(\REGISTERS[14][27] )
         );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(n234), .D(n299), .Q(\REGISTERS[14][26] )
         );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(n234), .D(n302), .Q(\REGISTERS[14][25] )
         );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(n234), .D(n305), .Q(\REGISTERS[14][24] )
         );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n234), .D(n308), .Q(\REGISTERS[14][23] )
         );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n234), .D(n311), .Q(\REGISTERS[14][22] )
         );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(n233), .D(n314), .Q(\REGISTERS[14][21] )
         );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(n233), .D(n317), .Q(\REGISTERS[14][20] )
         );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n233), .D(n320), .Q(\REGISTERS[14][19] )
         );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(n233), .D(n323), .Q(\REGISTERS[14][18] )
         );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n233), .D(n326), .Q(\REGISTERS[14][17] )
         );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(n233), .D(n329), .Q(\REGISTERS[14][16] )
         );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(n233), .D(n332), .Q(\REGISTERS[14][15] )
         );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(n233), .D(n335), .Q(\REGISTERS[14][14] )
         );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(n233), .D(n338), .Q(\REGISTERS[14][13] )
         );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(n233), .D(n341), .Q(\REGISTERS[14][12] )
         );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(n233), .D(n344), .Q(\REGISTERS[14][11] )
         );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n232), .D(n347), .Q(\REGISTERS[14][10] )
         );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(n232), .D(n350), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(n232), .D(n353), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n232), .D(n356), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(n232), .D(n359), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(n232), .D(n362), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(n232), .D(n365), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(n232), .D(n368), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(n232), .D(n371), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(n232), .D(n374), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(n232), .D(n377), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(n237), .D(n284), .Q(\REGISTERS[15][31] )
         );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(n237), .D(n287), .Q(\REGISTERS[15][30] )
         );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(n237), .D(n290), .Q(\REGISTERS[15][29] )
         );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(n237), .D(n293), .Q(\REGISTERS[15][28] )
         );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(n237), .D(n296), .Q(\REGISTERS[15][27] )
         );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(n237), .D(n299), .Q(\REGISTERS[15][26] )
         );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(n237), .D(n302), .Q(\REGISTERS[15][25] )
         );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(n237), .D(n305), .Q(\REGISTERS[15][24] )
         );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n237), .D(n308), .Q(\REGISTERS[15][23] )
         );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n237), .D(n311), .Q(\REGISTERS[15][22] )
         );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(n236), .D(n314), .Q(\REGISTERS[15][21] )
         );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(n236), .D(n317), .Q(\REGISTERS[15][20] )
         );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n236), .D(n320), .Q(\REGISTERS[15][19] )
         );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(n236), .D(n323), .Q(\REGISTERS[15][18] )
         );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n236), .D(n326), .Q(\REGISTERS[15][17] )
         );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(n236), .D(n329), .Q(\REGISTERS[15][16] )
         );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(n236), .D(n332), .Q(\REGISTERS[15][15] )
         );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(n236), .D(n335), .Q(\REGISTERS[15][14] )
         );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(n236), .D(n338), .Q(\REGISTERS[15][13] )
         );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(n236), .D(n341), .Q(\REGISTERS[15][12] )
         );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(n236), .D(n344), .Q(\REGISTERS[15][11] )
         );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n235), .D(n347), .Q(\REGISTERS[15][10] )
         );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(n235), .D(n350), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(n235), .D(n353), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n235), .D(n356), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(n235), .D(n359), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(n235), .D(n362), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(n235), .D(n365), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(n235), .D(n368), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(n235), .D(n371), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(n235), .D(n374), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(n235), .D(n377), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(n240), .D(n284), .Q(\REGISTERS[16][31] )
         );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(n240), .D(n287), .Q(\REGISTERS[16][30] )
         );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(n240), .D(n290), .Q(\REGISTERS[16][29] )
         );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(n240), .D(n293), .Q(\REGISTERS[16][28] )
         );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(n240), .D(n296), .Q(\REGISTERS[16][27] )
         );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(n240), .D(n299), .Q(\REGISTERS[16][26] )
         );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(n240), .D(n302), .Q(\REGISTERS[16][25] )
         );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(n240), .D(n305), .Q(\REGISTERS[16][24] )
         );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n240), .D(n308), .Q(\REGISTERS[16][23] )
         );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n240), .D(n311), .Q(\REGISTERS[16][22] )
         );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(n239), .D(n314), .Q(\REGISTERS[16][21] )
         );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(n239), .D(n317), .Q(\REGISTERS[16][20] )
         );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n239), .D(n320), .Q(\REGISTERS[16][19] )
         );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(n239), .D(n323), .Q(\REGISTERS[16][18] )
         );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n239), .D(n326), .Q(\REGISTERS[16][17] )
         );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(n239), .D(n329), .Q(\REGISTERS[16][16] )
         );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(n239), .D(n332), .Q(\REGISTERS[16][15] )
         );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(n239), .D(n335), .Q(\REGISTERS[16][14] )
         );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(n239), .D(n338), .Q(\REGISTERS[16][13] )
         );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(n239), .D(n341), .Q(\REGISTERS[16][12] )
         );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(n239), .D(n344), .Q(\REGISTERS[16][11] )
         );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n238), .D(n347), .Q(\REGISTERS[16][10] )
         );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(n238), .D(n350), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(n238), .D(n353), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n238), .D(n356), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(n238), .D(n359), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(n238), .D(n362), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(n238), .D(n365), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(n238), .D(n368), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(n238), .D(n371), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(n238), .D(n374), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(n238), .D(n377), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(n243), .D(n284), .Q(\REGISTERS[17][31] )
         );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(n243), .D(n287), .Q(\REGISTERS[17][30] )
         );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(n243), .D(n290), .Q(\REGISTERS[17][29] )
         );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(n243), .D(n293), .Q(\REGISTERS[17][28] )
         );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(n243), .D(n296), .Q(\REGISTERS[17][27] )
         );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(n243), .D(n299), .Q(\REGISTERS[17][26] )
         );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(n243), .D(n302), .Q(\REGISTERS[17][25] )
         );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(n243), .D(n305), .Q(\REGISTERS[17][24] )
         );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n243), .D(n308), .Q(\REGISTERS[17][23] )
         );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n243), .D(n311), .Q(\REGISTERS[17][22] )
         );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(n242), .D(n314), .Q(\REGISTERS[17][21] )
         );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(n242), .D(n317), .Q(\REGISTERS[17][20] )
         );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n242), .D(n320), .Q(\REGISTERS[17][19] )
         );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(n242), .D(n323), .Q(\REGISTERS[17][18] )
         );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n242), .D(n326), .Q(\REGISTERS[17][17] )
         );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(n242), .D(n329), .Q(\REGISTERS[17][16] )
         );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(n242), .D(n332), .Q(\REGISTERS[17][15] )
         );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(n242), .D(n335), .Q(\REGISTERS[17][14] )
         );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(n242), .D(n338), .Q(\REGISTERS[17][13] )
         );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(n242), .D(n341), .Q(\REGISTERS[17][12] )
         );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(n242), .D(n344), .Q(\REGISTERS[17][11] )
         );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n241), .D(n347), .Q(\REGISTERS[17][10] )
         );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(n241), .D(n350), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(n241), .D(n353), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n241), .D(n356), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(n241), .D(n359), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(n241), .D(n362), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(n241), .D(n365), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(n241), .D(n368), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(n241), .D(n371), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(n241), .D(n374), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(n241), .D(n377), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(n246), .D(n284), .Q(\REGISTERS[18][31] )
         );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(n246), .D(n287), .Q(\REGISTERS[18][30] )
         );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(n246), .D(n290), .Q(\REGISTERS[18][29] )
         );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(n246), .D(n293), .Q(\REGISTERS[18][28] )
         );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(n246), .D(n296), .Q(\REGISTERS[18][27] )
         );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(n246), .D(n299), .Q(\REGISTERS[18][26] )
         );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(n246), .D(n302), .Q(\REGISTERS[18][25] )
         );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(n246), .D(n305), .Q(\REGISTERS[18][24] )
         );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n246), .D(n308), .Q(\REGISTERS[18][23] )
         );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n246), .D(n311), .Q(\REGISTERS[18][22] )
         );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(n245), .D(n314), .Q(\REGISTERS[18][21] )
         );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(n245), .D(n317), .Q(\REGISTERS[18][20] )
         );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n245), .D(n320), .Q(\REGISTERS[18][19] )
         );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(n245), .D(n323), .Q(\REGISTERS[18][18] )
         );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n245), .D(n326), .Q(\REGISTERS[18][17] )
         );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(n245), .D(n329), .Q(\REGISTERS[18][16] )
         );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(n245), .D(n332), .Q(\REGISTERS[18][15] )
         );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(n245), .D(n335), .Q(\REGISTERS[18][14] )
         );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(n245), .D(n338), .Q(\REGISTERS[18][13] )
         );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(n245), .D(n341), .Q(\REGISTERS[18][12] )
         );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(n245), .D(n344), .Q(\REGISTERS[18][11] )
         );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n244), .D(n347), .Q(\REGISTERS[18][10] )
         );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(n244), .D(n350), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(n244), .D(n353), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n244), .D(n356), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(n244), .D(n359), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(n244), .D(n362), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(n244), .D(n365), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(n244), .D(n368), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(n244), .D(n371), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(n244), .D(n374), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(n244), .D(n377), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(n249), .D(n284), .Q(\REGISTERS[19][31] )
         );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(n249), .D(n287), .Q(\REGISTERS[19][30] )
         );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(n249), .D(n290), .Q(\REGISTERS[19][29] )
         );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(n249), .D(n293), .Q(\REGISTERS[19][28] )
         );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(n249), .D(n296), .Q(\REGISTERS[19][27] )
         );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(n249), .D(n299), .Q(\REGISTERS[19][26] )
         );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(n249), .D(n302), .Q(\REGISTERS[19][25] )
         );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(n249), .D(n305), .Q(\REGISTERS[19][24] )
         );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n249), .D(n308), .Q(\REGISTERS[19][23] )
         );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n249), .D(n311), .Q(\REGISTERS[19][22] )
         );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(n248), .D(n314), .Q(\REGISTERS[19][21] )
         );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(n248), .D(n317), .Q(\REGISTERS[19][20] )
         );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n248), .D(n320), .Q(\REGISTERS[19][19] )
         );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(n248), .D(n323), .Q(\REGISTERS[19][18] )
         );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n248), .D(n326), .Q(\REGISTERS[19][17] )
         );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(n248), .D(n329), .Q(\REGISTERS[19][16] )
         );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(n248), .D(n332), .Q(\REGISTERS[19][15] )
         );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(n248), .D(n335), .Q(\REGISTERS[19][14] )
         );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(n248), .D(n338), .Q(\REGISTERS[19][13] )
         );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(n248), .D(n341), .Q(\REGISTERS[19][12] )
         );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(n248), .D(n344), .Q(\REGISTERS[19][11] )
         );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n247), .D(n347), .Q(\REGISTERS[19][10] )
         );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(n247), .D(n350), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(n247), .D(n353), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n247), .D(n356), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(n247), .D(n359), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(n247), .D(n362), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(n247), .D(n365), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(n247), .D(n368), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(n247), .D(n371), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(n247), .D(n374), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(n247), .D(n377), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(n252), .D(n284), .Q(\REGISTERS[20][31] )
         );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(n252), .D(n287), .Q(\REGISTERS[20][30] )
         );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(n252), .D(n290), .Q(\REGISTERS[20][29] )
         );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(n252), .D(n293), .Q(\REGISTERS[20][28] )
         );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(n252), .D(n296), .Q(\REGISTERS[20][27] )
         );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(n252), .D(n299), .Q(\REGISTERS[20][26] )
         );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(n252), .D(n302), .Q(\REGISTERS[20][25] )
         );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(n252), .D(n305), .Q(\REGISTERS[20][24] )
         );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n252), .D(n308), .Q(\REGISTERS[20][23] )
         );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n252), .D(n311), .Q(\REGISTERS[20][22] )
         );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(n251), .D(n314), .Q(\REGISTERS[20][21] )
         );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(n251), .D(n317), .Q(\REGISTERS[20][20] )
         );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n251), .D(n320), .Q(\REGISTERS[20][19] )
         );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(n251), .D(n323), .Q(\REGISTERS[20][18] )
         );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n251), .D(n326), .Q(\REGISTERS[20][17] )
         );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(n251), .D(n329), .Q(\REGISTERS[20][16] )
         );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(n251), .D(n332), .Q(\REGISTERS[20][15] )
         );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(n251), .D(n335), .Q(\REGISTERS[20][14] )
         );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(n251), .D(n338), .Q(\REGISTERS[20][13] )
         );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(n251), .D(n341), .Q(\REGISTERS[20][12] )
         );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(n251), .D(n344), .Q(\REGISTERS[20][11] )
         );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n250), .D(n347), .Q(\REGISTERS[20][10] )
         );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(n250), .D(n350), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(n250), .D(n353), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n250), .D(n356), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(n250), .D(n359), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(n250), .D(n362), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(n250), .D(n365), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(n250), .D(n368), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(n250), .D(n371), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(n250), .D(n374), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(n250), .D(n377), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(n255), .D(n284), .Q(\REGISTERS[21][31] )
         );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(n255), .D(n287), .Q(\REGISTERS[21][30] )
         );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(n255), .D(n290), .Q(\REGISTERS[21][29] )
         );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(n255), .D(n293), .Q(\REGISTERS[21][28] )
         );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(n255), .D(n296), .Q(\REGISTERS[21][27] )
         );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(n255), .D(n299), .Q(\REGISTERS[21][26] )
         );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(n255), .D(n302), .Q(\REGISTERS[21][25] )
         );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(n255), .D(n305), .Q(\REGISTERS[21][24] )
         );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n255), .D(n308), .Q(\REGISTERS[21][23] )
         );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n255), .D(n311), .Q(\REGISTERS[21][22] )
         );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(n254), .D(n314), .Q(\REGISTERS[21][21] )
         );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(n254), .D(n317), .Q(\REGISTERS[21][20] )
         );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n254), .D(n320), .Q(\REGISTERS[21][19] )
         );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(n254), .D(n323), .Q(\REGISTERS[21][18] )
         );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n254), .D(n326), .Q(\REGISTERS[21][17] )
         );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(n254), .D(n329), .Q(\REGISTERS[21][16] )
         );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(n254), .D(n332), .Q(\REGISTERS[21][15] )
         );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(n254), .D(n335), .Q(\REGISTERS[21][14] )
         );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(n254), .D(n338), .Q(\REGISTERS[21][13] )
         );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(n254), .D(n341), .Q(\REGISTERS[21][12] )
         );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(n254), .D(n344), .Q(\REGISTERS[21][11] )
         );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n253), .D(n347), .Q(\REGISTERS[21][10] )
         );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(n253), .D(n350), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(n253), .D(n353), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n253), .D(n356), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(n253), .D(n359), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(n253), .D(n362), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(n253), .D(n365), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(n253), .D(n368), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(n253), .D(n371), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(n253), .D(n374), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(n253), .D(n377), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(n258), .D(n284), .Q(\REGISTERS[22][31] )
         );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(n258), .D(n287), .Q(\REGISTERS[22][30] )
         );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(n258), .D(n290), .Q(\REGISTERS[22][29] )
         );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(n258), .D(n293), .Q(\REGISTERS[22][28] )
         );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(n258), .D(n296), .Q(\REGISTERS[22][27] )
         );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(n258), .D(n299), .Q(\REGISTERS[22][26] )
         );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(n258), .D(n302), .Q(\REGISTERS[22][25] )
         );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(n258), .D(n305), .Q(\REGISTERS[22][24] )
         );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n258), .D(n308), .Q(\REGISTERS[22][23] )
         );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n258), .D(n311), .Q(\REGISTERS[22][22] )
         );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(n257), .D(n314), .Q(\REGISTERS[22][21] )
         );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(n257), .D(n317), .Q(\REGISTERS[22][20] )
         );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n257), .D(n320), .Q(\REGISTERS[22][19] )
         );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(n257), .D(n323), .Q(\REGISTERS[22][18] )
         );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n257), .D(n326), .Q(\REGISTERS[22][17] )
         );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(n257), .D(n329), .Q(\REGISTERS[22][16] )
         );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(n257), .D(n332), .Q(\REGISTERS[22][15] )
         );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(n257), .D(n335), .Q(\REGISTERS[22][14] )
         );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(n257), .D(n338), .Q(\REGISTERS[22][13] )
         );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(n257), .D(n341), .Q(\REGISTERS[22][12] )
         );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(n257), .D(n344), .Q(\REGISTERS[22][11] )
         );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n256), .D(n347), .Q(\REGISTERS[22][10] )
         );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(n256), .D(n350), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(n256), .D(n353), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n256), .D(n356), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(n256), .D(n359), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(n256), .D(n362), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(n256), .D(n365), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(n256), .D(n368), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(n256), .D(n371), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(n256), .D(n374), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(n256), .D(n377), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(n261), .D(n285), .Q(\REGISTERS[23][31] )
         );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(n261), .D(n288), .Q(\REGISTERS[23][30] )
         );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(n261), .D(n291), .Q(\REGISTERS[23][29] )
         );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(n261), .D(n294), .Q(\REGISTERS[23][28] )
         );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(n261), .D(n297), .Q(\REGISTERS[23][27] )
         );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(n261), .D(n300), .Q(\REGISTERS[23][26] )
         );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(n261), .D(n303), .Q(\REGISTERS[23][25] )
         );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(n261), .D(n306), .Q(\REGISTERS[23][24] )
         );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n261), .D(n309), .Q(\REGISTERS[23][23] )
         );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n261), .D(n312), .Q(\REGISTERS[23][22] )
         );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(n260), .D(n315), .Q(\REGISTERS[23][21] )
         );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(n260), .D(n318), .Q(\REGISTERS[23][20] )
         );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n260), .D(n321), .Q(\REGISTERS[23][19] )
         );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(n260), .D(n324), .Q(\REGISTERS[23][18] )
         );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n260), .D(n327), .Q(\REGISTERS[23][17] )
         );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(n260), .D(n330), .Q(\REGISTERS[23][16] )
         );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(n260), .D(n333), .Q(\REGISTERS[23][15] )
         );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(n260), .D(n336), .Q(\REGISTERS[23][14] )
         );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(n260), .D(n339), .Q(\REGISTERS[23][13] )
         );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(n260), .D(n342), .Q(\REGISTERS[23][12] )
         );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(n260), .D(n345), .Q(\REGISTERS[23][11] )
         );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n259), .D(n348), .Q(\REGISTERS[23][10] )
         );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(n259), .D(n351), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(n259), .D(n354), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n259), .D(n357), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(n259), .D(n360), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(n259), .D(n363), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(n259), .D(n366), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(n259), .D(n369), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(n259), .D(n372), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(n259), .D(n375), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(n259), .D(n378), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(n264), .D(n285), .Q(\REGISTERS[24][31] )
         );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(n264), .D(n288), .Q(\REGISTERS[24][30] )
         );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(n264), .D(n291), .Q(\REGISTERS[24][29] )
         );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(n264), .D(n294), .Q(\REGISTERS[24][28] )
         );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(n264), .D(n297), .Q(\REGISTERS[24][27] )
         );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(n264), .D(n300), .Q(\REGISTERS[24][26] )
         );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(n264), .D(n303), .Q(\REGISTERS[24][25] )
         );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n264), .D(n306), .Q(\REGISTERS[24][24] )
         );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n264), .D(n309), .Q(\REGISTERS[24][23] )
         );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(n264), .D(n312), .Q(\REGISTERS[24][22] )
         );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n263), .D(n315), .Q(\REGISTERS[24][21] )
         );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n263), .D(n318), .Q(\REGISTERS[24][20] )
         );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(n263), .D(n321), .Q(\REGISTERS[24][19] )
         );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(n263), .D(n324), .Q(\REGISTERS[24][18] )
         );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(n263), .D(n327), .Q(\REGISTERS[24][17] )
         );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(n263), .D(n330), .Q(\REGISTERS[24][16] )
         );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n263), .D(n333), .Q(\REGISTERS[24][15] )
         );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(n263), .D(n336), .Q(\REGISTERS[24][14] )
         );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(n263), .D(n339), .Q(\REGISTERS[24][13] )
         );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(n263), .D(n342), .Q(\REGISTERS[24][12] )
         );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(n263), .D(n345), .Q(\REGISTERS[24][11] )
         );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(n262), .D(n348), .Q(\REGISTERS[24][10] )
         );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(n262), .D(n351), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(n262), .D(n354), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(n262), .D(n357), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n262), .D(n360), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(n262), .D(n363), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(n262), .D(n366), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(n262), .D(n369), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(n262), .D(n372), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(n262), .D(n375), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(n262), .D(n378), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(n267), .D(n285), .Q(\REGISTERS[25][31] )
         );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(n267), .D(n288), .Q(\REGISTERS[25][30] )
         );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(n267), .D(n291), .Q(\REGISTERS[25][29] )
         );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(n267), .D(n294), .Q(\REGISTERS[25][28] )
         );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(n267), .D(n297), .Q(\REGISTERS[25][27] )
         );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(n267), .D(n300), .Q(\REGISTERS[25][26] )
         );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(n267), .D(n303), .Q(\REGISTERS[25][25] )
         );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(n267), .D(n306), .Q(\REGISTERS[25][24] )
         );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n267), .D(n309), .Q(\REGISTERS[25][23] )
         );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n267), .D(n312), .Q(\REGISTERS[25][22] )
         );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(n266), .D(n315), .Q(\REGISTERS[25][21] )
         );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(n266), .D(n318), .Q(\REGISTERS[25][20] )
         );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n266), .D(n321), .Q(\REGISTERS[25][19] )
         );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(n266), .D(n324), .Q(\REGISTERS[25][18] )
         );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n266), .D(n327), .Q(\REGISTERS[25][17] )
         );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(n266), .D(n330), .Q(\REGISTERS[25][16] )
         );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(n266), .D(n333), .Q(\REGISTERS[25][15] )
         );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(n266), .D(n336), .Q(\REGISTERS[25][14] )
         );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(n266), .D(n339), .Q(\REGISTERS[25][13] )
         );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(n266), .D(n342), .Q(\REGISTERS[25][12] )
         );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(n266), .D(n345), .Q(\REGISTERS[25][11] )
         );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n265), .D(n348), .Q(\REGISTERS[25][10] )
         );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(n265), .D(n351), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(n265), .D(n354), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n265), .D(n357), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(n265), .D(n360), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(n265), .D(n363), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(n265), .D(n366), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(n265), .D(n369), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(n265), .D(n372), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(n265), .D(n375), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(n265), .D(n378), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(n270), .D(n285), .Q(\REGISTERS[26][31] )
         );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(n270), .D(n288), .Q(\REGISTERS[26][30] )
         );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(n270), .D(n291), .Q(\REGISTERS[26][29] )
         );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(n270), .D(n294), .Q(\REGISTERS[26][28] )
         );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(n270), .D(n297), .Q(\REGISTERS[26][27] )
         );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(n270), .D(n300), .Q(\REGISTERS[26][26] )
         );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(n270), .D(n303), .Q(\REGISTERS[26][25] )
         );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(n270), .D(n306), .Q(\REGISTERS[26][24] )
         );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n270), .D(n309), .Q(\REGISTERS[26][23] )
         );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n270), .D(n312), .Q(\REGISTERS[26][22] )
         );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(n269), .D(n315), .Q(\REGISTERS[26][21] )
         );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(n269), .D(n318), .Q(\REGISTERS[26][20] )
         );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n269), .D(n321), .Q(\REGISTERS[26][19] )
         );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(n269), .D(n324), .Q(\REGISTERS[26][18] )
         );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n269), .D(n327), .Q(\REGISTERS[26][17] )
         );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(n269), .D(n330), .Q(\REGISTERS[26][16] )
         );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(n269), .D(n333), .Q(\REGISTERS[26][15] )
         );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(n269), .D(n336), .Q(\REGISTERS[26][14] )
         );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(n269), .D(n339), .Q(\REGISTERS[26][13] )
         );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(n269), .D(n342), .Q(\REGISTERS[26][12] )
         );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(n269), .D(n345), .Q(\REGISTERS[26][11] )
         );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n268), .D(n348), .Q(\REGISTERS[26][10] )
         );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(n268), .D(n351), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(n268), .D(n354), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n268), .D(n357), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(n268), .D(n360), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(n268), .D(n363), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(n268), .D(n366), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(n268), .D(n369), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(n268), .D(n372), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(n268), .D(n375), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(n268), .D(n378), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(n273), .D(n285), .Q(\REGISTERS[27][31] )
         );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(n273), .D(n288), .Q(\REGISTERS[27][30] )
         );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(n273), .D(n291), .Q(\REGISTERS[27][29] )
         );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(n273), .D(n294), .Q(\REGISTERS[27][28] )
         );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(n273), .D(n297), .Q(\REGISTERS[27][27] )
         );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(n273), .D(n300), .Q(\REGISTERS[27][26] )
         );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(n273), .D(n303), .Q(\REGISTERS[27][25] )
         );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(n273), .D(n306), .Q(\REGISTERS[27][24] )
         );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n273), .D(n309), .Q(\REGISTERS[27][23] )
         );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n273), .D(n312), .Q(\REGISTERS[27][22] )
         );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(n272), .D(n315), .Q(\REGISTERS[27][21] )
         );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(n272), .D(n318), .Q(\REGISTERS[27][20] )
         );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n272), .D(n321), .Q(\REGISTERS[27][19] )
         );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(n272), .D(n324), .Q(\REGISTERS[27][18] )
         );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n272), .D(n327), .Q(\REGISTERS[27][17] )
         );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(n272), .D(n330), .Q(\REGISTERS[27][16] )
         );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(n272), .D(n333), .Q(\REGISTERS[27][15] )
         );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(n272), .D(n336), .Q(\REGISTERS[27][14] )
         );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(n272), .D(n339), .Q(\REGISTERS[27][13] )
         );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(n272), .D(n342), .Q(\REGISTERS[27][12] )
         );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(n272), .D(n345), .Q(\REGISTERS[27][11] )
         );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n271), .D(n348), .Q(\REGISTERS[27][10] )
         );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(n271), .D(n351), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(n271), .D(n354), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n271), .D(n357), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(n271), .D(n360), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(n271), .D(n363), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(n271), .D(n366), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(n271), .D(n369), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(n271), .D(n372), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(n271), .D(n375), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(n271), .D(n378), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(n276), .D(n285), .Q(\REGISTERS[28][31] )
         );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(n276), .D(n288), .Q(\REGISTERS[28][30] )
         );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(n276), .D(n291), .Q(\REGISTERS[28][29] )
         );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(n276), .D(n294), .Q(\REGISTERS[28][28] )
         );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(n276), .D(n297), .Q(\REGISTERS[28][27] )
         );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(n276), .D(n300), .Q(\REGISTERS[28][26] )
         );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(n276), .D(n303), .Q(\REGISTERS[28][25] )
         );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(n276), .D(n306), .Q(\REGISTERS[28][24] )
         );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n276), .D(n309), .Q(\REGISTERS[28][23] )
         );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n276), .D(n312), .Q(\REGISTERS[28][22] )
         );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(n275), .D(n315), .Q(\REGISTERS[28][21] )
         );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(n275), .D(n318), .Q(\REGISTERS[28][20] )
         );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n275), .D(n321), .Q(\REGISTERS[28][19] )
         );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(n275), .D(n324), .Q(\REGISTERS[28][18] )
         );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n275), .D(n327), .Q(\REGISTERS[28][17] )
         );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(n275), .D(n330), .Q(\REGISTERS[28][16] )
         );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(n275), .D(n333), .Q(\REGISTERS[28][15] )
         );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(n275), .D(n336), .Q(\REGISTERS[28][14] )
         );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(n275), .D(n339), .Q(\REGISTERS[28][13] )
         );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(n275), .D(n342), .Q(\REGISTERS[28][12] )
         );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(n275), .D(n345), .Q(\REGISTERS[28][11] )
         );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n274), .D(n348), .Q(\REGISTERS[28][10] )
         );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(n274), .D(n351), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(n274), .D(n354), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n274), .D(n357), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(n274), .D(n360), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(n274), .D(n363), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(n274), .D(n366), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(n274), .D(n369), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(n274), .D(n372), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(n274), .D(n375), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(n274), .D(n378), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(n279), .D(n285), .Q(\REGISTERS[29][31] )
         );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(n279), .D(n288), .Q(\REGISTERS[29][30] )
         );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(n279), .D(n291), .Q(\REGISTERS[29][29] )
         );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(n279), .D(n294), .Q(\REGISTERS[29][28] )
         );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(n279), .D(n297), .Q(\REGISTERS[29][27] )
         );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(n279), .D(n300), .Q(\REGISTERS[29][26] )
         );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(n279), .D(n303), .Q(\REGISTERS[29][25] )
         );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(n279), .D(n306), .Q(\REGISTERS[29][24] )
         );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n279), .D(n309), .Q(\REGISTERS[29][23] )
         );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n279), .D(n312), .Q(\REGISTERS[29][22] )
         );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(n278), .D(n315), .Q(\REGISTERS[29][21] )
         );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(n278), .D(n318), .Q(\REGISTERS[29][20] )
         );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n278), .D(n321), .Q(\REGISTERS[29][19] )
         );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(n278), .D(n324), .Q(\REGISTERS[29][18] )
         );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n278), .D(n327), .Q(\REGISTERS[29][17] )
         );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(n278), .D(n330), .Q(\REGISTERS[29][16] )
         );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(n278), .D(n333), .Q(\REGISTERS[29][15] )
         );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(n278), .D(n336), .Q(\REGISTERS[29][14] )
         );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(n278), .D(n339), .Q(\REGISTERS[29][13] )
         );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(n278), .D(n342), .Q(\REGISTERS[29][12] )
         );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(n278), .D(n345), .Q(\REGISTERS[29][11] )
         );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n277), .D(n348), .Q(\REGISTERS[29][10] )
         );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(n277), .D(n351), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(n277), .D(n354), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n277), .D(n357), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(n277), .D(n360), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(n277), .D(n363), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(n277), .D(n366), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(n277), .D(n369), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(n277), .D(n372), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(n277), .D(n375), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(n277), .D(n378), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(n282), .D(n285), .Q(\REGISTERS[30][31] )
         );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(n282), .D(n288), .Q(\REGISTERS[30][30] )
         );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(n282), .D(n291), .Q(\REGISTERS[30][29] )
         );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(n282), .D(n294), .Q(\REGISTERS[30][28] )
         );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(n282), .D(n297), .Q(\REGISTERS[30][27] )
         );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(n282), .D(n300), .Q(\REGISTERS[30][26] )
         );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(n282), .D(n303), .Q(\REGISTERS[30][25] )
         );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(n282), .D(n306), .Q(\REGISTERS[30][24] )
         );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n282), .D(n309), .Q(\REGISTERS[30][23] )
         );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n282), .D(n312), .Q(\REGISTERS[30][22] )
         );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(n281), .D(n315), .Q(\REGISTERS[30][21] )
         );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(n281), .D(n318), .Q(\REGISTERS[30][20] )
         );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n281), .D(n321), .Q(\REGISTERS[30][19] )
         );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(n281), .D(n324), .Q(\REGISTERS[30][18] )
         );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n281), .D(n327), .Q(\REGISTERS[30][17] )
         );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(n281), .D(n330), .Q(\REGISTERS[30][16] )
         );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(n281), .D(n333), .Q(\REGISTERS[30][15] )
         );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(n281), .D(n336), .Q(\REGISTERS[30][14] )
         );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(n281), .D(n339), .Q(\REGISTERS[30][13] )
         );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(n281), .D(n342), .Q(\REGISTERS[30][12] )
         );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(n281), .D(n345), .Q(\REGISTERS[30][11] )
         );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n280), .D(n348), .Q(\REGISTERS[30][10] )
         );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(n280), .D(n351), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(n280), .D(n354), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n280), .D(n357), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(n280), .D(n360), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(n280), .D(n363), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(n280), .D(n366), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(n280), .D(n369), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(n280), .D(n372), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(n280), .D(n375), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(n280), .D(n378), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(n381), .D(n285), .Q(\REGISTERS[31][31] )
         );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(n381), .D(n288), .Q(\REGISTERS[31][30] )
         );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(n381), .D(n291), .Q(\REGISTERS[31][29] )
         );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(n381), .D(n294), .Q(\REGISTERS[31][28] )
         );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(n381), .D(n297), .Q(\REGISTERS[31][27] )
         );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(n381), .D(n300), .Q(\REGISTERS[31][26] )
         );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(n381), .D(n303), .Q(\REGISTERS[31][25] )
         );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(n381), .D(n306), .Q(\REGISTERS[31][24] )
         );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(n381), .D(n309), .Q(\REGISTERS[31][23] )
         );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(n381), .D(n312), .Q(\REGISTERS[31][22] )
         );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n380), .D(n315), .Q(\REGISTERS[31][21] )
         );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(n380), .D(n318), .Q(\REGISTERS[31][20] )
         );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n380), .D(n321), .Q(\REGISTERS[31][19] )
         );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(n380), .D(n324), .Q(\REGISTERS[31][18] )
         );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n380), .D(n327), .Q(\REGISTERS[31][17] )
         );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(n380), .D(n330), .Q(\REGISTERS[31][16] )
         );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(n380), .D(n333), .Q(\REGISTERS[31][15] )
         );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(n380), .D(n336), .Q(\REGISTERS[31][14] )
         );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(n380), .D(n339), .Q(\REGISTERS[31][13] )
         );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(n380), .D(n342), .Q(\REGISTERS[31][12] )
         );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n380), .D(n345), .Q(\REGISTERS[31][11] )
         );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n379), .D(n348), .Q(\REGISTERS[31][10] )
         );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(n379), .D(n351), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(n379), .D(n354), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(n379), .D(n357), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(n379), .D(n360), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(n379), .D(n363), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(n379), .D(n366), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(n379), .D(n369), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(n379), .D(n372), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(n379), .D(n375), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n379), .D(n378), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUTA_reg[31]  ( .G(n187), .D(N339), .Q(OUTA[31]) );
  DLH_X1 \OUTA_reg[30]  ( .G(n187), .D(N338), .Q(OUTA[30]) );
  DLH_X1 \OUTA_reg[29]  ( .G(n187), .D(N337), .Q(OUTA[29]) );
  DLH_X1 \OUTA_reg[28]  ( .G(n187), .D(N336), .Q(OUTA[28]) );
  DLH_X1 \OUTA_reg[27]  ( .G(n187), .D(N335), .Q(OUTA[27]) );
  DLH_X1 \OUTA_reg[26]  ( .G(n187), .D(N334), .Q(OUTA[26]) );
  DLH_X1 \OUTA_reg[25]  ( .G(n187), .D(N333), .Q(OUTA[25]) );
  DLH_X1 \OUTA_reg[24]  ( .G(n187), .D(N332), .Q(OUTA[24]) );
  DLH_X1 \OUTA_reg[23]  ( .G(n187), .D(N331), .Q(OUTA[23]) );
  DLH_X1 \OUTA_reg[22]  ( .G(n187), .D(N330), .Q(OUTA[22]) );
  DLH_X1 \OUTA_reg[21]  ( .G(n187), .D(N329), .Q(OUTA[21]) );
  DLH_X1 \OUTA_reg[20]  ( .G(n188), .D(N328), .Q(OUTA[20]) );
  DLH_X1 \OUTA_reg[19]  ( .G(n188), .D(N327), .Q(OUTA[19]) );
  DLH_X1 \OUTA_reg[18]  ( .G(n188), .D(N326), .Q(OUTA[18]) );
  DLH_X1 \OUTA_reg[17]  ( .G(n188), .D(N325), .Q(OUTA[17]) );
  DLH_X1 \OUTA_reg[16]  ( .G(n188), .D(N324), .Q(OUTA[16]) );
  DLH_X1 \OUTA_reg[15]  ( .G(n188), .D(N323), .Q(OUTA[15]) );
  DLH_X1 \OUTA_reg[14]  ( .G(n188), .D(N322), .Q(OUTA[14]) );
  DLH_X1 \OUTA_reg[13]  ( .G(n188), .D(N321), .Q(OUTA[13]) );
  DLH_X1 \OUTA_reg[12]  ( .G(n188), .D(N320), .Q(OUTA[12]) );
  DLH_X1 \OUTA_reg[11]  ( .G(n188), .D(N319), .Q(OUTA[11]) );
  DLH_X1 \OUTA_reg[10]  ( .G(n188), .D(N318), .Q(OUTA[10]) );
  DLH_X1 \OUTA_reg[9]  ( .G(n189), .D(N317), .Q(OUTA[9]) );
  DLH_X1 \OUTA_reg[8]  ( .G(n189), .D(N316), .Q(OUTA[8]) );
  DLH_X1 \OUTA_reg[7]  ( .G(n189), .D(N315), .Q(OUTA[7]) );
  DLH_X1 \OUTA_reg[6]  ( .G(n189), .D(N314), .Q(OUTA[6]) );
  DLH_X1 \OUTA_reg[5]  ( .G(n189), .D(N313), .Q(OUTA[5]) );
  DLH_X1 \OUTA_reg[4]  ( .G(n189), .D(N312), .Q(OUTA[4]) );
  DLH_X1 \OUTA_reg[3]  ( .G(n189), .D(N311), .Q(OUTA[3]) );
  DLH_X1 \OUTA_reg[2]  ( .G(n189), .D(N310), .Q(OUTA[2]) );
  DLH_X1 \OUTA_reg[1]  ( .G(n189), .D(N309), .Q(OUTA[1]) );
  DLH_X1 \OUTA_reg[0]  ( .G(n189), .D(N308), .Q(OUTA[0]) );
  DLH_X1 \OUTB_reg[31]  ( .G(n189), .D(N371), .Q(OUTB[31]) );
  DLH_X1 \OUTB_reg[30]  ( .G(n190), .D(N370), .Q(OUTB[30]) );
  DLH_X1 \OUTB_reg[29]  ( .G(n190), .D(N369), .Q(OUTB[29]) );
  DLH_X1 \OUTB_reg[28]  ( .G(n190), .D(N368), .Q(OUTB[28]) );
  DLH_X1 \OUTB_reg[27]  ( .G(n190), .D(N367), .Q(OUTB[27]) );
  DLH_X1 \OUTB_reg[26]  ( .G(n190), .D(N366), .Q(OUTB[26]) );
  DLH_X1 \OUTB_reg[25]  ( .G(n190), .D(N365), .Q(OUTB[25]) );
  DLH_X1 \OUTB_reg[24]  ( .G(n190), .D(N364), .Q(OUTB[24]) );
  DLH_X1 \OUTB_reg[23]  ( .G(n190), .D(N363), .Q(OUTB[23]) );
  DLH_X1 \OUTB_reg[22]  ( .G(n190), .D(N362), .Q(OUTB[22]) );
  DLH_X1 \OUTB_reg[21]  ( .G(n190), .D(N361), .Q(OUTB[21]) );
  DLH_X1 \OUTB_reg[20]  ( .G(n190), .D(N360), .Q(OUTB[20]) );
  DLH_X1 \OUTB_reg[19]  ( .G(n191), .D(N359), .Q(OUTB[19]) );
  DLH_X1 \OUTB_reg[18]  ( .G(n191), .D(N358), .Q(OUTB[18]) );
  DLH_X1 \OUTB_reg[17]  ( .G(n191), .D(N357), .Q(OUTB[17]) );
  DLH_X1 \OUTB_reg[16]  ( .G(n191), .D(N356), .Q(OUTB[16]) );
  DLH_X1 \OUTB_reg[15]  ( .G(n191), .D(N355), .Q(OUTB[15]) );
  DLH_X1 \OUTB_reg[14]  ( .G(n191), .D(N354), .Q(OUTB[14]) );
  DLH_X1 \OUTB_reg[13]  ( .G(n191), .D(N353), .Q(OUTB[13]) );
  DLH_X1 \OUTB_reg[12]  ( .G(n191), .D(N352), .Q(OUTB[12]) );
  DLH_X1 \OUTB_reg[11]  ( .G(n191), .D(N351), .Q(OUTB[11]) );
  DLH_X1 \OUTB_reg[10]  ( .G(n191), .D(N350), .Q(OUTB[10]) );
  DLH_X1 \OUTB_reg[9]  ( .G(n191), .D(N349), .Q(OUTB[9]) );
  DLH_X1 \OUTB_reg[8]  ( .G(n192), .D(N348), .Q(OUTB[8]) );
  DLH_X1 \OUTB_reg[7]  ( .G(n192), .D(N347), .Q(OUTB[7]) );
  DLH_X1 \OUTB_reg[6]  ( .G(n192), .D(N346), .Q(OUTB[6]) );
  DLH_X1 \OUTB_reg[5]  ( .G(n192), .D(N345), .Q(OUTB[5]) );
  DLH_X1 \OUTB_reg[4]  ( .G(n192), .D(N344), .Q(OUTB[4]) );
  DLH_X1 \OUTB_reg[3]  ( .G(n192), .D(N343), .Q(OUTB[3]) );
  DLH_X1 \OUTB_reg[2]  ( .G(n192), .D(N342), .Q(OUTB[2]) );
  DLH_X1 \OUTB_reg[1]  ( .G(n192), .D(N341), .Q(OUTB[1]) );
  DLH_X1 \OUTB_reg[0]  ( .G(n192), .D(N340), .Q(OUTB[0]) );
  NAND3_X1 U1905 ( .A1(n408), .A2(n407), .A3(WE), .ZN(n1775) );
  NAND3_X1 U1906 ( .A1(WE), .A2(n407), .A3(ADD_WR[3]), .ZN(n1783) );
  NAND3_X1 U1907 ( .A1(WE), .A2(n408), .A3(ADD_WR[4]), .ZN(n1785) );
  NAND3_X1 U1908 ( .A1(n410), .A2(n409), .A3(n411), .ZN(n1784) );
  NAND3_X1 U1909 ( .A1(n410), .A2(n409), .A3(ADD_WR[0]), .ZN(n1776) );
  NAND3_X1 U1910 ( .A1(n411), .A2(n409), .A3(ADD_WR[1]), .ZN(n1777) );
  NAND3_X1 U1911 ( .A1(ADD_WR[0]), .A2(n409), .A3(ADD_WR[1]), .ZN(n1778) );
  NAND3_X1 U1912 ( .A1(n411), .A2(n410), .A3(ADD_WR[2]), .ZN(n1779) );
  NAND3_X1 U1913 ( .A1(ADD_WR[0]), .A2(n410), .A3(ADD_WR[2]), .ZN(n1780) );
  NAND3_X1 U1914 ( .A1(ADD_WR[1]), .A2(n411), .A3(ADD_WR[2]), .ZN(n1781) );
  NAND3_X1 U1915 ( .A1(ADD_WR[3]), .A2(WE), .A3(ADD_WR[4]), .ZN(n1786) );
  NAND3_X1 U1916 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n1782)
         );
  NOR2_X1 U3 ( .A1(n2152), .A2(ADD_RDB[1]), .ZN(n1130) );
  NOR2_X1 U4 ( .A1(n2155), .A2(ADD_RDA[1]), .ZN(n1754) );
  BUF_X1 U5 ( .A(n542), .Z(n163) );
  BUF_X1 U6 ( .A(n566), .Z(n118) );
  BUF_X1 U7 ( .A(n576), .Z(n94) );
  BUF_X1 U8 ( .A(n542), .Z(n164) );
  BUF_X1 U9 ( .A(n566), .Z(n119) );
  BUF_X1 U10 ( .A(n576), .Z(n95) );
  BUF_X1 U11 ( .A(n542), .Z(n165) );
  BUF_X1 U12 ( .A(n566), .Z(n120) );
  BUF_X1 U13 ( .A(n576), .Z(n96) );
  BUF_X1 U14 ( .A(n549), .Z(n145) );
  BUF_X1 U15 ( .A(n549), .Z(n146) );
  BUF_X1 U16 ( .A(n549), .Z(n147) );
  BUF_X1 U17 ( .A(n536), .Z(n178) );
  BUF_X1 U18 ( .A(n541), .Z(n166) );
  BUF_X1 U19 ( .A(n546), .Z(n154) );
  BUF_X1 U20 ( .A(n551), .Z(n142) );
  BUF_X1 U21 ( .A(n570), .Z(n109) );
  BUF_X1 U22 ( .A(n565), .Z(n121) );
  BUF_X1 U23 ( .A(n575), .Z(n97) );
  BUF_X1 U24 ( .A(n560), .Z(n133) );
  BUF_X1 U25 ( .A(n536), .Z(n179) );
  BUF_X1 U26 ( .A(n541), .Z(n167) );
  BUF_X1 U27 ( .A(n546), .Z(n155) );
  BUF_X1 U28 ( .A(n551), .Z(n143) );
  BUF_X1 U29 ( .A(n570), .Z(n110) );
  BUF_X1 U30 ( .A(n565), .Z(n122) );
  BUF_X1 U31 ( .A(n575), .Z(n98) );
  BUF_X1 U32 ( .A(n560), .Z(n134) );
  BUF_X1 U33 ( .A(n533), .Z(n184) );
  BUF_X1 U34 ( .A(n538), .Z(n172) );
  BUF_X1 U35 ( .A(n543), .Z(n160) );
  BUF_X1 U36 ( .A(n548), .Z(n148) );
  BUF_X1 U37 ( .A(n567), .Z(n115) );
  BUF_X1 U38 ( .A(n562), .Z(n127) );
  BUF_X1 U39 ( .A(n572), .Z(n103) );
  BUF_X1 U40 ( .A(n533), .Z(n185) );
  BUF_X1 U41 ( .A(n538), .Z(n173) );
  BUF_X1 U42 ( .A(n543), .Z(n161) );
  BUF_X1 U43 ( .A(n548), .Z(n149) );
  BUF_X1 U44 ( .A(n567), .Z(n116) );
  BUF_X1 U45 ( .A(n562), .Z(n128) );
  BUF_X1 U46 ( .A(n572), .Z(n104) );
  BUF_X1 U47 ( .A(n537), .Z(n175) );
  BUF_X1 U48 ( .A(n547), .Z(n151) );
  BUF_X1 U49 ( .A(n552), .Z(n139) );
  BUF_X1 U50 ( .A(n571), .Z(n106) );
  BUF_X1 U51 ( .A(n561), .Z(n130) );
  BUF_X1 U52 ( .A(n537), .Z(n176) );
  BUF_X1 U53 ( .A(n547), .Z(n152) );
  BUF_X1 U54 ( .A(n552), .Z(n140) );
  BUF_X1 U55 ( .A(n571), .Z(n107) );
  BUF_X1 U56 ( .A(n561), .Z(n131) );
  BUF_X1 U57 ( .A(n1173), .Z(n52) );
  BUF_X1 U58 ( .A(n1173), .Z(n53) );
  BUF_X1 U59 ( .A(n533), .Z(n186) );
  BUF_X1 U60 ( .A(n538), .Z(n174) );
  BUF_X1 U61 ( .A(n567), .Z(n117) );
  BUF_X1 U62 ( .A(n562), .Z(n129) );
  BUF_X1 U63 ( .A(n572), .Z(n105) );
  BUF_X1 U64 ( .A(n536), .Z(n180) );
  BUF_X1 U65 ( .A(n541), .Z(n168) );
  BUF_X1 U66 ( .A(n546), .Z(n156) );
  BUF_X1 U67 ( .A(n551), .Z(n144) );
  BUF_X1 U68 ( .A(n570), .Z(n111) );
  BUF_X1 U69 ( .A(n565), .Z(n123) );
  BUF_X1 U70 ( .A(n575), .Z(n99) );
  BUF_X1 U71 ( .A(n560), .Z(n135) );
  BUF_X1 U72 ( .A(n543), .Z(n162) );
  BUF_X1 U73 ( .A(n548), .Z(n150) );
  BUF_X1 U74 ( .A(n557), .Z(n136) );
  BUF_X1 U75 ( .A(n557), .Z(n137) );
  BUF_X1 U76 ( .A(n537), .Z(n177) );
  BUF_X1 U77 ( .A(n547), .Z(n153) );
  BUF_X1 U78 ( .A(n552), .Z(n141) );
  BUF_X1 U79 ( .A(n571), .Z(n108) );
  BUF_X1 U80 ( .A(n561), .Z(n132) );
  BUF_X1 U81 ( .A(n534), .Z(n181) );
  BUF_X1 U82 ( .A(n539), .Z(n169) );
  BUF_X1 U83 ( .A(n544), .Z(n157) );
  BUF_X1 U84 ( .A(n568), .Z(n112) );
  BUF_X1 U85 ( .A(n563), .Z(n124) );
  BUF_X1 U86 ( .A(n573), .Z(n100) );
  BUF_X1 U87 ( .A(n534), .Z(n182) );
  BUF_X1 U88 ( .A(n539), .Z(n170) );
  BUF_X1 U89 ( .A(n544), .Z(n158) );
  BUF_X1 U90 ( .A(n568), .Z(n113) );
  BUF_X1 U91 ( .A(n563), .Z(n125) );
  BUF_X1 U92 ( .A(n573), .Z(n101) );
  BUF_X1 U93 ( .A(n1166), .Z(n71) );
  BUF_X1 U94 ( .A(n1190), .Z(n26) );
  BUF_X1 U95 ( .A(n1200), .Z(n2) );
  BUF_X1 U96 ( .A(n1166), .Z(n70) );
  BUF_X1 U97 ( .A(n1190), .Z(n25) );
  BUF_X1 U98 ( .A(n1200), .Z(n1) );
  BUF_X1 U99 ( .A(n1173), .Z(n54) );
  BUF_X1 U100 ( .A(n557), .Z(n138) );
  BUF_X1 U101 ( .A(n534), .Z(n183) );
  BUF_X1 U102 ( .A(n539), .Z(n171) );
  BUF_X1 U103 ( .A(n568), .Z(n114) );
  BUF_X1 U104 ( .A(n563), .Z(n126) );
  BUF_X1 U105 ( .A(n573), .Z(n102) );
  BUF_X1 U106 ( .A(n544), .Z(n159) );
  BUF_X1 U107 ( .A(n1166), .Z(n72) );
  BUF_X1 U108 ( .A(n1190), .Z(n27) );
  BUF_X1 U109 ( .A(n1200), .Z(n3) );
  NAND2_X1 U110 ( .A1(n1133), .A2(n1129), .ZN(n549) );
  AND2_X1 U111 ( .A1(n1124), .A2(n1129), .ZN(n542) );
  AND2_X1 U112 ( .A1(n1142), .A2(n1129), .ZN(n566) );
  AND2_X1 U113 ( .A1(n1147), .A2(n1129), .ZN(n576) );
  INV_X1 U114 ( .A(n406), .ZN(n390) );
  INV_X1 U115 ( .A(n406), .ZN(n389) );
  INV_X1 U116 ( .A(n406), .ZN(n393) );
  INV_X1 U117 ( .A(n406), .ZN(n392) );
  INV_X1 U118 ( .A(n406), .ZN(n391) );
  NOR2_X1 U119 ( .A1(n2152), .A2(n2151), .ZN(n1129) );
  BUF_X1 U120 ( .A(n1181), .Z(n43) );
  BUF_X1 U121 ( .A(n1181), .Z(n44) );
  BUF_X1 U122 ( .A(n1158), .Z(n88) );
  BUF_X1 U123 ( .A(n1163), .Z(n76) );
  BUF_X1 U124 ( .A(n1168), .Z(n64) );
  BUF_X1 U125 ( .A(n1187), .Z(n31) );
  BUF_X1 U126 ( .A(n1192), .Z(n19) );
  BUF_X1 U127 ( .A(n1197), .Z(n7) );
  BUF_X1 U128 ( .A(n1158), .Z(n89) );
  BUF_X1 U129 ( .A(n1163), .Z(n77) );
  BUF_X1 U130 ( .A(n1168), .Z(n65) );
  BUF_X1 U131 ( .A(n1187), .Z(n32) );
  BUF_X1 U132 ( .A(n1192), .Z(n20) );
  BUF_X1 U133 ( .A(n1197), .Z(n8) );
  BUF_X1 U134 ( .A(n1160), .Z(n85) );
  BUF_X1 U135 ( .A(n1165), .Z(n73) );
  BUF_X1 U136 ( .A(n1170), .Z(n61) );
  BUF_X1 U137 ( .A(n1175), .Z(n49) );
  BUF_X1 U138 ( .A(n1189), .Z(n28) );
  BUF_X1 U139 ( .A(n1194), .Z(n16) );
  BUF_X1 U140 ( .A(n1184), .Z(n40) );
  BUF_X1 U141 ( .A(n1199), .Z(n4) );
  BUF_X1 U142 ( .A(n1160), .Z(n86) );
  BUF_X1 U143 ( .A(n1165), .Z(n74) );
  BUF_X1 U144 ( .A(n1170), .Z(n62) );
  BUF_X1 U145 ( .A(n1175), .Z(n50) );
  BUF_X1 U146 ( .A(n1189), .Z(n29) );
  BUF_X1 U147 ( .A(n1194), .Z(n17) );
  BUF_X1 U148 ( .A(n1184), .Z(n41) );
  BUF_X1 U149 ( .A(n1199), .Z(n5) );
  BUF_X1 U150 ( .A(n1157), .Z(n91) );
  BUF_X1 U151 ( .A(n1162), .Z(n79) );
  BUF_X1 U152 ( .A(n1167), .Z(n67) );
  BUF_X1 U153 ( .A(n1172), .Z(n55) );
  BUF_X1 U154 ( .A(n1186), .Z(n34) );
  BUF_X1 U155 ( .A(n1191), .Z(n22) );
  BUF_X1 U156 ( .A(n1196), .Z(n10) );
  BUF_X1 U157 ( .A(n1157), .Z(n92) );
  BUF_X1 U158 ( .A(n1162), .Z(n80) );
  BUF_X1 U159 ( .A(n1167), .Z(n68) );
  BUF_X1 U160 ( .A(n1172), .Z(n56) );
  BUF_X1 U161 ( .A(n1186), .Z(n35) );
  BUF_X1 U162 ( .A(n1191), .Z(n23) );
  BUF_X1 U163 ( .A(n1196), .Z(n11) );
  BUF_X1 U164 ( .A(n1181), .Z(n45) );
  BUF_X1 U165 ( .A(n1161), .Z(n83) );
  BUF_X1 U166 ( .A(n1171), .Z(n59) );
  BUF_X1 U167 ( .A(n1176), .Z(n47) );
  BUF_X1 U168 ( .A(n1195), .Z(n14) );
  BUF_X1 U169 ( .A(n1185), .Z(n38) );
  BUF_X1 U170 ( .A(n1161), .Z(n82) );
  BUF_X1 U171 ( .A(n1171), .Z(n58) );
  BUF_X1 U172 ( .A(n1176), .Z(n46) );
  BUF_X1 U173 ( .A(n1195), .Z(n13) );
  BUF_X1 U174 ( .A(n1185), .Z(n37) );
  BUF_X1 U175 ( .A(n1158), .Z(n90) );
  BUF_X1 U176 ( .A(n1163), .Z(n78) );
  BUF_X1 U177 ( .A(n1168), .Z(n66) );
  BUF_X1 U178 ( .A(n1187), .Z(n33) );
  BUF_X1 U179 ( .A(n1192), .Z(n21) );
  BUF_X1 U180 ( .A(n1197), .Z(n9) );
  BUF_X1 U181 ( .A(n1160), .Z(n87) );
  BUF_X1 U182 ( .A(n1165), .Z(n75) );
  BUF_X1 U183 ( .A(n1170), .Z(n63) );
  BUF_X1 U184 ( .A(n1175), .Z(n51) );
  BUF_X1 U185 ( .A(n1189), .Z(n30) );
  BUF_X1 U186 ( .A(n1194), .Z(n18) );
  BUF_X1 U187 ( .A(n1184), .Z(n42) );
  BUF_X1 U188 ( .A(n1199), .Z(n6) );
  BUF_X1 U189 ( .A(n1157), .Z(n93) );
  BUF_X1 U190 ( .A(n1162), .Z(n81) );
  BUF_X1 U191 ( .A(n1167), .Z(n69) );
  BUF_X1 U192 ( .A(n1172), .Z(n57) );
  BUF_X1 U193 ( .A(n1186), .Z(n36) );
  BUF_X1 U194 ( .A(n1191), .Z(n24) );
  BUF_X1 U195 ( .A(n1196), .Z(n12) );
  BUF_X1 U196 ( .A(n1176), .Z(n48) );
  BUF_X1 U197 ( .A(n1161), .Z(n84) );
  BUF_X1 U198 ( .A(n1171), .Z(n60) );
  BUF_X1 U199 ( .A(n1195), .Z(n15) );
  BUF_X1 U200 ( .A(n1185), .Z(n39) );
  NAND2_X1 U201 ( .A1(n1127), .A2(n1134), .ZN(n543) );
  NAND2_X1 U202 ( .A1(n1127), .A2(n1133), .ZN(n544) );
  NAND2_X1 U203 ( .A1(n1129), .A2(n1134), .ZN(n548) );
  NAND2_X1 U204 ( .A1(n1126), .A2(n1130), .ZN(n538) );
  NAND2_X1 U205 ( .A1(n1124), .A2(n1130), .ZN(n539) );
  NAND2_X1 U206 ( .A1(n1143), .A2(n1130), .ZN(n562) );
  NAND2_X1 U207 ( .A1(n1142), .A2(n1130), .ZN(n563) );
  NAND2_X1 U208 ( .A1(n1148), .A2(n1130), .ZN(n572) );
  NAND2_X1 U209 ( .A1(n1147), .A2(n1130), .ZN(n573) );
  NAND2_X1 U210 ( .A1(n1126), .A2(n1127), .ZN(n533) );
  NAND2_X1 U211 ( .A1(n1124), .A2(n1127), .ZN(n534) );
  NAND2_X1 U212 ( .A1(n1148), .A2(n1127), .ZN(n567) );
  NAND2_X1 U213 ( .A1(n1147), .A2(n1127), .ZN(n568) );
  NAND2_X1 U214 ( .A1(n1143), .A2(n1127), .ZN(n557) );
  AND2_X1 U215 ( .A1(n1136), .A2(n2150), .ZN(n1133) );
  NAND2_X1 U216 ( .A1(n1757), .A2(n1753), .ZN(n1173) );
  AND2_X1 U217 ( .A1(n1150), .A2(n2150), .ZN(n1147) );
  AND2_X1 U218 ( .A1(n1131), .A2(n2150), .ZN(n1124) );
  AND2_X1 U219 ( .A1(n1130), .A2(n1133), .ZN(n552) );
  AND2_X1 U220 ( .A1(n1130), .A2(n1134), .ZN(n551) );
  AND2_X1 U221 ( .A1(n1125), .A2(n1133), .ZN(n547) );
  AND2_X1 U222 ( .A1(n1125), .A2(n1134), .ZN(n546) );
  AND2_X1 U223 ( .A1(n1126), .A2(n1129), .ZN(n541) );
  AND2_X1 U224 ( .A1(n1143), .A2(n1129), .ZN(n565) );
  AND2_X1 U225 ( .A1(n1148), .A2(n1129), .ZN(n575) );
  AND2_X1 U226 ( .A1(n1748), .A2(n1753), .ZN(n1166) );
  AND2_X1 U227 ( .A1(n1766), .A2(n1753), .ZN(n1190) );
  AND2_X1 U228 ( .A1(n1771), .A2(n1753), .ZN(n1200) );
  AND2_X1 U229 ( .A1(n1124), .A2(n1125), .ZN(n537) );
  AND2_X1 U230 ( .A1(n1126), .A2(n1125), .ZN(n536) );
  AND2_X1 U231 ( .A1(n1147), .A2(n1125), .ZN(n571) );
  AND2_X1 U232 ( .A1(n1148), .A2(n1125), .ZN(n570) );
  AND2_X1 U233 ( .A1(n1142), .A2(n1125), .ZN(n561) );
  AND2_X1 U234 ( .A1(n1143), .A2(n1125), .ZN(n560) );
  AND2_X1 U235 ( .A1(n1145), .A2(n2150), .ZN(n1142) );
  BUF_X1 U236 ( .A(n386), .Z(n406) );
  BUF_X1 U237 ( .A(n385), .Z(n405) );
  BUF_X1 U238 ( .A(n385), .Z(n404) );
  BUF_X1 U239 ( .A(n385), .Z(n403) );
  BUF_X1 U240 ( .A(n384), .Z(n402) );
  BUF_X1 U241 ( .A(n384), .Z(n401) );
  BUF_X1 U242 ( .A(n384), .Z(n400) );
  BUF_X1 U243 ( .A(n383), .Z(n399) );
  BUF_X1 U244 ( .A(n383), .Z(n397) );
  BUF_X1 U245 ( .A(n382), .Z(n396) );
  BUF_X1 U246 ( .A(n382), .Z(n395) );
  BUF_X1 U247 ( .A(n382), .Z(n394) );
  BUF_X1 U248 ( .A(n383), .Z(n398) );
  NOR2_X1 U249 ( .A1(ADD_RDB[1]), .A2(ADD_RDB[2]), .ZN(n1127) );
  NOR2_X1 U250 ( .A1(n2155), .A2(n2156), .ZN(n1753) );
  NOR2_X1 U251 ( .A1(n2151), .A2(ADD_RDB[2]), .ZN(n1125) );
  NAND2_X1 U252 ( .A1(n1751), .A2(n1757), .ZN(n1168) );
  NAND2_X1 U253 ( .A1(n1751), .A2(n1758), .ZN(n1167) );
  NAND2_X1 U254 ( .A1(n1753), .A2(n1758), .ZN(n1172) );
  NAND2_X1 U255 ( .A1(n1750), .A2(n1754), .ZN(n1162) );
  NAND2_X1 U256 ( .A1(n1748), .A2(n1754), .ZN(n1163) );
  NAND2_X1 U257 ( .A1(n1767), .A2(n1754), .ZN(n1186) );
  NAND2_X1 U258 ( .A1(n1766), .A2(n1754), .ZN(n1187) );
  NAND2_X1 U259 ( .A1(n1772), .A2(n1754), .ZN(n1196) );
  NAND2_X1 U260 ( .A1(n1771), .A2(n1754), .ZN(n1197) );
  NAND2_X1 U261 ( .A1(n1750), .A2(n1751), .ZN(n1157) );
  NAND2_X1 U262 ( .A1(n1748), .A2(n1751), .ZN(n1158) );
  NAND2_X1 U263 ( .A1(n1771), .A2(n1751), .ZN(n1192) );
  NAND2_X1 U264 ( .A1(n1772), .A2(n1751), .ZN(n1191) );
  NAND2_X1 U265 ( .A1(n1767), .A2(n1751), .ZN(n1181) );
  AND2_X1 U266 ( .A1(ADD_RDB[0]), .A2(n1136), .ZN(n1134) );
  AND2_X1 U267 ( .A1(n1760), .A2(n2157), .ZN(n1757) );
  NOR2_X1 U268 ( .A1(ADD_RDB[3]), .A2(ADD_RDB[4]), .ZN(n1145) );
  NOR2_X1 U269 ( .A1(n2153), .A2(ADD_RDB[4]), .ZN(n1150) );
  AND2_X1 U270 ( .A1(n1131), .A2(ADD_RDB[0]), .ZN(n1126) );
  AND2_X1 U271 ( .A1(n1150), .A2(ADD_RDB[0]), .ZN(n1148) );
  AND2_X1 U272 ( .A1(n1145), .A2(ADD_RDB[0]), .ZN(n1143) );
  AND2_X1 U273 ( .A1(n1774), .A2(n2157), .ZN(n1771) );
  AND2_X1 U274 ( .A1(n1755), .A2(n2157), .ZN(n1748) );
  AND2_X1 U275 ( .A1(n1754), .A2(n1757), .ZN(n1176) );
  AND2_X1 U276 ( .A1(n1754), .A2(n1758), .ZN(n1175) );
  AND2_X1 U277 ( .A1(n1749), .A2(n1757), .ZN(n1171) );
  AND2_X1 U278 ( .A1(n1749), .A2(n1758), .ZN(n1170) );
  AND2_X1 U279 ( .A1(n1750), .A2(n1753), .ZN(n1165) );
  AND2_X1 U280 ( .A1(n1767), .A2(n1753), .ZN(n1189) );
  AND2_X1 U281 ( .A1(n1772), .A2(n1753), .ZN(n1199) );
  AND2_X1 U282 ( .A1(n1750), .A2(n1749), .ZN(n1160) );
  AND2_X1 U283 ( .A1(n1748), .A2(n1749), .ZN(n1161) );
  AND2_X1 U284 ( .A1(n1771), .A2(n1749), .ZN(n1195) );
  AND2_X1 U285 ( .A1(n1772), .A2(n1749), .ZN(n1194) );
  AND2_X1 U286 ( .A1(n1766), .A2(n1749), .ZN(n1185) );
  AND2_X1 U287 ( .A1(n1767), .A2(n1749), .ZN(n1184) );
  INV_X1 U288 ( .A(ADD_RDB[0]), .ZN(n2150) );
  AND2_X1 U289 ( .A1(n1769), .A2(n2157), .ZN(n1766) );
  INV_X1 U290 ( .A(ADD_RDB[1]), .ZN(n2151) );
  INV_X1 U291 ( .A(ADD_RDB[2]), .ZN(n2152) );
  AND2_X1 U292 ( .A1(ADD_RDB[4]), .A2(ADD_RDB[3]), .ZN(n1136) );
  AND2_X1 U293 ( .A1(ADD_RDB[4]), .A2(n2153), .ZN(n1131) );
  INV_X1 U294 ( .A(ADD_RDB[3]), .ZN(n2153) );
  BUF_X1 U295 ( .A(N298), .Z(n214) );
  BUF_X1 U296 ( .A(N298), .Z(n215) );
  BUF_X1 U297 ( .A(N299), .Z(n211) );
  BUF_X1 U298 ( .A(N299), .Z(n212) );
  BUF_X1 U299 ( .A(N300), .Z(n208) );
  BUF_X1 U300 ( .A(N300), .Z(n209) );
  BUF_X1 U301 ( .A(N301), .Z(n205) );
  BUF_X1 U302 ( .A(N301), .Z(n206) );
  BUF_X1 U303 ( .A(N302), .Z(n202) );
  BUF_X1 U304 ( .A(N302), .Z(n203) );
  BUF_X1 U305 ( .A(N303), .Z(n199) );
  BUF_X1 U306 ( .A(N303), .Z(n200) );
  BUF_X1 U307 ( .A(N304), .Z(n196) );
  BUF_X1 U308 ( .A(N304), .Z(n197) );
  BUF_X1 U309 ( .A(N305), .Z(n193) );
  BUF_X1 U310 ( .A(N305), .Z(n194) );
  BUF_X1 U311 ( .A(N243), .Z(n379) );
  BUF_X1 U312 ( .A(N243), .Z(n380) );
  BUF_X1 U313 ( .A(N276), .Z(n280) );
  BUF_X1 U314 ( .A(N276), .Z(n281) );
  BUF_X1 U315 ( .A(N277), .Z(n277) );
  BUF_X1 U316 ( .A(N277), .Z(n278) );
  BUF_X1 U317 ( .A(N278), .Z(n274) );
  BUF_X1 U318 ( .A(N278), .Z(n275) );
  BUF_X1 U319 ( .A(N279), .Z(n271) );
  BUF_X1 U320 ( .A(N279), .Z(n272) );
  BUF_X1 U321 ( .A(N280), .Z(n268) );
  BUF_X1 U322 ( .A(N280), .Z(n269) );
  BUF_X1 U323 ( .A(N281), .Z(n265) );
  BUF_X1 U324 ( .A(N281), .Z(n266) );
  BUF_X1 U325 ( .A(N282), .Z(n262) );
  BUF_X1 U326 ( .A(N282), .Z(n263) );
  BUF_X1 U327 ( .A(N283), .Z(n259) );
  BUF_X1 U328 ( .A(N283), .Z(n260) );
  BUF_X1 U329 ( .A(N284), .Z(n256) );
  BUF_X1 U330 ( .A(N284), .Z(n257) );
  BUF_X1 U331 ( .A(N285), .Z(n253) );
  BUF_X1 U332 ( .A(N285), .Z(n254) );
  BUF_X1 U333 ( .A(N286), .Z(n250) );
  BUF_X1 U334 ( .A(N286), .Z(n251) );
  BUF_X1 U335 ( .A(N287), .Z(n247) );
  BUF_X1 U336 ( .A(N287), .Z(n248) );
  BUF_X1 U337 ( .A(N288), .Z(n244) );
  BUF_X1 U338 ( .A(N288), .Z(n245) );
  BUF_X1 U339 ( .A(N289), .Z(n241) );
  BUF_X1 U340 ( .A(N289), .Z(n242) );
  BUF_X1 U341 ( .A(N290), .Z(n238) );
  BUF_X1 U342 ( .A(N290), .Z(n239) );
  BUF_X1 U343 ( .A(N291), .Z(n235) );
  BUF_X1 U344 ( .A(N291), .Z(n236) );
  BUF_X1 U345 ( .A(N292), .Z(n232) );
  BUF_X1 U346 ( .A(N292), .Z(n233) );
  BUF_X1 U347 ( .A(N293), .Z(n229) );
  BUF_X1 U348 ( .A(N293), .Z(n230) );
  BUF_X1 U349 ( .A(N294), .Z(n226) );
  BUF_X1 U350 ( .A(N294), .Z(n227) );
  BUF_X1 U351 ( .A(N295), .Z(n223) );
  BUF_X1 U352 ( .A(N295), .Z(n224) );
  BUF_X1 U353 ( .A(N296), .Z(n220) );
  BUF_X1 U354 ( .A(N296), .Z(n221) );
  BUF_X1 U355 ( .A(N297), .Z(n217) );
  BUF_X1 U356 ( .A(N297), .Z(n218) );
  BUF_X1 U357 ( .A(N298), .Z(n216) );
  BUF_X1 U358 ( .A(N299), .Z(n213) );
  BUF_X1 U359 ( .A(N300), .Z(n210) );
  BUF_X1 U360 ( .A(N301), .Z(n207) );
  BUF_X1 U361 ( .A(N302), .Z(n204) );
  BUF_X1 U362 ( .A(N303), .Z(n201) );
  BUF_X1 U363 ( .A(N304), .Z(n198) );
  BUF_X1 U364 ( .A(N305), .Z(n195) );
  BUF_X1 U365 ( .A(N243), .Z(n381) );
  BUF_X1 U366 ( .A(N276), .Z(n282) );
  BUF_X1 U367 ( .A(N277), .Z(n279) );
  BUF_X1 U368 ( .A(N278), .Z(n276) );
  BUF_X1 U369 ( .A(N279), .Z(n273) );
  BUF_X1 U370 ( .A(N280), .Z(n270) );
  BUF_X1 U371 ( .A(N281), .Z(n267) );
  BUF_X1 U372 ( .A(N282), .Z(n264) );
  BUF_X1 U373 ( .A(N283), .Z(n261) );
  BUF_X1 U374 ( .A(N284), .Z(n258) );
  BUF_X1 U375 ( .A(N285), .Z(n255) );
  BUF_X1 U376 ( .A(N286), .Z(n252) );
  BUF_X1 U377 ( .A(N287), .Z(n249) );
  BUF_X1 U378 ( .A(N288), .Z(n246) );
  BUF_X1 U379 ( .A(N289), .Z(n243) );
  BUF_X1 U380 ( .A(N290), .Z(n240) );
  BUF_X1 U381 ( .A(N291), .Z(n237) );
  BUF_X1 U382 ( .A(N292), .Z(n234) );
  BUF_X1 U383 ( .A(N293), .Z(n231) );
  BUF_X1 U384 ( .A(N294), .Z(n228) );
  BUF_X1 U385 ( .A(N295), .Z(n225) );
  BUF_X1 U386 ( .A(N296), .Z(n222) );
  BUF_X1 U387 ( .A(N297), .Z(n219) );
  BUF_X1 U388 ( .A(n387), .Z(n385) );
  BUF_X1 U389 ( .A(n387), .Z(n384) );
  BUF_X1 U390 ( .A(n388), .Z(n382) );
  BUF_X1 U391 ( .A(n388), .Z(n383) );
  BUF_X1 U392 ( .A(n387), .Z(n386) );
  NOR2_X1 U393 ( .A1(ADD_RDA[1]), .A2(ADD_RDA[2]), .ZN(n1751) );
  NOR2_X1 U394 ( .A1(n2156), .A2(ADD_RDA[2]), .ZN(n1749) );
  AND2_X1 U395 ( .A1(ADD_RDA[0]), .A2(n1760), .ZN(n1758) );
  NOR2_X1 U396 ( .A1(ADD_RDA[3]), .A2(ADD_RDA[4]), .ZN(n1769) );
  AOI21_X1 U397 ( .B1(n1117), .B2(n1118), .A(n391), .ZN(N340) );
  NOR4_X1 U398 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1117) );
  NOR4_X1 U399 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
  OAI21_X1 U400 ( .B1(n136), .B2(n443), .A(n1141), .ZN(n1140) );
  AOI21_X1 U401 ( .B1(n1099), .B2(n1100), .A(n391), .ZN(N341) );
  NOR4_X1 U402 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1099) );
  NOR4_X1 U403 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
  OAI21_X1 U404 ( .B1(n136), .B2(n442), .A(n1113), .ZN(n1112) );
  AOI21_X1 U405 ( .B1(n1081), .B2(n1082), .A(n391), .ZN(N342) );
  NOR4_X1 U406 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1081) );
  NOR4_X1 U407 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
  OAI21_X1 U408 ( .B1(n136), .B2(n441), .A(n1095), .ZN(n1094) );
  AOI21_X1 U409 ( .B1(n1063), .B2(n1064), .A(n391), .ZN(N343) );
  NOR4_X1 U410 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1063) );
  NOR4_X1 U411 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
  OAI21_X1 U412 ( .B1(n136), .B2(n440), .A(n1077), .ZN(n1076) );
  AOI21_X1 U413 ( .B1(n1045), .B2(n1046), .A(n391), .ZN(N344) );
  NOR4_X1 U414 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1045) );
  NOR4_X1 U415 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
  OAI21_X1 U416 ( .B1(n136), .B2(n439), .A(n1059), .ZN(n1058) );
  AOI21_X1 U417 ( .B1(n1027), .B2(n1028), .A(n391), .ZN(N345) );
  NOR4_X1 U418 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1027) );
  NOR4_X1 U419 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
  OAI21_X1 U420 ( .B1(n136), .B2(n438), .A(n1041), .ZN(n1040) );
  AOI21_X1 U421 ( .B1(n1009), .B2(n1010), .A(n391), .ZN(N346) );
  NOR4_X1 U422 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1009) );
  NOR4_X1 U423 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
  OAI21_X1 U424 ( .B1(n136), .B2(n437), .A(n1023), .ZN(n1022) );
  AOI21_X1 U425 ( .B1(n991), .B2(n992), .A(n391), .ZN(N347) );
  NOR4_X1 U426 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n991) );
  NOR4_X1 U427 ( .A1(n993), .A2(n994), .A3(n995), .A4(n996), .ZN(n992) );
  OAI21_X1 U428 ( .B1(n136), .B2(n436), .A(n1005), .ZN(n1004) );
  AOI21_X1 U429 ( .B1(n973), .B2(n974), .A(n390), .ZN(N348) );
  NOR4_X1 U430 ( .A1(n983), .A2(n984), .A3(n985), .A4(n986), .ZN(n973) );
  NOR4_X1 U431 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n974) );
  OAI21_X1 U432 ( .B1(n136), .B2(n435), .A(n987), .ZN(n986) );
  AOI21_X1 U433 ( .B1(n955), .B2(n956), .A(n390), .ZN(N349) );
  NOR4_X1 U434 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n955) );
  NOR4_X1 U435 ( .A1(n957), .A2(n958), .A3(n959), .A4(n960), .ZN(n956) );
  OAI21_X1 U436 ( .B1(n136), .B2(n434), .A(n969), .ZN(n968) );
  AOI21_X1 U437 ( .B1(n937), .B2(n938), .A(n390), .ZN(N350) );
  NOR4_X1 U438 ( .A1(n947), .A2(n948), .A3(n949), .A4(n950), .ZN(n937) );
  NOR4_X1 U439 ( .A1(n939), .A2(n940), .A3(n941), .A4(n942), .ZN(n938) );
  OAI21_X1 U440 ( .B1(n136), .B2(n433), .A(n951), .ZN(n950) );
  AOI21_X1 U441 ( .B1(n919), .B2(n920), .A(n390), .ZN(N351) );
  NOR4_X1 U442 ( .A1(n929), .A2(n930), .A3(n931), .A4(n932), .ZN(n919) );
  NOR4_X1 U443 ( .A1(n921), .A2(n922), .A3(n923), .A4(n924), .ZN(n920) );
  OAI21_X1 U444 ( .B1(n136), .B2(n432), .A(n933), .ZN(n932) );
  AOI21_X1 U445 ( .B1(n901), .B2(n902), .A(n390), .ZN(N352) );
  NOR4_X1 U446 ( .A1(n911), .A2(n912), .A3(n913), .A4(n914), .ZN(n901) );
  NOR4_X1 U447 ( .A1(n903), .A2(n904), .A3(n905), .A4(n906), .ZN(n902) );
  OAI21_X1 U448 ( .B1(n137), .B2(n431), .A(n915), .ZN(n914) );
  AOI21_X1 U449 ( .B1(n883), .B2(n884), .A(n390), .ZN(N353) );
  NOR4_X1 U450 ( .A1(n893), .A2(n894), .A3(n895), .A4(n896), .ZN(n883) );
  NOR4_X1 U451 ( .A1(n885), .A2(n886), .A3(n887), .A4(n888), .ZN(n884) );
  OAI21_X1 U452 ( .B1(n137), .B2(n430), .A(n897), .ZN(n896) );
  AOI21_X1 U453 ( .B1(n865), .B2(n866), .A(n390), .ZN(N354) );
  NOR4_X1 U454 ( .A1(n875), .A2(n876), .A3(n877), .A4(n878), .ZN(n865) );
  NOR4_X1 U455 ( .A1(n867), .A2(n868), .A3(n869), .A4(n870), .ZN(n866) );
  OAI21_X1 U456 ( .B1(n137), .B2(n429), .A(n879), .ZN(n878) );
  AOI21_X1 U457 ( .B1(n847), .B2(n848), .A(n390), .ZN(N355) );
  NOR4_X1 U458 ( .A1(n857), .A2(n858), .A3(n859), .A4(n860), .ZN(n847) );
  NOR4_X1 U459 ( .A1(n849), .A2(n850), .A3(n851), .A4(n852), .ZN(n848) );
  OAI21_X1 U460 ( .B1(n137), .B2(n428), .A(n861), .ZN(n860) );
  AOI21_X1 U461 ( .B1(n829), .B2(n830), .A(n390), .ZN(N356) );
  NOR4_X1 U462 ( .A1(n839), .A2(n840), .A3(n841), .A4(n842), .ZN(n829) );
  NOR4_X1 U463 ( .A1(n831), .A2(n832), .A3(n833), .A4(n834), .ZN(n830) );
  OAI21_X1 U464 ( .B1(n137), .B2(n427), .A(n843), .ZN(n842) );
  AOI21_X1 U465 ( .B1(n811), .B2(n812), .A(n390), .ZN(N357) );
  NOR4_X1 U466 ( .A1(n821), .A2(n822), .A3(n823), .A4(n824), .ZN(n811) );
  NOR4_X1 U467 ( .A1(n813), .A2(n814), .A3(n815), .A4(n816), .ZN(n812) );
  OAI21_X1 U468 ( .B1(n137), .B2(n426), .A(n825), .ZN(n824) );
  AOI21_X1 U469 ( .B1(n793), .B2(n794), .A(n390), .ZN(N358) );
  NOR4_X1 U470 ( .A1(n803), .A2(n804), .A3(n805), .A4(n806), .ZN(n793) );
  NOR4_X1 U471 ( .A1(n795), .A2(n796), .A3(n797), .A4(n798), .ZN(n794) );
  OAI21_X1 U472 ( .B1(n137), .B2(n425), .A(n807), .ZN(n806) );
  AOI21_X1 U473 ( .B1(n775), .B2(n776), .A(n390), .ZN(N359) );
  NOR4_X1 U474 ( .A1(n785), .A2(n786), .A3(n787), .A4(n788), .ZN(n775) );
  NOR4_X1 U475 ( .A1(n777), .A2(n778), .A3(n779), .A4(n780), .ZN(n776) );
  OAI21_X1 U476 ( .B1(n137), .B2(n424), .A(n789), .ZN(n788) );
  AOI21_X1 U477 ( .B1(n757), .B2(n758), .A(n389), .ZN(N360) );
  NOR4_X1 U478 ( .A1(n767), .A2(n768), .A3(n769), .A4(n770), .ZN(n757) );
  NOR4_X1 U479 ( .A1(n759), .A2(n760), .A3(n761), .A4(n762), .ZN(n758) );
  OAI21_X1 U480 ( .B1(n137), .B2(n423), .A(n771), .ZN(n770) );
  AOI21_X1 U481 ( .B1(n739), .B2(n740), .A(n389), .ZN(N361) );
  NOR4_X1 U482 ( .A1(n749), .A2(n750), .A3(n751), .A4(n752), .ZN(n739) );
  NOR4_X1 U483 ( .A1(n741), .A2(n742), .A3(n743), .A4(n744), .ZN(n740) );
  OAI21_X1 U484 ( .B1(n137), .B2(n422), .A(n753), .ZN(n752) );
  AOI21_X1 U485 ( .B1(n721), .B2(n722), .A(n389), .ZN(N362) );
  NOR4_X1 U486 ( .A1(n731), .A2(n732), .A3(n733), .A4(n734), .ZN(n721) );
  NOR4_X1 U487 ( .A1(n723), .A2(n724), .A3(n725), .A4(n726), .ZN(n722) );
  OAI21_X1 U488 ( .B1(n137), .B2(n421), .A(n735), .ZN(n734) );
  AOI21_X1 U489 ( .B1(n703), .B2(n704), .A(n389), .ZN(N363) );
  NOR4_X1 U490 ( .A1(n713), .A2(n714), .A3(n715), .A4(n716), .ZN(n703) );
  NOR4_X1 U491 ( .A1(n705), .A2(n706), .A3(n707), .A4(n708), .ZN(n704) );
  OAI21_X1 U492 ( .B1(n137), .B2(n420), .A(n717), .ZN(n716) );
  AOI21_X1 U493 ( .B1(n685), .B2(n686), .A(n389), .ZN(N364) );
  NOR4_X1 U494 ( .A1(n695), .A2(n696), .A3(n697), .A4(n698), .ZN(n685) );
  NOR4_X1 U495 ( .A1(n687), .A2(n688), .A3(n689), .A4(n690), .ZN(n686) );
  OAI21_X1 U496 ( .B1(n138), .B2(n419), .A(n699), .ZN(n698) );
  AOI21_X1 U497 ( .B1(n667), .B2(n668), .A(n389), .ZN(N365) );
  NOR4_X1 U498 ( .A1(n677), .A2(n678), .A3(n679), .A4(n680), .ZN(n667) );
  NOR4_X1 U499 ( .A1(n669), .A2(n670), .A3(n671), .A4(n672), .ZN(n668) );
  OAI21_X1 U500 ( .B1(n138), .B2(n418), .A(n681), .ZN(n680) );
  AOI21_X1 U501 ( .B1(n649), .B2(n650), .A(n389), .ZN(N366) );
  NOR4_X1 U502 ( .A1(n659), .A2(n660), .A3(n661), .A4(n662), .ZN(n649) );
  NOR4_X1 U503 ( .A1(n651), .A2(n652), .A3(n653), .A4(n654), .ZN(n650) );
  OAI21_X1 U504 ( .B1(n138), .B2(n417), .A(n663), .ZN(n662) );
  AOI21_X1 U505 ( .B1(n631), .B2(n632), .A(n389), .ZN(N367) );
  NOR4_X1 U506 ( .A1(n641), .A2(n642), .A3(n643), .A4(n644), .ZN(n631) );
  NOR4_X1 U507 ( .A1(n633), .A2(n634), .A3(n635), .A4(n636), .ZN(n632) );
  OAI21_X1 U508 ( .B1(n138), .B2(n416), .A(n645), .ZN(n644) );
  AOI21_X1 U509 ( .B1(n613), .B2(n614), .A(n389), .ZN(N368) );
  NOR4_X1 U510 ( .A1(n623), .A2(n624), .A3(n625), .A4(n626), .ZN(n613) );
  NOR4_X1 U511 ( .A1(n615), .A2(n616), .A3(n617), .A4(n618), .ZN(n614) );
  OAI21_X1 U512 ( .B1(n138), .B2(n415), .A(n627), .ZN(n626) );
  AOI21_X1 U513 ( .B1(n595), .B2(n596), .A(n389), .ZN(N369) );
  NOR4_X1 U514 ( .A1(n605), .A2(n606), .A3(n607), .A4(n608), .ZN(n595) );
  NOR4_X1 U515 ( .A1(n597), .A2(n598), .A3(n599), .A4(n600), .ZN(n596) );
  OAI21_X1 U516 ( .B1(n138), .B2(n414), .A(n609), .ZN(n608) );
  AOI21_X1 U517 ( .B1(n577), .B2(n578), .A(n389), .ZN(N370) );
  NOR4_X1 U518 ( .A1(n587), .A2(n588), .A3(n589), .A4(n590), .ZN(n577) );
  NOR4_X1 U519 ( .A1(n579), .A2(n580), .A3(n581), .A4(n582), .ZN(n578) );
  OAI21_X1 U520 ( .B1(n138), .B2(n413), .A(n591), .ZN(n590) );
  AOI21_X1 U521 ( .B1(n527), .B2(n528), .A(n389), .ZN(N371) );
  NOR4_X1 U522 ( .A1(n553), .A2(n554), .A3(n555), .A4(n556), .ZN(n527) );
  NOR4_X1 U523 ( .A1(n529), .A2(n530), .A3(n531), .A4(n532), .ZN(n528) );
  OAI21_X1 U524 ( .B1(n138), .B2(n412), .A(n559), .ZN(n556) );
  AOI21_X1 U525 ( .B1(n1669), .B2(n1670), .A(n393), .ZN(N312) );
  NOR4_X1 U526 ( .A1(n1679), .A2(n1680), .A3(n1681), .A4(n1682), .ZN(n1669) );
  NOR4_X1 U527 ( .A1(n1671), .A2(n1672), .A3(n1673), .A4(n1674), .ZN(n1670) );
  OAI221_X1 U528 ( .B1(n1889), .B2(n10), .C1(n1857), .C2(n7), .A(n1686), .ZN(
        n1679) );
  AOI21_X1 U529 ( .B1(n1651), .B2(n1652), .A(n393), .ZN(N313) );
  NOR4_X1 U530 ( .A1(n1661), .A2(n1662), .A3(n1663), .A4(n1664), .ZN(n1651) );
  NOR4_X1 U531 ( .A1(n1653), .A2(n1654), .A3(n1655), .A4(n1656), .ZN(n1652) );
  OAI221_X1 U532 ( .B1(n1888), .B2(n10), .C1(n1856), .C2(n7), .A(n1668), .ZN(
        n1661) );
  AOI21_X1 U533 ( .B1(n1633), .B2(n1634), .A(n393), .ZN(N314) );
  NOR4_X1 U534 ( .A1(n1643), .A2(n1644), .A3(n1645), .A4(n1646), .ZN(n1633) );
  NOR4_X1 U535 ( .A1(n1635), .A2(n1636), .A3(n1637), .A4(n1638), .ZN(n1634) );
  OAI221_X1 U536 ( .B1(n1887), .B2(n10), .C1(n1855), .C2(n7), .A(n1650), .ZN(
        n1643) );
  AOI21_X1 U537 ( .B1(n1615), .B2(n1616), .A(n393), .ZN(N315) );
  NOR4_X1 U538 ( .A1(n1625), .A2(n1626), .A3(n1627), .A4(n1628), .ZN(n1615) );
  NOR4_X1 U539 ( .A1(n1617), .A2(n1618), .A3(n1619), .A4(n1620), .ZN(n1616) );
  OAI221_X1 U540 ( .B1(n1886), .B2(n10), .C1(n1854), .C2(n7), .A(n1632), .ZN(
        n1625) );
  AOI21_X1 U541 ( .B1(n1597), .B2(n1598), .A(n393), .ZN(N316) );
  NOR4_X1 U542 ( .A1(n1607), .A2(n1608), .A3(n1609), .A4(n1610), .ZN(n1597) );
  NOR4_X1 U543 ( .A1(n1599), .A2(n1600), .A3(n1601), .A4(n1602), .ZN(n1598) );
  OAI221_X1 U544 ( .B1(n1885), .B2(n10), .C1(n1853), .C2(n7), .A(n1614), .ZN(
        n1607) );
  AOI21_X1 U545 ( .B1(n1579), .B2(n1580), .A(n393), .ZN(N317) );
  NOR4_X1 U546 ( .A1(n1589), .A2(n1590), .A3(n1591), .A4(n1592), .ZN(n1579) );
  NOR4_X1 U547 ( .A1(n1581), .A2(n1582), .A3(n1583), .A4(n1584), .ZN(n1580) );
  OAI221_X1 U548 ( .B1(n1884), .B2(n10), .C1(n1852), .C2(n7), .A(n1596), .ZN(
        n1589) );
  AOI21_X1 U549 ( .B1(n1561), .B2(n1562), .A(n393), .ZN(N318) );
  NOR4_X1 U550 ( .A1(n1571), .A2(n1572), .A3(n1573), .A4(n1574), .ZN(n1561) );
  NOR4_X1 U551 ( .A1(n1563), .A2(n1564), .A3(n1565), .A4(n1566), .ZN(n1562) );
  OAI221_X1 U552 ( .B1(n1883), .B2(n10), .C1(n1851), .C2(n7), .A(n1578), .ZN(
        n1571) );
  AOI21_X1 U553 ( .B1(n1543), .B2(n1544), .A(n393), .ZN(N319) );
  NOR4_X1 U554 ( .A1(n1553), .A2(n1554), .A3(n1555), .A4(n1556), .ZN(n1543) );
  NOR4_X1 U555 ( .A1(n1545), .A2(n1546), .A3(n1547), .A4(n1548), .ZN(n1544) );
  OAI221_X1 U556 ( .B1(n1882), .B2(n10), .C1(n1850), .C2(n7), .A(n1560), .ZN(
        n1553) );
  AOI21_X1 U557 ( .B1(n1525), .B2(n1526), .A(n393), .ZN(N320) );
  NOR4_X1 U558 ( .A1(n1535), .A2(n1536), .A3(n1537), .A4(n1538), .ZN(n1525) );
  NOR4_X1 U559 ( .A1(n1527), .A2(n1528), .A3(n1529), .A4(n1530), .ZN(n1526) );
  OAI221_X1 U560 ( .B1(n1881), .B2(n11), .C1(n1849), .C2(n8), .A(n1542), .ZN(
        n1535) );
  AOI21_X1 U561 ( .B1(n1507), .B2(n1508), .A(n393), .ZN(N321) );
  NOR4_X1 U562 ( .A1(n1517), .A2(n1518), .A3(n1519), .A4(n1520), .ZN(n1507) );
  NOR4_X1 U563 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .ZN(n1508) );
  OAI221_X1 U564 ( .B1(n1880), .B2(n11), .C1(n1848), .C2(n8), .A(n1524), .ZN(
        n1517) );
  AOI21_X1 U565 ( .B1(n1489), .B2(n1490), .A(n393), .ZN(N322) );
  NOR4_X1 U566 ( .A1(n1499), .A2(n1500), .A3(n1501), .A4(n1502), .ZN(n1489) );
  NOR4_X1 U567 ( .A1(n1491), .A2(n1492), .A3(n1493), .A4(n1494), .ZN(n1490) );
  OAI221_X1 U568 ( .B1(n1879), .B2(n11), .C1(n1847), .C2(n8), .A(n1506), .ZN(
        n1499) );
  AOI21_X1 U569 ( .B1(n1471), .B2(n1472), .A(n393), .ZN(N323) );
  NOR4_X1 U570 ( .A1(n1481), .A2(n1482), .A3(n1483), .A4(n1484), .ZN(n1471) );
  NOR4_X1 U571 ( .A1(n1473), .A2(n1474), .A3(n1475), .A4(n1476), .ZN(n1472) );
  OAI221_X1 U572 ( .B1(n1878), .B2(n11), .C1(n1846), .C2(n8), .A(n1488), .ZN(
        n1481) );
  AOI21_X1 U573 ( .B1(n1453), .B2(n1454), .A(n392), .ZN(N324) );
  NOR4_X1 U574 ( .A1(n1463), .A2(n1464), .A3(n1465), .A4(n1466), .ZN(n1453) );
  NOR4_X1 U575 ( .A1(n1455), .A2(n1456), .A3(n1457), .A4(n1458), .ZN(n1454) );
  OAI221_X1 U576 ( .B1(n1877), .B2(n11), .C1(n1845), .C2(n8), .A(n1470), .ZN(
        n1463) );
  AOI21_X1 U577 ( .B1(n1435), .B2(n1436), .A(n392), .ZN(N325) );
  NOR4_X1 U578 ( .A1(n1445), .A2(n1446), .A3(n1447), .A4(n1448), .ZN(n1435) );
  NOR4_X1 U579 ( .A1(n1437), .A2(n1438), .A3(n1439), .A4(n1440), .ZN(n1436) );
  OAI221_X1 U580 ( .B1(n1876), .B2(n11), .C1(n1844), .C2(n8), .A(n1452), .ZN(
        n1445) );
  AOI21_X1 U581 ( .B1(n1417), .B2(n1418), .A(n392), .ZN(N326) );
  NOR4_X1 U582 ( .A1(n1427), .A2(n1428), .A3(n1429), .A4(n1430), .ZN(n1417) );
  NOR4_X1 U583 ( .A1(n1419), .A2(n1420), .A3(n1421), .A4(n1422), .ZN(n1418) );
  OAI221_X1 U584 ( .B1(n1875), .B2(n11), .C1(n1843), .C2(n8), .A(n1434), .ZN(
        n1427) );
  AOI21_X1 U585 ( .B1(n1399), .B2(n1400), .A(n392), .ZN(N327) );
  NOR4_X1 U586 ( .A1(n1409), .A2(n1410), .A3(n1411), .A4(n1412), .ZN(n1399) );
  NOR4_X1 U587 ( .A1(n1401), .A2(n1402), .A3(n1403), .A4(n1404), .ZN(n1400) );
  OAI221_X1 U588 ( .B1(n1874), .B2(n11), .C1(n1842), .C2(n8), .A(n1416), .ZN(
        n1409) );
  AOI21_X1 U589 ( .B1(n1381), .B2(n1382), .A(n392), .ZN(N328) );
  NOR4_X1 U590 ( .A1(n1391), .A2(n1392), .A3(n1393), .A4(n1394), .ZN(n1381) );
  NOR4_X1 U591 ( .A1(n1383), .A2(n1384), .A3(n1385), .A4(n1386), .ZN(n1382) );
  OAI221_X1 U592 ( .B1(n1873), .B2(n11), .C1(n1841), .C2(n8), .A(n1398), .ZN(
        n1391) );
  AOI21_X1 U593 ( .B1(n1363), .B2(n1364), .A(n392), .ZN(N329) );
  NOR4_X1 U594 ( .A1(n1373), .A2(n1374), .A3(n1375), .A4(n1376), .ZN(n1363) );
  NOR4_X1 U595 ( .A1(n1365), .A2(n1366), .A3(n1367), .A4(n1368), .ZN(n1364) );
  OAI221_X1 U596 ( .B1(n1872), .B2(n11), .C1(n1840), .C2(n8), .A(n1380), .ZN(
        n1373) );
  AOI21_X1 U597 ( .B1(n1345), .B2(n1346), .A(n392), .ZN(N330) );
  NOR4_X1 U598 ( .A1(n1355), .A2(n1356), .A3(n1357), .A4(n1358), .ZN(n1345) );
  NOR4_X1 U599 ( .A1(n1347), .A2(n1348), .A3(n1349), .A4(n1350), .ZN(n1346) );
  OAI221_X1 U600 ( .B1(n1871), .B2(n11), .C1(n1839), .C2(n8), .A(n1362), .ZN(
        n1355) );
  AOI21_X1 U601 ( .B1(n1327), .B2(n1328), .A(n392), .ZN(N331) );
  NOR4_X1 U602 ( .A1(n1337), .A2(n1338), .A3(n1339), .A4(n1340), .ZN(n1327) );
  NOR4_X1 U603 ( .A1(n1329), .A2(n1330), .A3(n1331), .A4(n1332), .ZN(n1328) );
  OAI221_X1 U604 ( .B1(n1870), .B2(n11), .C1(n1838), .C2(n8), .A(n1344), .ZN(
        n1337) );
  AOI21_X1 U605 ( .B1(n1309), .B2(n1310), .A(n392), .ZN(N332) );
  NOR4_X1 U606 ( .A1(n1319), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1309) );
  NOR4_X1 U607 ( .A1(n1311), .A2(n1312), .A3(n1313), .A4(n1314), .ZN(n1310) );
  OAI221_X1 U608 ( .B1(n1869), .B2(n12), .C1(n1837), .C2(n9), .A(n1326), .ZN(
        n1319) );
  AOI21_X1 U609 ( .B1(n1291), .B2(n1292), .A(n392), .ZN(N333) );
  NOR4_X1 U610 ( .A1(n1301), .A2(n1302), .A3(n1303), .A4(n1304), .ZN(n1291) );
  NOR4_X1 U611 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1292) );
  OAI221_X1 U612 ( .B1(n1868), .B2(n12), .C1(n1836), .C2(n9), .A(n1308), .ZN(
        n1301) );
  AOI21_X1 U613 ( .B1(n1273), .B2(n1274), .A(n392), .ZN(N334) );
  NOR4_X1 U614 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1273) );
  NOR4_X1 U615 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1274) );
  OAI221_X1 U616 ( .B1(n1867), .B2(n12), .C1(n1835), .C2(n9), .A(n1290), .ZN(
        n1283) );
  AOI21_X1 U617 ( .B1(n1255), .B2(n1256), .A(n392), .ZN(N335) );
  NOR4_X1 U618 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1255) );
  NOR4_X1 U619 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1256) );
  OAI221_X1 U620 ( .B1(n1866), .B2(n12), .C1(n1834), .C2(n9), .A(n1272), .ZN(
        n1265) );
  AOI21_X1 U621 ( .B1(n1237), .B2(n1238), .A(n391), .ZN(N336) );
  NOR4_X1 U622 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1237) );
  NOR4_X1 U623 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1238) );
  OAI221_X1 U624 ( .B1(n1865), .B2(n12), .C1(n1833), .C2(n9), .A(n1254), .ZN(
        n1247) );
  AOI21_X1 U625 ( .B1(n1219), .B2(n1220), .A(n391), .ZN(N337) );
  NOR4_X1 U626 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1219) );
  NOR4_X1 U627 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
  OAI221_X1 U628 ( .B1(n1864), .B2(n12), .C1(n1832), .C2(n9), .A(n1236), .ZN(
        n1229) );
  AOI21_X1 U629 ( .B1(n1201), .B2(n1202), .A(n391), .ZN(N338) );
  NOR4_X1 U630 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1201) );
  NOR4_X1 U631 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
  OAI221_X1 U632 ( .B1(n1863), .B2(n12), .C1(n1831), .C2(n9), .A(n1218), .ZN(
        n1211) );
  AOI21_X1 U633 ( .B1(n1151), .B2(n1152), .A(n391), .ZN(N339) );
  NOR4_X1 U634 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1151) );
  NOR4_X1 U635 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1152) );
  OAI221_X1 U636 ( .B1(n1862), .B2(n12), .C1(n1830), .C2(n9), .A(n1198), .ZN(
        n1177) );
  NOR2_X1 U637 ( .A1(n2154), .A2(ADD_RDA[4]), .ZN(n1774) );
  AND2_X1 U638 ( .A1(n1755), .A2(ADD_RDA[0]), .ZN(n1750) );
  AND2_X1 U639 ( .A1(n1774), .A2(ADD_RDA[0]), .ZN(n1772) );
  AND2_X1 U640 ( .A1(n1769), .A2(ADD_RDA[0]), .ZN(n1767) );
  AOI21_X1 U641 ( .B1(n1741), .B2(n1742), .A(n390), .ZN(N308) );
  NOR4_X1 U642 ( .A1(n1761), .A2(n1762), .A3(n1763), .A4(n1764), .ZN(n1741) );
  NOR4_X1 U643 ( .A1(n1743), .A2(n1744), .A3(n1745), .A4(n1746), .ZN(n1742) );
  OAI221_X1 U644 ( .B1(n1893), .B2(n10), .C1(n1861), .C2(n7), .A(n1773), .ZN(
        n1761) );
  AOI21_X1 U645 ( .B1(n1723), .B2(n1724), .A(n389), .ZN(N309) );
  NOR4_X1 U646 ( .A1(n1733), .A2(n1734), .A3(n1735), .A4(n1736), .ZN(n1723) );
  NOR4_X1 U647 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(n1724) );
  OAI221_X1 U648 ( .B1(n1892), .B2(n10), .C1(n1860), .C2(n7), .A(n1740), .ZN(
        n1733) );
  AOI21_X1 U649 ( .B1(n1705), .B2(n1706), .A(n393), .ZN(N310) );
  NOR4_X1 U650 ( .A1(n1715), .A2(n1716), .A3(n1717), .A4(n1718), .ZN(n1705) );
  NOR4_X1 U651 ( .A1(n1707), .A2(n1708), .A3(n1709), .A4(n1710), .ZN(n1706) );
  OAI221_X1 U652 ( .B1(n1891), .B2(n10), .C1(n1859), .C2(n7), .A(n1722), .ZN(
        n1715) );
  AOI21_X1 U653 ( .B1(n1687), .B2(n1688), .A(n392), .ZN(N311) );
  NOR4_X1 U654 ( .A1(n1697), .A2(n1698), .A3(n1699), .A4(n1700), .ZN(n1687) );
  NOR4_X1 U655 ( .A1(n1689), .A2(n1690), .A3(n1691), .A4(n1692), .ZN(n1688) );
  OAI221_X1 U656 ( .B1(n1890), .B2(n10), .C1(n1858), .C2(n7), .A(n1704), .ZN(
        n1697) );
  INV_X1 U657 ( .A(ADD_RDA[0]), .ZN(n2157) );
  INV_X1 U658 ( .A(ADD_RDA[1]), .ZN(n2156) );
  INV_X1 U659 ( .A(ADD_RDA[2]), .ZN(n2155) );
  INV_X1 U660 ( .A(ADD_RDA[3]), .ZN(n2154) );
  AND2_X1 U661 ( .A1(ADD_RDA[4]), .A2(ADD_RDA[3]), .ZN(n1760) );
  AND2_X1 U662 ( .A1(ADD_RDA[4]), .A2(n2154), .ZN(n1755) );
  OAI21_X1 U663 ( .B1(n1783), .B2(n1784), .A(n395), .ZN(N298) );
  OAI21_X1 U664 ( .B1(n1775), .B2(n1782), .A(n395), .ZN(N299) );
  OAI21_X1 U665 ( .B1(n1775), .B2(n1781), .A(n395), .ZN(N300) );
  OAI21_X1 U666 ( .B1(n1775), .B2(n1780), .A(n394), .ZN(N301) );
  OAI21_X1 U667 ( .B1(n1775), .B2(n1779), .A(n394), .ZN(N302) );
  OAI21_X1 U668 ( .B1(n1775), .B2(n1778), .A(n394), .ZN(N303) );
  OAI21_X1 U669 ( .B1(n1775), .B2(n1777), .A(n394), .ZN(N304) );
  OAI21_X1 U670 ( .B1(n1775), .B2(n1776), .A(n398), .ZN(N305) );
  OAI21_X1 U671 ( .B1(n1782), .B2(n1786), .A(n395), .ZN(N243) );
  OAI21_X1 U672 ( .B1(n1781), .B2(n1786), .A(n401), .ZN(N276) );
  OAI21_X1 U673 ( .B1(n1780), .B2(n1786), .A(n401), .ZN(N277) );
  OAI21_X1 U674 ( .B1(n1779), .B2(n1786), .A(n401), .ZN(N278) );
  OAI21_X1 U675 ( .B1(n1778), .B2(n1786), .A(n400), .ZN(N279) );
  OAI21_X1 U676 ( .B1(n1777), .B2(n1786), .A(n400), .ZN(N280) );
  OAI21_X1 U677 ( .B1(n1776), .B2(n1786), .A(n400), .ZN(N281) );
  OAI21_X1 U678 ( .B1(n1784), .B2(n1786), .A(n400), .ZN(N282) );
  OAI21_X1 U679 ( .B1(n1782), .B2(n1785), .A(n399), .ZN(N283) );
  OAI21_X1 U680 ( .B1(n1781), .B2(n1785), .A(n399), .ZN(N284) );
  OAI21_X1 U681 ( .B1(n1780), .B2(n1785), .A(n399), .ZN(N285) );
  OAI21_X1 U682 ( .B1(n1779), .B2(n1785), .A(n399), .ZN(N286) );
  OAI21_X1 U683 ( .B1(n1778), .B2(n1785), .A(n398), .ZN(N287) );
  OAI21_X1 U684 ( .B1(n1777), .B2(n1785), .A(n398), .ZN(N288) );
  OAI21_X1 U685 ( .B1(n1776), .B2(n1785), .A(n398), .ZN(N289) );
  OAI21_X1 U686 ( .B1(n1784), .B2(n1785), .A(n397), .ZN(N290) );
  OAI21_X1 U687 ( .B1(n1782), .B2(n1783), .A(n397), .ZN(N291) );
  OAI21_X1 U688 ( .B1(n1781), .B2(n1783), .A(n397), .ZN(N292) );
  OAI21_X1 U689 ( .B1(n1780), .B2(n1783), .A(n397), .ZN(N293) );
  OAI21_X1 U690 ( .B1(n1779), .B2(n1783), .A(n396), .ZN(N294) );
  OAI21_X1 U691 ( .B1(n1778), .B2(n1783), .A(n396), .ZN(N295) );
  OAI21_X1 U692 ( .B1(n1777), .B2(n1783), .A(n396), .ZN(N296) );
  OAI21_X1 U693 ( .B1(n1776), .B2(n1783), .A(n396), .ZN(N297) );
  BUF_X1 U694 ( .A(N244), .Z(n377) );
  BUF_X1 U695 ( .A(N245), .Z(n374) );
  BUF_X1 U696 ( .A(N246), .Z(n371) );
  BUF_X1 U697 ( .A(N247), .Z(n368) );
  BUF_X1 U698 ( .A(N248), .Z(n365) );
  BUF_X1 U699 ( .A(N249), .Z(n362) );
  BUF_X1 U700 ( .A(N250), .Z(n359) );
  BUF_X1 U701 ( .A(N251), .Z(n356) );
  BUF_X1 U702 ( .A(N252), .Z(n353) );
  BUF_X1 U703 ( .A(N253), .Z(n350) );
  BUF_X1 U704 ( .A(N254), .Z(n347) );
  BUF_X1 U705 ( .A(N255), .Z(n344) );
  BUF_X1 U706 ( .A(N256), .Z(n341) );
  BUF_X1 U707 ( .A(N257), .Z(n338) );
  BUF_X1 U708 ( .A(N258), .Z(n335) );
  BUF_X1 U709 ( .A(N259), .Z(n332) );
  BUF_X1 U710 ( .A(N260), .Z(n329) );
  BUF_X1 U711 ( .A(N261), .Z(n326) );
  BUF_X1 U712 ( .A(N262), .Z(n323) );
  BUF_X1 U713 ( .A(N263), .Z(n320) );
  BUF_X1 U714 ( .A(N264), .Z(n317) );
  BUF_X1 U715 ( .A(N265), .Z(n314) );
  BUF_X1 U716 ( .A(N266), .Z(n311) );
  BUF_X1 U717 ( .A(N267), .Z(n308) );
  BUF_X1 U718 ( .A(N268), .Z(n305) );
  BUF_X1 U719 ( .A(N269), .Z(n302) );
  BUF_X1 U720 ( .A(N270), .Z(n299) );
  BUF_X1 U721 ( .A(N271), .Z(n296) );
  BUF_X1 U722 ( .A(N272), .Z(n293) );
  BUF_X1 U723 ( .A(N273), .Z(n290) );
  BUF_X1 U724 ( .A(N274), .Z(n287) );
  BUF_X1 U725 ( .A(N275), .Z(n284) );
  BUF_X1 U726 ( .A(N244), .Z(n376) );
  BUF_X1 U727 ( .A(N245), .Z(n373) );
  BUF_X1 U728 ( .A(N246), .Z(n370) );
  BUF_X1 U729 ( .A(N247), .Z(n367) );
  BUF_X1 U730 ( .A(N248), .Z(n364) );
  BUF_X1 U731 ( .A(N249), .Z(n361) );
  BUF_X1 U732 ( .A(N250), .Z(n358) );
  BUF_X1 U733 ( .A(N251), .Z(n355) );
  BUF_X1 U734 ( .A(N252), .Z(n352) );
  BUF_X1 U735 ( .A(N253), .Z(n349) );
  BUF_X1 U736 ( .A(N254), .Z(n346) );
  BUF_X1 U737 ( .A(N255), .Z(n343) );
  BUF_X1 U738 ( .A(N256), .Z(n340) );
  BUF_X1 U739 ( .A(N257), .Z(n337) );
  BUF_X1 U740 ( .A(N258), .Z(n334) );
  BUF_X1 U741 ( .A(N259), .Z(n331) );
  BUF_X1 U742 ( .A(N260), .Z(n328) );
  BUF_X1 U743 ( .A(N261), .Z(n325) );
  BUF_X1 U744 ( .A(N262), .Z(n322) );
  BUF_X1 U745 ( .A(N263), .Z(n319) );
  BUF_X1 U746 ( .A(N264), .Z(n316) );
  BUF_X1 U747 ( .A(N265), .Z(n313) );
  BUF_X1 U748 ( .A(N266), .Z(n310) );
  BUF_X1 U749 ( .A(N267), .Z(n307) );
  BUF_X1 U750 ( .A(N268), .Z(n304) );
  BUF_X1 U751 ( .A(N269), .Z(n301) );
  BUF_X1 U752 ( .A(N270), .Z(n298) );
  BUF_X1 U753 ( .A(N271), .Z(n295) );
  BUF_X1 U754 ( .A(N272), .Z(n292) );
  BUF_X1 U755 ( .A(N273), .Z(n289) );
  BUF_X1 U756 ( .A(N274), .Z(n286) );
  BUF_X1 U757 ( .A(N275), .Z(n283) );
  BUF_X1 U758 ( .A(N244), .Z(n378) );
  BUF_X1 U759 ( .A(N245), .Z(n375) );
  BUF_X1 U760 ( .A(N246), .Z(n372) );
  BUF_X1 U761 ( .A(N247), .Z(n369) );
  BUF_X1 U762 ( .A(N248), .Z(n366) );
  BUF_X1 U763 ( .A(N249), .Z(n363) );
  BUF_X1 U764 ( .A(N250), .Z(n360) );
  BUF_X1 U765 ( .A(N251), .Z(n357) );
  BUF_X1 U766 ( .A(N252), .Z(n354) );
  BUF_X1 U767 ( .A(N253), .Z(n351) );
  BUF_X1 U768 ( .A(N254), .Z(n348) );
  BUF_X1 U769 ( .A(N255), .Z(n345) );
  BUF_X1 U770 ( .A(N256), .Z(n342) );
  BUF_X1 U771 ( .A(N257), .Z(n339) );
  BUF_X1 U772 ( .A(N258), .Z(n336) );
  BUF_X1 U773 ( .A(N259), .Z(n333) );
  BUF_X1 U774 ( .A(N260), .Z(n330) );
  BUF_X1 U775 ( .A(N261), .Z(n327) );
  BUF_X1 U776 ( .A(N262), .Z(n324) );
  BUF_X1 U777 ( .A(N263), .Z(n321) );
  BUF_X1 U778 ( .A(N264), .Z(n318) );
  BUF_X1 U779 ( .A(N265), .Z(n315) );
  BUF_X1 U780 ( .A(N266), .Z(n312) );
  BUF_X1 U781 ( .A(N267), .Z(n309) );
  BUF_X1 U782 ( .A(N268), .Z(n306) );
  BUF_X1 U783 ( .A(N269), .Z(n303) );
  BUF_X1 U784 ( .A(N270), .Z(n300) );
  BUF_X1 U785 ( .A(N271), .Z(n297) );
  BUF_X1 U786 ( .A(N272), .Z(n294) );
  BUF_X1 U787 ( .A(N273), .Z(n291) );
  BUF_X1 U788 ( .A(N274), .Z(n288) );
  BUF_X1 U789 ( .A(N275), .Z(n285) );
  BUF_X1 U790 ( .A(RESET), .Z(n387) );
  BUF_X1 U791 ( .A(RESET), .Z(n388) );
  OAI221_X1 U792 ( .B1(n1933), .B2(n93), .C1(n1901), .C2(n90), .A(n1315), .ZN(
        n1314) );
  AOI22_X1 U793 ( .A1(n87), .A2(\REGISTERS[19][24] ), .B1(n82), .B2(
        \REGISTERS[18][24] ), .ZN(n1315) );
  OAI221_X1 U794 ( .B1(n1932), .B2(n93), .C1(n1900), .C2(n90), .A(n1297), .ZN(
        n1296) );
  AOI22_X1 U795 ( .A1(n87), .A2(\REGISTERS[19][25] ), .B1(n82), .B2(
        \REGISTERS[18][25] ), .ZN(n1297) );
  OAI221_X1 U796 ( .B1(n1931), .B2(n93), .C1(n1899), .C2(n90), .A(n1279), .ZN(
        n1278) );
  AOI22_X1 U797 ( .A1(n87), .A2(\REGISTERS[19][26] ), .B1(n82), .B2(
        \REGISTERS[18][26] ), .ZN(n1279) );
  OAI221_X1 U798 ( .B1(n1930), .B2(n93), .C1(n1898), .C2(n90), .A(n1261), .ZN(
        n1260) );
  AOI22_X1 U799 ( .A1(n87), .A2(\REGISTERS[19][27] ), .B1(n82), .B2(
        \REGISTERS[18][27] ), .ZN(n1261) );
  OAI221_X1 U800 ( .B1(n1929), .B2(n93), .C1(n1897), .C2(n90), .A(n1243), .ZN(
        n1242) );
  AOI22_X1 U801 ( .A1(n87), .A2(\REGISTERS[19][28] ), .B1(n82), .B2(
        \REGISTERS[18][28] ), .ZN(n1243) );
  OAI221_X1 U802 ( .B1(n1928), .B2(n93), .C1(n1896), .C2(n90), .A(n1225), .ZN(
        n1224) );
  AOI22_X1 U803 ( .A1(n87), .A2(\REGISTERS[19][29] ), .B1(n82), .B2(
        \REGISTERS[18][29] ), .ZN(n1225) );
  OAI221_X1 U804 ( .B1(n1927), .B2(n93), .C1(n1895), .C2(n90), .A(n1207), .ZN(
        n1206) );
  AOI22_X1 U805 ( .A1(n87), .A2(\REGISTERS[19][30] ), .B1(n82), .B2(
        \REGISTERS[18][30] ), .ZN(n1207) );
  OAI221_X1 U806 ( .B1(n1926), .B2(n93), .C1(n1894), .C2(n90), .A(n1159), .ZN(
        n1156) );
  AOI22_X1 U807 ( .A1(n87), .A2(\REGISTERS[19][31] ), .B1(n82), .B2(
        \REGISTERS[18][31] ), .ZN(n1159) );
  OAI221_X1 U808 ( .B1(n1997), .B2(n81), .C1(n1965), .C2(n78), .A(n1316), .ZN(
        n1313) );
  AOI22_X1 U809 ( .A1(n75), .A2(\REGISTERS[23][24] ), .B1(n70), .B2(
        \REGISTERS[22][24] ), .ZN(n1316) );
  OAI221_X1 U810 ( .B1(n483), .B2(n36), .C1(n451), .C2(n33), .A(n1324), .ZN(
        n1321) );
  AOI22_X1 U811 ( .A1(n30), .A2(\REGISTERS[7][24] ), .B1(n25), .B2(
        \REGISTERS[6][24] ), .ZN(n1324) );
  OAI221_X1 U812 ( .B1(n1996), .B2(n81), .C1(n1964), .C2(n78), .A(n1298), .ZN(
        n1295) );
  AOI22_X1 U813 ( .A1(n75), .A2(\REGISTERS[23][25] ), .B1(n70), .B2(
        \REGISTERS[22][25] ), .ZN(n1298) );
  OAI221_X1 U814 ( .B1(n482), .B2(n36), .C1(n450), .C2(n33), .A(n1306), .ZN(
        n1303) );
  AOI22_X1 U815 ( .A1(n30), .A2(\REGISTERS[7][25] ), .B1(n25), .B2(
        \REGISTERS[6][25] ), .ZN(n1306) );
  OAI221_X1 U816 ( .B1(n1995), .B2(n81), .C1(n1963), .C2(n78), .A(n1280), .ZN(
        n1277) );
  AOI22_X1 U817 ( .A1(n75), .A2(\REGISTERS[23][26] ), .B1(n70), .B2(
        \REGISTERS[22][26] ), .ZN(n1280) );
  OAI221_X1 U818 ( .B1(n481), .B2(n36), .C1(n449), .C2(n33), .A(n1288), .ZN(
        n1285) );
  AOI22_X1 U819 ( .A1(n30), .A2(\REGISTERS[7][26] ), .B1(n25), .B2(
        \REGISTERS[6][26] ), .ZN(n1288) );
  OAI221_X1 U820 ( .B1(n1994), .B2(n81), .C1(n1962), .C2(n78), .A(n1262), .ZN(
        n1259) );
  AOI22_X1 U821 ( .A1(n75), .A2(\REGISTERS[23][27] ), .B1(n70), .B2(
        \REGISTERS[22][27] ), .ZN(n1262) );
  OAI221_X1 U822 ( .B1(n480), .B2(n36), .C1(n448), .C2(n33), .A(n1270), .ZN(
        n1267) );
  AOI22_X1 U823 ( .A1(n30), .A2(\REGISTERS[7][27] ), .B1(n25), .B2(
        \REGISTERS[6][27] ), .ZN(n1270) );
  OAI221_X1 U824 ( .B1(n1993), .B2(n81), .C1(n1961), .C2(n78), .A(n1244), .ZN(
        n1241) );
  AOI22_X1 U825 ( .A1(n75), .A2(\REGISTERS[23][28] ), .B1(n70), .B2(
        \REGISTERS[22][28] ), .ZN(n1244) );
  OAI221_X1 U826 ( .B1(n479), .B2(n36), .C1(n447), .C2(n33), .A(n1252), .ZN(
        n1249) );
  AOI22_X1 U827 ( .A1(n30), .A2(\REGISTERS[7][28] ), .B1(n25), .B2(
        \REGISTERS[6][28] ), .ZN(n1252) );
  OAI221_X1 U828 ( .B1(n1992), .B2(n81), .C1(n1960), .C2(n78), .A(n1226), .ZN(
        n1223) );
  AOI22_X1 U829 ( .A1(n75), .A2(\REGISTERS[23][29] ), .B1(n70), .B2(
        \REGISTERS[22][29] ), .ZN(n1226) );
  OAI221_X1 U830 ( .B1(n478), .B2(n36), .C1(n446), .C2(n33), .A(n1234), .ZN(
        n1231) );
  AOI22_X1 U831 ( .A1(n30), .A2(\REGISTERS[7][29] ), .B1(n25), .B2(
        \REGISTERS[6][29] ), .ZN(n1234) );
  OAI221_X1 U832 ( .B1(n1991), .B2(n81), .C1(n1959), .C2(n78), .A(n1208), .ZN(
        n1205) );
  AOI22_X1 U833 ( .A1(n75), .A2(\REGISTERS[23][30] ), .B1(n70), .B2(
        \REGISTERS[22][30] ), .ZN(n1208) );
  OAI221_X1 U834 ( .B1(n477), .B2(n36), .C1(n445), .C2(n33), .A(n1216), .ZN(
        n1213) );
  AOI22_X1 U835 ( .A1(n30), .A2(\REGISTERS[7][30] ), .B1(n25), .B2(
        \REGISTERS[6][30] ), .ZN(n1216) );
  OAI221_X1 U836 ( .B1(n1990), .B2(n81), .C1(n1958), .C2(n78), .A(n1164), .ZN(
        n1155) );
  AOI22_X1 U837 ( .A1(n75), .A2(\REGISTERS[23][31] ), .B1(n70), .B2(
        \REGISTERS[22][31] ), .ZN(n1164) );
  OAI221_X1 U838 ( .B1(n476), .B2(n36), .C1(n444), .C2(n33), .A(n1188), .ZN(
        n1179) );
  AOI22_X1 U839 ( .A1(n30), .A2(\REGISTERS[7][31] ), .B1(n25), .B2(
        \REGISTERS[6][31] ), .ZN(n1188) );
  OAI221_X1 U840 ( .B1(n499), .B2(n34), .C1(n467), .C2(n31), .A(n1612), .ZN(
        n1609) );
  AOI22_X1 U841 ( .A1(n28), .A2(\REGISTERS[7][8] ), .B1(n26), .B2(
        \REGISTERS[6][8] ), .ZN(n1612) );
  OAI221_X1 U842 ( .B1(n498), .B2(n34), .C1(n466), .C2(n31), .A(n1594), .ZN(
        n1591) );
  AOI22_X1 U843 ( .A1(n28), .A2(\REGISTERS[7][9] ), .B1(n26), .B2(
        \REGISTERS[6][9] ), .ZN(n1594) );
  OAI221_X1 U844 ( .B1(n497), .B2(n34), .C1(n465), .C2(n31), .A(n1576), .ZN(
        n1573) );
  AOI22_X1 U845 ( .A1(n28), .A2(\REGISTERS[7][10] ), .B1(n26), .B2(
        \REGISTERS[6][10] ), .ZN(n1576) );
  OAI221_X1 U846 ( .B1(n496), .B2(n34), .C1(n464), .C2(n31), .A(n1558), .ZN(
        n1555) );
  AOI22_X1 U847 ( .A1(n28), .A2(\REGISTERS[7][11] ), .B1(n26), .B2(
        \REGISTERS[6][11] ), .ZN(n1558) );
  OAI221_X1 U848 ( .B1(n495), .B2(n35), .C1(n463), .C2(n32), .A(n1540), .ZN(
        n1537) );
  AOI22_X1 U849 ( .A1(n29), .A2(\REGISTERS[7][12] ), .B1(n26), .B2(
        \REGISTERS[6][12] ), .ZN(n1540) );
  OAI221_X1 U850 ( .B1(n494), .B2(n35), .C1(n462), .C2(n32), .A(n1522), .ZN(
        n1519) );
  AOI22_X1 U851 ( .A1(n29), .A2(\REGISTERS[7][13] ), .B1(n26), .B2(
        \REGISTERS[6][13] ), .ZN(n1522) );
  OAI221_X1 U852 ( .B1(n493), .B2(n35), .C1(n461), .C2(n32), .A(n1504), .ZN(
        n1501) );
  AOI22_X1 U853 ( .A1(n29), .A2(\REGISTERS[7][14] ), .B1(n26), .B2(
        \REGISTERS[6][14] ), .ZN(n1504) );
  OAI221_X1 U854 ( .B1(n492), .B2(n35), .C1(n460), .C2(n32), .A(n1486), .ZN(
        n1483) );
  AOI22_X1 U855 ( .A1(n29), .A2(\REGISTERS[7][15] ), .B1(n26), .B2(
        \REGISTERS[6][15] ), .ZN(n1486) );
  OAI221_X1 U856 ( .B1(n491), .B2(n35), .C1(n459), .C2(n32), .A(n1468), .ZN(
        n1465) );
  AOI22_X1 U857 ( .A1(n29), .A2(\REGISTERS[7][16] ), .B1(n26), .B2(
        \REGISTERS[6][16] ), .ZN(n1468) );
  OAI221_X1 U858 ( .B1(n490), .B2(n35), .C1(n458), .C2(n32), .A(n1450), .ZN(
        n1447) );
  AOI22_X1 U859 ( .A1(n29), .A2(\REGISTERS[7][17] ), .B1(n26), .B2(
        \REGISTERS[6][17] ), .ZN(n1450) );
  OAI221_X1 U860 ( .B1(n489), .B2(n35), .C1(n457), .C2(n32), .A(n1432), .ZN(
        n1429) );
  AOI22_X1 U861 ( .A1(n29), .A2(\REGISTERS[7][18] ), .B1(n26), .B2(
        \REGISTERS[6][18] ), .ZN(n1432) );
  OAI221_X1 U862 ( .B1(n488), .B2(n35), .C1(n456), .C2(n32), .A(n1414), .ZN(
        n1411) );
  AOI22_X1 U863 ( .A1(n29), .A2(\REGISTERS[7][19] ), .B1(n26), .B2(
        \REGISTERS[6][19] ), .ZN(n1414) );
  OAI221_X1 U864 ( .B1(n487), .B2(n35), .C1(n455), .C2(n32), .A(n1396), .ZN(
        n1393) );
  AOI22_X1 U865 ( .A1(n29), .A2(\REGISTERS[7][20] ), .B1(n25), .B2(
        \REGISTERS[6][20] ), .ZN(n1396) );
  OAI221_X1 U866 ( .B1(n486), .B2(n35), .C1(n454), .C2(n32), .A(n1378), .ZN(
        n1375) );
  AOI22_X1 U867 ( .A1(n29), .A2(\REGISTERS[7][21] ), .B1(n25), .B2(
        \REGISTERS[6][21] ), .ZN(n1378) );
  OAI221_X1 U868 ( .B1(n485), .B2(n35), .C1(n453), .C2(n32), .A(n1360), .ZN(
        n1357) );
  AOI22_X1 U869 ( .A1(n29), .A2(\REGISTERS[7][22] ), .B1(n25), .B2(
        \REGISTERS[6][22] ), .ZN(n1360) );
  OAI221_X1 U870 ( .B1(n484), .B2(n35), .C1(n452), .C2(n32), .A(n1342), .ZN(
        n1339) );
  AOI22_X1 U871 ( .A1(n29), .A2(\REGISTERS[7][23] ), .B1(n25), .B2(
        \REGISTERS[6][23] ), .ZN(n1342) );
  OAI221_X1 U872 ( .B1(n186), .B2(n1933), .C1(n183), .C2(n1901), .A(n691), 
        .ZN(n690) );
  AOI22_X1 U873 ( .A1(\REGISTERS[19][24] ), .A2(n180), .B1(\REGISTERS[18][24] ), .B2(n177), .ZN(n691) );
  OAI221_X1 U874 ( .B1(n174), .B2(n1997), .C1(n171), .C2(n1965), .A(n692), 
        .ZN(n689) );
  AOI22_X1 U875 ( .A1(\REGISTERS[23][24] ), .A2(n168), .B1(\REGISTERS[22][24] ), .B2(n165), .ZN(n692) );
  OAI221_X1 U876 ( .B1(n162), .B2(n2061), .C1(n159), .C2(n2029), .A(n693), 
        .ZN(n688) );
  AOI22_X1 U877 ( .A1(\REGISTERS[27][24] ), .A2(n156), .B1(\REGISTERS[26][24] ), .B2(n153), .ZN(n693) );
  OAI221_X1 U878 ( .B1(n150), .B2(n2125), .C1(n147), .C2(n2093), .A(n694), 
        .ZN(n687) );
  AOI22_X1 U879 ( .A1(\REGISTERS[29][24] ), .A2(n144), .B1(\REGISTERS[28][24] ), .B2(n141), .ZN(n694) );
  OAI221_X1 U880 ( .B1(n117), .B2(n1805), .C1(n114), .C2(n515), .A(n701), .ZN(
        n696) );
  AOI22_X1 U881 ( .A1(\REGISTERS[11][24] ), .A2(n111), .B1(\REGISTERS[10][24] ), .B2(n108), .ZN(n701) );
  OAI221_X1 U882 ( .B1(n129), .B2(n483), .C1(n126), .C2(n451), .A(n700), .ZN(
        n697) );
  AOI22_X1 U883 ( .A1(\REGISTERS[7][24] ), .A2(n123), .B1(\REGISTERS[6][24] ), 
        .B2(n120), .ZN(n700) );
  OAI221_X1 U884 ( .B1(n105), .B2(n1869), .C1(n102), .C2(n1837), .A(n702), 
        .ZN(n695) );
  AOI22_X1 U885 ( .A1(\REGISTERS[15][24] ), .A2(n99), .B1(\REGISTERS[14][24] ), 
        .B2(n96), .ZN(n702) );
  OAI221_X1 U886 ( .B1(n186), .B2(n1932), .C1(n183), .C2(n1900), .A(n673), 
        .ZN(n672) );
  AOI22_X1 U887 ( .A1(\REGISTERS[19][25] ), .A2(n180), .B1(\REGISTERS[18][25] ), .B2(n177), .ZN(n673) );
  OAI221_X1 U888 ( .B1(n174), .B2(n1996), .C1(n171), .C2(n1964), .A(n674), 
        .ZN(n671) );
  AOI22_X1 U889 ( .A1(\REGISTERS[23][25] ), .A2(n168), .B1(\REGISTERS[22][25] ), .B2(n165), .ZN(n674) );
  OAI221_X1 U890 ( .B1(n162), .B2(n2060), .C1(n159), .C2(n2028), .A(n675), 
        .ZN(n670) );
  AOI22_X1 U891 ( .A1(\REGISTERS[27][25] ), .A2(n156), .B1(\REGISTERS[26][25] ), .B2(n153), .ZN(n675) );
  OAI221_X1 U892 ( .B1(n150), .B2(n2124), .C1(n147), .C2(n2092), .A(n676), 
        .ZN(n669) );
  AOI22_X1 U893 ( .A1(\REGISTERS[29][25] ), .A2(n144), .B1(\REGISTERS[28][25] ), .B2(n141), .ZN(n676) );
  OAI221_X1 U894 ( .B1(n117), .B2(n1804), .C1(n114), .C2(n514), .A(n683), .ZN(
        n678) );
  AOI22_X1 U895 ( .A1(\REGISTERS[11][25] ), .A2(n111), .B1(\REGISTERS[10][25] ), .B2(n108), .ZN(n683) );
  OAI221_X1 U896 ( .B1(n129), .B2(n482), .C1(n126), .C2(n450), .A(n682), .ZN(
        n679) );
  AOI22_X1 U897 ( .A1(\REGISTERS[7][25] ), .A2(n123), .B1(\REGISTERS[6][25] ), 
        .B2(n120), .ZN(n682) );
  OAI221_X1 U898 ( .B1(n105), .B2(n1868), .C1(n102), .C2(n1836), .A(n684), 
        .ZN(n677) );
  AOI22_X1 U899 ( .A1(\REGISTERS[15][25] ), .A2(n99), .B1(\REGISTERS[14][25] ), 
        .B2(n96), .ZN(n684) );
  OAI221_X1 U900 ( .B1(n186), .B2(n1931), .C1(n183), .C2(n1899), .A(n655), 
        .ZN(n654) );
  AOI22_X1 U901 ( .A1(\REGISTERS[19][26] ), .A2(n180), .B1(\REGISTERS[18][26] ), .B2(n177), .ZN(n655) );
  OAI221_X1 U902 ( .B1(n174), .B2(n1995), .C1(n171), .C2(n1963), .A(n656), 
        .ZN(n653) );
  AOI22_X1 U903 ( .A1(\REGISTERS[23][26] ), .A2(n168), .B1(\REGISTERS[22][26] ), .B2(n165), .ZN(n656) );
  OAI221_X1 U904 ( .B1(n162), .B2(n2059), .C1(n159), .C2(n2027), .A(n657), 
        .ZN(n652) );
  AOI22_X1 U905 ( .A1(\REGISTERS[27][26] ), .A2(n156), .B1(\REGISTERS[26][26] ), .B2(n153), .ZN(n657) );
  OAI221_X1 U906 ( .B1(n150), .B2(n2123), .C1(n147), .C2(n2091), .A(n658), 
        .ZN(n651) );
  AOI22_X1 U907 ( .A1(\REGISTERS[29][26] ), .A2(n144), .B1(\REGISTERS[28][26] ), .B2(n141), .ZN(n658) );
  OAI221_X1 U908 ( .B1(n117), .B2(n1803), .C1(n114), .C2(n513), .A(n665), .ZN(
        n660) );
  AOI22_X1 U909 ( .A1(\REGISTERS[11][26] ), .A2(n111), .B1(\REGISTERS[10][26] ), .B2(n108), .ZN(n665) );
  OAI221_X1 U910 ( .B1(n129), .B2(n481), .C1(n126), .C2(n449), .A(n664), .ZN(
        n661) );
  AOI22_X1 U911 ( .A1(\REGISTERS[7][26] ), .A2(n123), .B1(\REGISTERS[6][26] ), 
        .B2(n120), .ZN(n664) );
  OAI221_X1 U912 ( .B1(n105), .B2(n1867), .C1(n102), .C2(n1835), .A(n666), 
        .ZN(n659) );
  AOI22_X1 U913 ( .A1(\REGISTERS[15][26] ), .A2(n99), .B1(\REGISTERS[14][26] ), 
        .B2(n96), .ZN(n666) );
  OAI221_X1 U914 ( .B1(n186), .B2(n1930), .C1(n183), .C2(n1898), .A(n637), 
        .ZN(n636) );
  AOI22_X1 U915 ( .A1(\REGISTERS[19][27] ), .A2(n180), .B1(\REGISTERS[18][27] ), .B2(n177), .ZN(n637) );
  OAI221_X1 U916 ( .B1(n174), .B2(n1994), .C1(n171), .C2(n1962), .A(n638), 
        .ZN(n635) );
  AOI22_X1 U917 ( .A1(\REGISTERS[23][27] ), .A2(n168), .B1(\REGISTERS[22][27] ), .B2(n165), .ZN(n638) );
  OAI221_X1 U918 ( .B1(n162), .B2(n2058), .C1(n159), .C2(n2026), .A(n639), 
        .ZN(n634) );
  AOI22_X1 U919 ( .A1(\REGISTERS[27][27] ), .A2(n156), .B1(\REGISTERS[26][27] ), .B2(n153), .ZN(n639) );
  OAI221_X1 U920 ( .B1(n150), .B2(n2122), .C1(n147), .C2(n2090), .A(n640), 
        .ZN(n633) );
  AOI22_X1 U921 ( .A1(\REGISTERS[29][27] ), .A2(n144), .B1(\REGISTERS[28][27] ), .B2(n141), .ZN(n640) );
  OAI221_X1 U922 ( .B1(n117), .B2(n1802), .C1(n114), .C2(n512), .A(n647), .ZN(
        n642) );
  AOI22_X1 U923 ( .A1(\REGISTERS[11][27] ), .A2(n111), .B1(\REGISTERS[10][27] ), .B2(n108), .ZN(n647) );
  OAI221_X1 U924 ( .B1(n129), .B2(n480), .C1(n126), .C2(n448), .A(n646), .ZN(
        n643) );
  AOI22_X1 U925 ( .A1(\REGISTERS[7][27] ), .A2(n123), .B1(\REGISTERS[6][27] ), 
        .B2(n120), .ZN(n646) );
  OAI221_X1 U926 ( .B1(n105), .B2(n1866), .C1(n102), .C2(n1834), .A(n648), 
        .ZN(n641) );
  AOI22_X1 U927 ( .A1(\REGISTERS[15][27] ), .A2(n99), .B1(\REGISTERS[14][27] ), 
        .B2(n96), .ZN(n648) );
  OAI221_X1 U928 ( .B1(n186), .B2(n1929), .C1(n183), .C2(n1897), .A(n619), 
        .ZN(n618) );
  AOI22_X1 U929 ( .A1(\REGISTERS[19][28] ), .A2(n180), .B1(\REGISTERS[18][28] ), .B2(n177), .ZN(n619) );
  OAI221_X1 U930 ( .B1(n174), .B2(n1993), .C1(n171), .C2(n1961), .A(n620), 
        .ZN(n617) );
  AOI22_X1 U931 ( .A1(\REGISTERS[23][28] ), .A2(n168), .B1(\REGISTERS[22][28] ), .B2(n165), .ZN(n620) );
  OAI221_X1 U932 ( .B1(n162), .B2(n2057), .C1(n159), .C2(n2025), .A(n621), 
        .ZN(n616) );
  AOI22_X1 U933 ( .A1(\REGISTERS[27][28] ), .A2(n156), .B1(\REGISTERS[26][28] ), .B2(n153), .ZN(n621) );
  OAI221_X1 U934 ( .B1(n150), .B2(n2121), .C1(n147), .C2(n2089), .A(n622), 
        .ZN(n615) );
  AOI22_X1 U935 ( .A1(\REGISTERS[29][28] ), .A2(n144), .B1(\REGISTERS[28][28] ), .B2(n141), .ZN(n622) );
  OAI221_X1 U936 ( .B1(n117), .B2(n1801), .C1(n114), .C2(n511), .A(n629), .ZN(
        n624) );
  AOI22_X1 U937 ( .A1(\REGISTERS[11][28] ), .A2(n111), .B1(\REGISTERS[10][28] ), .B2(n108), .ZN(n629) );
  OAI221_X1 U938 ( .B1(n129), .B2(n479), .C1(n126), .C2(n447), .A(n628), .ZN(
        n625) );
  AOI22_X1 U939 ( .A1(\REGISTERS[7][28] ), .A2(n123), .B1(\REGISTERS[6][28] ), 
        .B2(n120), .ZN(n628) );
  OAI221_X1 U940 ( .B1(n105), .B2(n1865), .C1(n102), .C2(n1833), .A(n630), 
        .ZN(n623) );
  AOI22_X1 U941 ( .A1(\REGISTERS[15][28] ), .A2(n99), .B1(\REGISTERS[14][28] ), 
        .B2(n96), .ZN(n630) );
  OAI221_X1 U942 ( .B1(n186), .B2(n1928), .C1(n183), .C2(n1896), .A(n601), 
        .ZN(n600) );
  AOI22_X1 U943 ( .A1(\REGISTERS[19][29] ), .A2(n180), .B1(\REGISTERS[18][29] ), .B2(n177), .ZN(n601) );
  OAI221_X1 U944 ( .B1(n174), .B2(n1992), .C1(n171), .C2(n1960), .A(n602), 
        .ZN(n599) );
  AOI22_X1 U945 ( .A1(\REGISTERS[23][29] ), .A2(n168), .B1(\REGISTERS[22][29] ), .B2(n165), .ZN(n602) );
  OAI221_X1 U946 ( .B1(n162), .B2(n2056), .C1(n159), .C2(n2024), .A(n603), 
        .ZN(n598) );
  AOI22_X1 U947 ( .A1(\REGISTERS[27][29] ), .A2(n156), .B1(\REGISTERS[26][29] ), .B2(n153), .ZN(n603) );
  OAI221_X1 U948 ( .B1(n150), .B2(n2120), .C1(n147), .C2(n2088), .A(n604), 
        .ZN(n597) );
  AOI22_X1 U949 ( .A1(\REGISTERS[29][29] ), .A2(n144), .B1(\REGISTERS[28][29] ), .B2(n141), .ZN(n604) );
  OAI221_X1 U950 ( .B1(n117), .B2(n1800), .C1(n114), .C2(n510), .A(n611), .ZN(
        n606) );
  AOI22_X1 U951 ( .A1(\REGISTERS[11][29] ), .A2(n111), .B1(\REGISTERS[10][29] ), .B2(n108), .ZN(n611) );
  OAI221_X1 U952 ( .B1(n129), .B2(n478), .C1(n126), .C2(n446), .A(n610), .ZN(
        n607) );
  AOI22_X1 U953 ( .A1(\REGISTERS[7][29] ), .A2(n123), .B1(\REGISTERS[6][29] ), 
        .B2(n120), .ZN(n610) );
  OAI221_X1 U954 ( .B1(n105), .B2(n1864), .C1(n102), .C2(n1832), .A(n612), 
        .ZN(n605) );
  AOI22_X1 U955 ( .A1(\REGISTERS[15][29] ), .A2(n99), .B1(\REGISTERS[14][29] ), 
        .B2(n96), .ZN(n612) );
  OAI221_X1 U956 ( .B1(n186), .B2(n1927), .C1(n183), .C2(n1895), .A(n583), 
        .ZN(n582) );
  AOI22_X1 U957 ( .A1(\REGISTERS[19][30] ), .A2(n180), .B1(\REGISTERS[18][30] ), .B2(n177), .ZN(n583) );
  OAI221_X1 U958 ( .B1(n174), .B2(n1991), .C1(n171), .C2(n1959), .A(n584), 
        .ZN(n581) );
  AOI22_X1 U959 ( .A1(\REGISTERS[23][30] ), .A2(n168), .B1(\REGISTERS[22][30] ), .B2(n165), .ZN(n584) );
  OAI221_X1 U960 ( .B1(n162), .B2(n2055), .C1(n159), .C2(n2023), .A(n585), 
        .ZN(n580) );
  AOI22_X1 U961 ( .A1(\REGISTERS[27][30] ), .A2(n156), .B1(\REGISTERS[26][30] ), .B2(n153), .ZN(n585) );
  OAI221_X1 U962 ( .B1(n150), .B2(n2119), .C1(n147), .C2(n2087), .A(n586), 
        .ZN(n579) );
  AOI22_X1 U963 ( .A1(\REGISTERS[29][30] ), .A2(n144), .B1(\REGISTERS[28][30] ), .B2(n141), .ZN(n586) );
  OAI221_X1 U964 ( .B1(n117), .B2(n1799), .C1(n114), .C2(n509), .A(n593), .ZN(
        n588) );
  AOI22_X1 U965 ( .A1(\REGISTERS[11][30] ), .A2(n111), .B1(\REGISTERS[10][30] ), .B2(n108), .ZN(n593) );
  OAI221_X1 U966 ( .B1(n129), .B2(n477), .C1(n126), .C2(n445), .A(n592), .ZN(
        n589) );
  AOI22_X1 U967 ( .A1(\REGISTERS[7][30] ), .A2(n123), .B1(\REGISTERS[6][30] ), 
        .B2(n120), .ZN(n592) );
  OAI221_X1 U968 ( .B1(n105), .B2(n1863), .C1(n102), .C2(n1831), .A(n594), 
        .ZN(n587) );
  AOI22_X1 U969 ( .A1(\REGISTERS[15][30] ), .A2(n99), .B1(\REGISTERS[14][30] ), 
        .B2(n96), .ZN(n594) );
  OAI221_X1 U970 ( .B1(n186), .B2(n1926), .C1(n183), .C2(n1894), .A(n535), 
        .ZN(n532) );
  AOI22_X1 U971 ( .A1(\REGISTERS[19][31] ), .A2(n180), .B1(\REGISTERS[18][31] ), .B2(n177), .ZN(n535) );
  OAI221_X1 U972 ( .B1(n174), .B2(n1990), .C1(n171), .C2(n1958), .A(n540), 
        .ZN(n531) );
  AOI22_X1 U973 ( .A1(\REGISTERS[23][31] ), .A2(n168), .B1(\REGISTERS[22][31] ), .B2(n165), .ZN(n540) );
  OAI221_X1 U974 ( .B1(n162), .B2(n2054), .C1(n159), .C2(n2022), .A(n545), 
        .ZN(n530) );
  AOI22_X1 U975 ( .A1(\REGISTERS[27][31] ), .A2(n156), .B1(\REGISTERS[26][31] ), .B2(n153), .ZN(n545) );
  OAI221_X1 U976 ( .B1(n150), .B2(n2118), .C1(n147), .C2(n2086), .A(n550), 
        .ZN(n529) );
  AOI22_X1 U977 ( .A1(\REGISTERS[29][31] ), .A2(n144), .B1(\REGISTERS[28][31] ), .B2(n141), .ZN(n550) );
  OAI221_X1 U978 ( .B1(n117), .B2(n1798), .C1(n114), .C2(n508), .A(n569), .ZN(
        n554) );
  AOI22_X1 U979 ( .A1(\REGISTERS[11][31] ), .A2(n111), .B1(\REGISTERS[10][31] ), .B2(n108), .ZN(n569) );
  OAI221_X1 U980 ( .B1(n129), .B2(n476), .C1(n126), .C2(n444), .A(n564), .ZN(
        n555) );
  AOI22_X1 U981 ( .A1(\REGISTERS[7][31] ), .A2(n123), .B1(\REGISTERS[6][31] ), 
        .B2(n120), .ZN(n564) );
  OAI221_X1 U982 ( .B1(n105), .B2(n1862), .C1(n102), .C2(n1830), .A(n574), 
        .ZN(n553) );
  AOI22_X1 U983 ( .A1(\REGISTERS[15][31] ), .A2(n99), .B1(\REGISTERS[14][31] ), 
        .B2(n96), .ZN(n574) );
  AOI22_X1 U984 ( .A1(n4), .A2(\REGISTERS[15][0] ), .B1(n3), .B2(
        \REGISTERS[14][0] ), .ZN(n1773) );
  AOI22_X1 U985 ( .A1(n4), .A2(\REGISTERS[15][1] ), .B1(n3), .B2(
        \REGISTERS[14][1] ), .ZN(n1740) );
  AOI22_X1 U986 ( .A1(n4), .A2(\REGISTERS[15][2] ), .B1(n3), .B2(
        \REGISTERS[14][2] ), .ZN(n1722) );
  AOI22_X1 U987 ( .A1(n4), .A2(\REGISTERS[15][3] ), .B1(n3), .B2(
        \REGISTERS[14][3] ), .ZN(n1704) );
  AOI22_X1 U988 ( .A1(n4), .A2(\REGISTERS[15][4] ), .B1(n3), .B2(
        \REGISTERS[14][4] ), .ZN(n1686) );
  AOI22_X1 U989 ( .A1(n4), .A2(\REGISTERS[15][5] ), .B1(n3), .B2(
        \REGISTERS[14][5] ), .ZN(n1668) );
  AOI22_X1 U990 ( .A1(n4), .A2(\REGISTERS[15][6] ), .B1(n3), .B2(
        \REGISTERS[14][6] ), .ZN(n1650) );
  AOI22_X1 U991 ( .A1(n4), .A2(\REGISTERS[15][7] ), .B1(n3), .B2(
        \REGISTERS[14][7] ), .ZN(n1632) );
  AOI22_X1 U992 ( .A1(n4), .A2(\REGISTERS[15][8] ), .B1(n2), .B2(
        \REGISTERS[14][8] ), .ZN(n1614) );
  AOI22_X1 U993 ( .A1(n4), .A2(\REGISTERS[15][9] ), .B1(n2), .B2(
        \REGISTERS[14][9] ), .ZN(n1596) );
  AOI22_X1 U994 ( .A1(n4), .A2(\REGISTERS[15][10] ), .B1(n2), .B2(
        \REGISTERS[14][10] ), .ZN(n1578) );
  AOI22_X1 U995 ( .A1(n4), .A2(\REGISTERS[15][11] ), .B1(n2), .B2(
        \REGISTERS[14][11] ), .ZN(n1560) );
  AOI22_X1 U996 ( .A1(n5), .A2(\REGISTERS[15][12] ), .B1(n2), .B2(
        \REGISTERS[14][12] ), .ZN(n1542) );
  AOI22_X1 U997 ( .A1(n5), .A2(\REGISTERS[15][13] ), .B1(n2), .B2(
        \REGISTERS[14][13] ), .ZN(n1524) );
  AOI22_X1 U998 ( .A1(n5), .A2(\REGISTERS[15][14] ), .B1(n2), .B2(
        \REGISTERS[14][14] ), .ZN(n1506) );
  AOI22_X1 U999 ( .A1(n5), .A2(\REGISTERS[15][15] ), .B1(n2), .B2(
        \REGISTERS[14][15] ), .ZN(n1488) );
  AOI22_X1 U1000 ( .A1(n5), .A2(\REGISTERS[15][16] ), .B1(n2), .B2(
        \REGISTERS[14][16] ), .ZN(n1470) );
  AOI22_X1 U1001 ( .A1(n5), .A2(\REGISTERS[15][17] ), .B1(n2), .B2(
        \REGISTERS[14][17] ), .ZN(n1452) );
  AOI22_X1 U1002 ( .A1(n5), .A2(\REGISTERS[15][18] ), .B1(n2), .B2(
        \REGISTERS[14][18] ), .ZN(n1434) );
  AOI22_X1 U1003 ( .A1(n5), .A2(\REGISTERS[15][19] ), .B1(n2), .B2(
        \REGISTERS[14][19] ), .ZN(n1416) );
  AOI22_X1 U1004 ( .A1(n5), .A2(\REGISTERS[15][20] ), .B1(n1), .B2(
        \REGISTERS[14][20] ), .ZN(n1398) );
  AOI22_X1 U1005 ( .A1(n5), .A2(\REGISTERS[15][21] ), .B1(n1), .B2(
        \REGISTERS[14][21] ), .ZN(n1380) );
  AOI22_X1 U1006 ( .A1(n5), .A2(\REGISTERS[15][22] ), .B1(n1), .B2(
        \REGISTERS[14][22] ), .ZN(n1362) );
  AOI22_X1 U1007 ( .A1(n5), .A2(\REGISTERS[15][23] ), .B1(n1), .B2(
        \REGISTERS[14][23] ), .ZN(n1344) );
  AOI22_X1 U1008 ( .A1(n6), .A2(\REGISTERS[15][24] ), .B1(n1), .B2(
        \REGISTERS[14][24] ), .ZN(n1326) );
  AOI22_X1 U1009 ( .A1(n6), .A2(\REGISTERS[15][25] ), .B1(n1), .B2(
        \REGISTERS[14][25] ), .ZN(n1308) );
  AOI22_X1 U1010 ( .A1(n6), .A2(\REGISTERS[15][26] ), .B1(n1), .B2(
        \REGISTERS[14][26] ), .ZN(n1290) );
  AOI22_X1 U1011 ( .A1(n6), .A2(\REGISTERS[15][27] ), .B1(n1), .B2(
        \REGISTERS[14][27] ), .ZN(n1272) );
  AOI22_X1 U1012 ( .A1(n6), .A2(\REGISTERS[15][28] ), .B1(n1), .B2(
        \REGISTERS[14][28] ), .ZN(n1254) );
  AOI22_X1 U1013 ( .A1(n6), .A2(\REGISTERS[15][29] ), .B1(n1), .B2(
        \REGISTERS[14][29] ), .ZN(n1236) );
  AOI22_X1 U1014 ( .A1(n6), .A2(\REGISTERS[15][30] ), .B1(n1), .B2(
        \REGISTERS[14][30] ), .ZN(n1218) );
  AOI22_X1 U1015 ( .A1(n6), .A2(\REGISTERS[15][31] ), .B1(n1), .B2(
        \REGISTERS[14][31] ), .ZN(n1198) );
  OAI221_X1 U1016 ( .B1(n184), .B2(n1957), .C1(n181), .C2(n1925), .A(n1123), 
        .ZN(n1122) );
  AOI22_X1 U1017 ( .A1(\REGISTERS[19][0] ), .A2(n178), .B1(\REGISTERS[18][0] ), 
        .B2(n175), .ZN(n1123) );
  OAI221_X1 U1018 ( .B1(n172), .B2(n2021), .C1(n169), .C2(n1989), .A(n1128), 
        .ZN(n1121) );
  AOI22_X1 U1019 ( .A1(\REGISTERS[23][0] ), .A2(n166), .B1(\REGISTERS[22][0] ), 
        .B2(n163), .ZN(n1128) );
  OAI221_X1 U1020 ( .B1(n160), .B2(n2085), .C1(n157), .C2(n2053), .A(n1132), 
        .ZN(n1120) );
  AOI22_X1 U1021 ( .A1(\REGISTERS[27][0] ), .A2(n154), .B1(\REGISTERS[26][0] ), 
        .B2(n151), .ZN(n1132) );
  OAI221_X1 U1022 ( .B1(n148), .B2(n2149), .C1(n145), .C2(n2117), .A(n1135), 
        .ZN(n1119) );
  AOI22_X1 U1023 ( .A1(\REGISTERS[29][0] ), .A2(n142), .B1(\REGISTERS[28][0] ), 
        .B2(n139), .ZN(n1135) );
  OAI221_X1 U1024 ( .B1(n115), .B2(n1829), .C1(n112), .C2(n1797), .A(n1146), 
        .ZN(n1138) );
  AOI22_X1 U1025 ( .A1(\REGISTERS[11][0] ), .A2(n109), .B1(\REGISTERS[10][0] ), 
        .B2(n106), .ZN(n1146) );
  OAI221_X1 U1026 ( .B1(n127), .B2(n507), .C1(n124), .C2(n475), .A(n1144), 
        .ZN(n1139) );
  AOI22_X1 U1027 ( .A1(\REGISTERS[7][0] ), .A2(n121), .B1(\REGISTERS[6][0] ), 
        .B2(n118), .ZN(n1144) );
  OAI221_X1 U1028 ( .B1(n103), .B2(n1893), .C1(n100), .C2(n1861), .A(n1149), 
        .ZN(n1137) );
  AOI22_X1 U1029 ( .A1(\REGISTERS[15][0] ), .A2(n97), .B1(\REGISTERS[14][0] ), 
        .B2(n94), .ZN(n1149) );
  OAI221_X1 U1030 ( .B1(n184), .B2(n1956), .C1(n181), .C2(n1924), .A(n1105), 
        .ZN(n1104) );
  AOI22_X1 U1031 ( .A1(\REGISTERS[19][1] ), .A2(n178), .B1(\REGISTERS[18][1] ), 
        .B2(n175), .ZN(n1105) );
  OAI221_X1 U1032 ( .B1(n172), .B2(n2020), .C1(n169), .C2(n1988), .A(n1106), 
        .ZN(n1103) );
  AOI22_X1 U1033 ( .A1(\REGISTERS[23][1] ), .A2(n166), .B1(\REGISTERS[22][1] ), 
        .B2(n163), .ZN(n1106) );
  OAI221_X1 U1034 ( .B1(n160), .B2(n2084), .C1(n157), .C2(n2052), .A(n1107), 
        .ZN(n1102) );
  AOI22_X1 U1035 ( .A1(\REGISTERS[27][1] ), .A2(n154), .B1(\REGISTERS[26][1] ), 
        .B2(n151), .ZN(n1107) );
  OAI221_X1 U1036 ( .B1(n148), .B2(n2148), .C1(n145), .C2(n2116), .A(n1108), 
        .ZN(n1101) );
  AOI22_X1 U1037 ( .A1(\REGISTERS[29][1] ), .A2(n142), .B1(\REGISTERS[28][1] ), 
        .B2(n139), .ZN(n1108) );
  OAI221_X1 U1038 ( .B1(n115), .B2(n1828), .C1(n112), .C2(n1796), .A(n1115), 
        .ZN(n1110) );
  AOI22_X1 U1039 ( .A1(\REGISTERS[11][1] ), .A2(n109), .B1(\REGISTERS[10][1] ), 
        .B2(n106), .ZN(n1115) );
  OAI221_X1 U1040 ( .B1(n127), .B2(n506), .C1(n124), .C2(n474), .A(n1114), 
        .ZN(n1111) );
  AOI22_X1 U1041 ( .A1(\REGISTERS[7][1] ), .A2(n121), .B1(\REGISTERS[6][1] ), 
        .B2(n118), .ZN(n1114) );
  OAI221_X1 U1042 ( .B1(n103), .B2(n1892), .C1(n100), .C2(n1860), .A(n1116), 
        .ZN(n1109) );
  AOI22_X1 U1043 ( .A1(\REGISTERS[15][1] ), .A2(n97), .B1(\REGISTERS[14][1] ), 
        .B2(n94), .ZN(n1116) );
  OAI221_X1 U1044 ( .B1(n184), .B2(n1955), .C1(n181), .C2(n1923), .A(n1087), 
        .ZN(n1086) );
  AOI22_X1 U1045 ( .A1(\REGISTERS[19][2] ), .A2(n178), .B1(\REGISTERS[18][2] ), 
        .B2(n175), .ZN(n1087) );
  OAI221_X1 U1046 ( .B1(n172), .B2(n2019), .C1(n169), .C2(n1987), .A(n1088), 
        .ZN(n1085) );
  AOI22_X1 U1047 ( .A1(\REGISTERS[23][2] ), .A2(n166), .B1(\REGISTERS[22][2] ), 
        .B2(n163), .ZN(n1088) );
  OAI221_X1 U1048 ( .B1(n160), .B2(n2083), .C1(n157), .C2(n2051), .A(n1089), 
        .ZN(n1084) );
  AOI22_X1 U1049 ( .A1(\REGISTERS[27][2] ), .A2(n154), .B1(\REGISTERS[26][2] ), 
        .B2(n151), .ZN(n1089) );
  OAI221_X1 U1050 ( .B1(n148), .B2(n2147), .C1(n145), .C2(n2115), .A(n1090), 
        .ZN(n1083) );
  AOI22_X1 U1051 ( .A1(\REGISTERS[29][2] ), .A2(n142), .B1(\REGISTERS[28][2] ), 
        .B2(n139), .ZN(n1090) );
  OAI221_X1 U1052 ( .B1(n115), .B2(n1827), .C1(n112), .C2(n1795), .A(n1097), 
        .ZN(n1092) );
  AOI22_X1 U1053 ( .A1(\REGISTERS[11][2] ), .A2(n109), .B1(\REGISTERS[10][2] ), 
        .B2(n106), .ZN(n1097) );
  OAI221_X1 U1054 ( .B1(n127), .B2(n505), .C1(n124), .C2(n473), .A(n1096), 
        .ZN(n1093) );
  AOI22_X1 U1055 ( .A1(\REGISTERS[7][2] ), .A2(n121), .B1(\REGISTERS[6][2] ), 
        .B2(n118), .ZN(n1096) );
  OAI221_X1 U1056 ( .B1(n103), .B2(n1891), .C1(n100), .C2(n1859), .A(n1098), 
        .ZN(n1091) );
  AOI22_X1 U1057 ( .A1(\REGISTERS[15][2] ), .A2(n97), .B1(\REGISTERS[14][2] ), 
        .B2(n94), .ZN(n1098) );
  OAI221_X1 U1058 ( .B1(n184), .B2(n1954), .C1(n181), .C2(n1922), .A(n1069), 
        .ZN(n1068) );
  AOI22_X1 U1059 ( .A1(\REGISTERS[19][3] ), .A2(n178), .B1(\REGISTERS[18][3] ), 
        .B2(n175), .ZN(n1069) );
  OAI221_X1 U1060 ( .B1(n172), .B2(n2018), .C1(n169), .C2(n1986), .A(n1070), 
        .ZN(n1067) );
  AOI22_X1 U1061 ( .A1(\REGISTERS[23][3] ), .A2(n166), .B1(\REGISTERS[22][3] ), 
        .B2(n163), .ZN(n1070) );
  OAI221_X1 U1062 ( .B1(n160), .B2(n2082), .C1(n157), .C2(n2050), .A(n1071), 
        .ZN(n1066) );
  AOI22_X1 U1063 ( .A1(\REGISTERS[27][3] ), .A2(n154), .B1(\REGISTERS[26][3] ), 
        .B2(n151), .ZN(n1071) );
  OAI221_X1 U1064 ( .B1(n148), .B2(n2146), .C1(n145), .C2(n2114), .A(n1072), 
        .ZN(n1065) );
  AOI22_X1 U1065 ( .A1(\REGISTERS[29][3] ), .A2(n142), .B1(\REGISTERS[28][3] ), 
        .B2(n139), .ZN(n1072) );
  OAI221_X1 U1066 ( .B1(n115), .B2(n1826), .C1(n112), .C2(n1794), .A(n1079), 
        .ZN(n1074) );
  AOI22_X1 U1067 ( .A1(\REGISTERS[11][3] ), .A2(n109), .B1(\REGISTERS[10][3] ), 
        .B2(n106), .ZN(n1079) );
  OAI221_X1 U1068 ( .B1(n127), .B2(n504), .C1(n124), .C2(n472), .A(n1078), 
        .ZN(n1075) );
  AOI22_X1 U1069 ( .A1(\REGISTERS[7][3] ), .A2(n121), .B1(\REGISTERS[6][3] ), 
        .B2(n118), .ZN(n1078) );
  OAI221_X1 U1070 ( .B1(n103), .B2(n1890), .C1(n100), .C2(n1858), .A(n1080), 
        .ZN(n1073) );
  AOI22_X1 U1071 ( .A1(\REGISTERS[15][3] ), .A2(n97), .B1(\REGISTERS[14][3] ), 
        .B2(n94), .ZN(n1080) );
  OAI221_X1 U1072 ( .B1(n184), .B2(n1953), .C1(n181), .C2(n1921), .A(n1051), 
        .ZN(n1050) );
  AOI22_X1 U1073 ( .A1(\REGISTERS[19][4] ), .A2(n178), .B1(\REGISTERS[18][4] ), 
        .B2(n175), .ZN(n1051) );
  OAI221_X1 U1074 ( .B1(n172), .B2(n2017), .C1(n169), .C2(n1985), .A(n1052), 
        .ZN(n1049) );
  AOI22_X1 U1075 ( .A1(\REGISTERS[23][4] ), .A2(n166), .B1(\REGISTERS[22][4] ), 
        .B2(n163), .ZN(n1052) );
  OAI221_X1 U1076 ( .B1(n160), .B2(n2081), .C1(n157), .C2(n2049), .A(n1053), 
        .ZN(n1048) );
  AOI22_X1 U1077 ( .A1(\REGISTERS[27][4] ), .A2(n154), .B1(\REGISTERS[26][4] ), 
        .B2(n151), .ZN(n1053) );
  OAI221_X1 U1078 ( .B1(n148), .B2(n2145), .C1(n145), .C2(n2113), .A(n1054), 
        .ZN(n1047) );
  AOI22_X1 U1079 ( .A1(\REGISTERS[29][4] ), .A2(n142), .B1(\REGISTERS[28][4] ), 
        .B2(n139), .ZN(n1054) );
  OAI221_X1 U1080 ( .B1(n115), .B2(n1825), .C1(n112), .C2(n1793), .A(n1061), 
        .ZN(n1056) );
  AOI22_X1 U1081 ( .A1(\REGISTERS[11][4] ), .A2(n109), .B1(\REGISTERS[10][4] ), 
        .B2(n106), .ZN(n1061) );
  OAI221_X1 U1082 ( .B1(n127), .B2(n503), .C1(n124), .C2(n471), .A(n1060), 
        .ZN(n1057) );
  AOI22_X1 U1083 ( .A1(\REGISTERS[7][4] ), .A2(n121), .B1(\REGISTERS[6][4] ), 
        .B2(n118), .ZN(n1060) );
  OAI221_X1 U1084 ( .B1(n103), .B2(n1889), .C1(n100), .C2(n1857), .A(n1062), 
        .ZN(n1055) );
  AOI22_X1 U1085 ( .A1(\REGISTERS[15][4] ), .A2(n97), .B1(\REGISTERS[14][4] ), 
        .B2(n94), .ZN(n1062) );
  OAI221_X1 U1086 ( .B1(n184), .B2(n1952), .C1(n181), .C2(n1920), .A(n1033), 
        .ZN(n1032) );
  AOI22_X1 U1087 ( .A1(\REGISTERS[19][5] ), .A2(n178), .B1(\REGISTERS[18][5] ), 
        .B2(n175), .ZN(n1033) );
  OAI221_X1 U1088 ( .B1(n172), .B2(n2016), .C1(n169), .C2(n1984), .A(n1034), 
        .ZN(n1031) );
  AOI22_X1 U1089 ( .A1(\REGISTERS[23][5] ), .A2(n166), .B1(\REGISTERS[22][5] ), 
        .B2(n163), .ZN(n1034) );
  OAI221_X1 U1090 ( .B1(n160), .B2(n2080), .C1(n157), .C2(n2048), .A(n1035), 
        .ZN(n1030) );
  AOI22_X1 U1091 ( .A1(\REGISTERS[27][5] ), .A2(n154), .B1(\REGISTERS[26][5] ), 
        .B2(n151), .ZN(n1035) );
  OAI221_X1 U1092 ( .B1(n148), .B2(n2144), .C1(n145), .C2(n2112), .A(n1036), 
        .ZN(n1029) );
  AOI22_X1 U1093 ( .A1(\REGISTERS[29][5] ), .A2(n142), .B1(\REGISTERS[28][5] ), 
        .B2(n139), .ZN(n1036) );
  OAI221_X1 U1094 ( .B1(n115), .B2(n1824), .C1(n112), .C2(n1792), .A(n1043), 
        .ZN(n1038) );
  AOI22_X1 U1095 ( .A1(\REGISTERS[11][5] ), .A2(n109), .B1(\REGISTERS[10][5] ), 
        .B2(n106), .ZN(n1043) );
  OAI221_X1 U1096 ( .B1(n127), .B2(n502), .C1(n124), .C2(n470), .A(n1042), 
        .ZN(n1039) );
  AOI22_X1 U1097 ( .A1(\REGISTERS[7][5] ), .A2(n121), .B1(\REGISTERS[6][5] ), 
        .B2(n118), .ZN(n1042) );
  OAI221_X1 U1098 ( .B1(n103), .B2(n1888), .C1(n100), .C2(n1856), .A(n1044), 
        .ZN(n1037) );
  AOI22_X1 U1099 ( .A1(\REGISTERS[15][5] ), .A2(n97), .B1(\REGISTERS[14][5] ), 
        .B2(n94), .ZN(n1044) );
  OAI221_X1 U1100 ( .B1(n184), .B2(n1951), .C1(n181), .C2(n1919), .A(n1015), 
        .ZN(n1014) );
  AOI22_X1 U1101 ( .A1(\REGISTERS[19][6] ), .A2(n178), .B1(\REGISTERS[18][6] ), 
        .B2(n175), .ZN(n1015) );
  OAI221_X1 U1102 ( .B1(n172), .B2(n2015), .C1(n169), .C2(n1983), .A(n1016), 
        .ZN(n1013) );
  AOI22_X1 U1103 ( .A1(\REGISTERS[23][6] ), .A2(n166), .B1(\REGISTERS[22][6] ), 
        .B2(n163), .ZN(n1016) );
  OAI221_X1 U1104 ( .B1(n160), .B2(n2079), .C1(n157), .C2(n2047), .A(n1017), 
        .ZN(n1012) );
  AOI22_X1 U1105 ( .A1(\REGISTERS[27][6] ), .A2(n154), .B1(\REGISTERS[26][6] ), 
        .B2(n151), .ZN(n1017) );
  OAI221_X1 U1106 ( .B1(n148), .B2(n2143), .C1(n145), .C2(n2111), .A(n1018), 
        .ZN(n1011) );
  AOI22_X1 U1107 ( .A1(\REGISTERS[29][6] ), .A2(n142), .B1(\REGISTERS[28][6] ), 
        .B2(n139), .ZN(n1018) );
  OAI221_X1 U1108 ( .B1(n115), .B2(n1823), .C1(n112), .C2(n1791), .A(n1025), 
        .ZN(n1020) );
  AOI22_X1 U1109 ( .A1(\REGISTERS[11][6] ), .A2(n109), .B1(\REGISTERS[10][6] ), 
        .B2(n106), .ZN(n1025) );
  OAI221_X1 U1110 ( .B1(n127), .B2(n501), .C1(n124), .C2(n469), .A(n1024), 
        .ZN(n1021) );
  AOI22_X1 U1111 ( .A1(\REGISTERS[7][6] ), .A2(n121), .B1(\REGISTERS[6][6] ), 
        .B2(n118), .ZN(n1024) );
  OAI221_X1 U1112 ( .B1(n103), .B2(n1887), .C1(n100), .C2(n1855), .A(n1026), 
        .ZN(n1019) );
  AOI22_X1 U1113 ( .A1(\REGISTERS[15][6] ), .A2(n97), .B1(\REGISTERS[14][6] ), 
        .B2(n94), .ZN(n1026) );
  OAI221_X1 U1114 ( .B1(n184), .B2(n1950), .C1(n181), .C2(n1918), .A(n997), 
        .ZN(n996) );
  AOI22_X1 U1115 ( .A1(\REGISTERS[19][7] ), .A2(n178), .B1(\REGISTERS[18][7] ), 
        .B2(n175), .ZN(n997) );
  OAI221_X1 U1116 ( .B1(n172), .B2(n2014), .C1(n169), .C2(n1982), .A(n998), 
        .ZN(n995) );
  AOI22_X1 U1117 ( .A1(\REGISTERS[23][7] ), .A2(n166), .B1(\REGISTERS[22][7] ), 
        .B2(n163), .ZN(n998) );
  OAI221_X1 U1118 ( .B1(n160), .B2(n2078), .C1(n157), .C2(n2046), .A(n999), 
        .ZN(n994) );
  AOI22_X1 U1119 ( .A1(\REGISTERS[27][7] ), .A2(n154), .B1(\REGISTERS[26][7] ), 
        .B2(n151), .ZN(n999) );
  OAI221_X1 U1120 ( .B1(n148), .B2(n2142), .C1(n145), .C2(n2110), .A(n1000), 
        .ZN(n993) );
  AOI22_X1 U1121 ( .A1(\REGISTERS[29][7] ), .A2(n142), .B1(\REGISTERS[28][7] ), 
        .B2(n139), .ZN(n1000) );
  OAI221_X1 U1122 ( .B1(n115), .B2(n1822), .C1(n112), .C2(n1790), .A(n1007), 
        .ZN(n1002) );
  AOI22_X1 U1123 ( .A1(\REGISTERS[11][7] ), .A2(n109), .B1(\REGISTERS[10][7] ), 
        .B2(n106), .ZN(n1007) );
  OAI221_X1 U1124 ( .B1(n127), .B2(n500), .C1(n124), .C2(n468), .A(n1006), 
        .ZN(n1003) );
  AOI22_X1 U1125 ( .A1(\REGISTERS[7][7] ), .A2(n121), .B1(\REGISTERS[6][7] ), 
        .B2(n118), .ZN(n1006) );
  OAI221_X1 U1126 ( .B1(n103), .B2(n1886), .C1(n100), .C2(n1854), .A(n1008), 
        .ZN(n1001) );
  AOI22_X1 U1127 ( .A1(\REGISTERS[15][7] ), .A2(n97), .B1(\REGISTERS[14][7] ), 
        .B2(n94), .ZN(n1008) );
  OAI221_X1 U1128 ( .B1(n184), .B2(n1949), .C1(n181), .C2(n1917), .A(n979), 
        .ZN(n978) );
  AOI22_X1 U1129 ( .A1(\REGISTERS[19][8] ), .A2(n178), .B1(\REGISTERS[18][8] ), 
        .B2(n175), .ZN(n979) );
  OAI221_X1 U1130 ( .B1(n172), .B2(n2013), .C1(n169), .C2(n1981), .A(n980), 
        .ZN(n977) );
  AOI22_X1 U1131 ( .A1(\REGISTERS[23][8] ), .A2(n166), .B1(\REGISTERS[22][8] ), 
        .B2(n163), .ZN(n980) );
  OAI221_X1 U1132 ( .B1(n160), .B2(n2077), .C1(n157), .C2(n2045), .A(n981), 
        .ZN(n976) );
  AOI22_X1 U1133 ( .A1(\REGISTERS[27][8] ), .A2(n154), .B1(\REGISTERS[26][8] ), 
        .B2(n151), .ZN(n981) );
  OAI221_X1 U1134 ( .B1(n148), .B2(n2141), .C1(n145), .C2(n2109), .A(n982), 
        .ZN(n975) );
  AOI22_X1 U1135 ( .A1(\REGISTERS[29][8] ), .A2(n142), .B1(\REGISTERS[28][8] ), 
        .B2(n139), .ZN(n982) );
  OAI221_X1 U1136 ( .B1(n115), .B2(n1821), .C1(n112), .C2(n1789), .A(n989), 
        .ZN(n984) );
  AOI22_X1 U1137 ( .A1(\REGISTERS[11][8] ), .A2(n109), .B1(\REGISTERS[10][8] ), 
        .B2(n106), .ZN(n989) );
  OAI221_X1 U1138 ( .B1(n127), .B2(n499), .C1(n124), .C2(n467), .A(n988), .ZN(
        n985) );
  AOI22_X1 U1139 ( .A1(\REGISTERS[7][8] ), .A2(n121), .B1(\REGISTERS[6][8] ), 
        .B2(n118), .ZN(n988) );
  OAI221_X1 U1140 ( .B1(n103), .B2(n1885), .C1(n100), .C2(n1853), .A(n990), 
        .ZN(n983) );
  AOI22_X1 U1141 ( .A1(\REGISTERS[15][8] ), .A2(n97), .B1(\REGISTERS[14][8] ), 
        .B2(n94), .ZN(n990) );
  OAI221_X1 U1142 ( .B1(n184), .B2(n1948), .C1(n181), .C2(n1916), .A(n961), 
        .ZN(n960) );
  AOI22_X1 U1143 ( .A1(\REGISTERS[19][9] ), .A2(n178), .B1(\REGISTERS[18][9] ), 
        .B2(n175), .ZN(n961) );
  OAI221_X1 U1144 ( .B1(n172), .B2(n2012), .C1(n169), .C2(n1980), .A(n962), 
        .ZN(n959) );
  AOI22_X1 U1145 ( .A1(\REGISTERS[23][9] ), .A2(n166), .B1(\REGISTERS[22][9] ), 
        .B2(n163), .ZN(n962) );
  OAI221_X1 U1146 ( .B1(n160), .B2(n2076), .C1(n157), .C2(n2044), .A(n963), 
        .ZN(n958) );
  AOI22_X1 U1147 ( .A1(\REGISTERS[27][9] ), .A2(n154), .B1(\REGISTERS[26][9] ), 
        .B2(n151), .ZN(n963) );
  OAI221_X1 U1148 ( .B1(n148), .B2(n2140), .C1(n145), .C2(n2108), .A(n964), 
        .ZN(n957) );
  AOI22_X1 U1149 ( .A1(\REGISTERS[29][9] ), .A2(n142), .B1(\REGISTERS[28][9] ), 
        .B2(n139), .ZN(n964) );
  OAI221_X1 U1150 ( .B1(n115), .B2(n1820), .C1(n112), .C2(n1788), .A(n971), 
        .ZN(n966) );
  AOI22_X1 U1151 ( .A1(\REGISTERS[11][9] ), .A2(n109), .B1(\REGISTERS[10][9] ), 
        .B2(n106), .ZN(n971) );
  OAI221_X1 U1152 ( .B1(n127), .B2(n498), .C1(n124), .C2(n466), .A(n970), .ZN(
        n967) );
  AOI22_X1 U1153 ( .A1(\REGISTERS[7][9] ), .A2(n121), .B1(\REGISTERS[6][9] ), 
        .B2(n118), .ZN(n970) );
  OAI221_X1 U1154 ( .B1(n103), .B2(n1884), .C1(n100), .C2(n1852), .A(n972), 
        .ZN(n965) );
  AOI22_X1 U1155 ( .A1(\REGISTERS[15][9] ), .A2(n97), .B1(\REGISTERS[14][9] ), 
        .B2(n94), .ZN(n972) );
  OAI221_X1 U1156 ( .B1(n184), .B2(n1947), .C1(n181), .C2(n1915), .A(n943), 
        .ZN(n942) );
  AOI22_X1 U1157 ( .A1(\REGISTERS[19][10] ), .A2(n178), .B1(
        \REGISTERS[18][10] ), .B2(n175), .ZN(n943) );
  OAI221_X1 U1158 ( .B1(n172), .B2(n2011), .C1(n169), .C2(n1979), .A(n944), 
        .ZN(n941) );
  AOI22_X1 U1159 ( .A1(\REGISTERS[23][10] ), .A2(n166), .B1(
        \REGISTERS[22][10] ), .B2(n163), .ZN(n944) );
  OAI221_X1 U1160 ( .B1(n160), .B2(n2075), .C1(n157), .C2(n2043), .A(n945), 
        .ZN(n940) );
  AOI22_X1 U1161 ( .A1(\REGISTERS[27][10] ), .A2(n154), .B1(
        \REGISTERS[26][10] ), .B2(n151), .ZN(n945) );
  OAI221_X1 U1162 ( .B1(n148), .B2(n2139), .C1(n145), .C2(n2107), .A(n946), 
        .ZN(n939) );
  AOI22_X1 U1163 ( .A1(\REGISTERS[29][10] ), .A2(n142), .B1(
        \REGISTERS[28][10] ), .B2(n139), .ZN(n946) );
  OAI221_X1 U1164 ( .B1(n115), .B2(n1819), .C1(n112), .C2(n1787), .A(n953), 
        .ZN(n948) );
  AOI22_X1 U1165 ( .A1(\REGISTERS[11][10] ), .A2(n109), .B1(
        \REGISTERS[10][10] ), .B2(n106), .ZN(n953) );
  OAI221_X1 U1166 ( .B1(n127), .B2(n497), .C1(n124), .C2(n465), .A(n952), .ZN(
        n949) );
  AOI22_X1 U1167 ( .A1(\REGISTERS[7][10] ), .A2(n121), .B1(\REGISTERS[6][10] ), 
        .B2(n118), .ZN(n952) );
  OAI221_X1 U1168 ( .B1(n103), .B2(n1883), .C1(n100), .C2(n1851), .A(n954), 
        .ZN(n947) );
  AOI22_X1 U1169 ( .A1(\REGISTERS[15][10] ), .A2(n97), .B1(\REGISTERS[14][10] ), .B2(n94), .ZN(n954) );
  OAI221_X1 U1170 ( .B1(n184), .B2(n1946), .C1(n181), .C2(n1914), .A(n925), 
        .ZN(n924) );
  AOI22_X1 U1171 ( .A1(\REGISTERS[19][11] ), .A2(n178), .B1(
        \REGISTERS[18][11] ), .B2(n175), .ZN(n925) );
  OAI221_X1 U1172 ( .B1(n172), .B2(n2010), .C1(n169), .C2(n1978), .A(n926), 
        .ZN(n923) );
  AOI22_X1 U1173 ( .A1(\REGISTERS[23][11] ), .A2(n166), .B1(
        \REGISTERS[22][11] ), .B2(n163), .ZN(n926) );
  OAI221_X1 U1174 ( .B1(n160), .B2(n2074), .C1(n157), .C2(n2042), .A(n927), 
        .ZN(n922) );
  AOI22_X1 U1175 ( .A1(\REGISTERS[27][11] ), .A2(n154), .B1(
        \REGISTERS[26][11] ), .B2(n151), .ZN(n927) );
  OAI221_X1 U1176 ( .B1(n148), .B2(n2138), .C1(n145), .C2(n2106), .A(n928), 
        .ZN(n921) );
  AOI22_X1 U1177 ( .A1(\REGISTERS[29][11] ), .A2(n142), .B1(
        \REGISTERS[28][11] ), .B2(n139), .ZN(n928) );
  OAI221_X1 U1178 ( .B1(n115), .B2(n1818), .C1(n112), .C2(n1182), .A(n935), 
        .ZN(n930) );
  AOI22_X1 U1179 ( .A1(\REGISTERS[11][11] ), .A2(n109), .B1(
        \REGISTERS[10][11] ), .B2(n106), .ZN(n935) );
  OAI221_X1 U1180 ( .B1(n127), .B2(n496), .C1(n124), .C2(n464), .A(n934), .ZN(
        n931) );
  AOI22_X1 U1181 ( .A1(\REGISTERS[7][11] ), .A2(n121), .B1(\REGISTERS[6][11] ), 
        .B2(n118), .ZN(n934) );
  OAI221_X1 U1182 ( .B1(n103), .B2(n1882), .C1(n100), .C2(n1850), .A(n936), 
        .ZN(n929) );
  AOI22_X1 U1183 ( .A1(\REGISTERS[15][11] ), .A2(n97), .B1(\REGISTERS[14][11] ), .B2(n94), .ZN(n936) );
  OAI221_X1 U1184 ( .B1(n185), .B2(n1945), .C1(n182), .C2(n1913), .A(n907), 
        .ZN(n906) );
  AOI22_X1 U1185 ( .A1(\REGISTERS[19][12] ), .A2(n179), .B1(
        \REGISTERS[18][12] ), .B2(n176), .ZN(n907) );
  OAI221_X1 U1186 ( .B1(n173), .B2(n2009), .C1(n170), .C2(n1977), .A(n908), 
        .ZN(n905) );
  AOI22_X1 U1187 ( .A1(\REGISTERS[23][12] ), .A2(n167), .B1(
        \REGISTERS[22][12] ), .B2(n164), .ZN(n908) );
  OAI221_X1 U1188 ( .B1(n161), .B2(n2073), .C1(n158), .C2(n2041), .A(n909), 
        .ZN(n904) );
  AOI22_X1 U1189 ( .A1(\REGISTERS[27][12] ), .A2(n155), .B1(
        \REGISTERS[26][12] ), .B2(n152), .ZN(n909) );
  OAI221_X1 U1190 ( .B1(n149), .B2(n2137), .C1(n146), .C2(n2105), .A(n910), 
        .ZN(n903) );
  AOI22_X1 U1191 ( .A1(\REGISTERS[29][12] ), .A2(n143), .B1(
        \REGISTERS[28][12] ), .B2(n140), .ZN(n910) );
  OAI221_X1 U1192 ( .B1(n116), .B2(n1817), .C1(n113), .C2(n558), .A(n917), 
        .ZN(n912) );
  AOI22_X1 U1193 ( .A1(\REGISTERS[11][12] ), .A2(n110), .B1(
        \REGISTERS[10][12] ), .B2(n107), .ZN(n917) );
  OAI221_X1 U1194 ( .B1(n128), .B2(n495), .C1(n125), .C2(n463), .A(n916), .ZN(
        n913) );
  AOI22_X1 U1195 ( .A1(\REGISTERS[7][12] ), .A2(n122), .B1(\REGISTERS[6][12] ), 
        .B2(n119), .ZN(n916) );
  OAI221_X1 U1196 ( .B1(n104), .B2(n1881), .C1(n101), .C2(n1849), .A(n918), 
        .ZN(n911) );
  AOI22_X1 U1197 ( .A1(\REGISTERS[15][12] ), .A2(n98), .B1(\REGISTERS[14][12] ), .B2(n95), .ZN(n918) );
  OAI221_X1 U1198 ( .B1(n185), .B2(n1944), .C1(n182), .C2(n1912), .A(n889), 
        .ZN(n888) );
  AOI22_X1 U1199 ( .A1(\REGISTERS[19][13] ), .A2(n179), .B1(
        \REGISTERS[18][13] ), .B2(n176), .ZN(n889) );
  OAI221_X1 U1200 ( .B1(n173), .B2(n2008), .C1(n170), .C2(n1976), .A(n890), 
        .ZN(n887) );
  AOI22_X1 U1201 ( .A1(\REGISTERS[23][13] ), .A2(n167), .B1(
        \REGISTERS[22][13] ), .B2(n164), .ZN(n890) );
  OAI221_X1 U1202 ( .B1(n161), .B2(n2072), .C1(n158), .C2(n2040), .A(n891), 
        .ZN(n886) );
  AOI22_X1 U1203 ( .A1(\REGISTERS[27][13] ), .A2(n155), .B1(
        \REGISTERS[26][13] ), .B2(n152), .ZN(n891) );
  OAI221_X1 U1204 ( .B1(n149), .B2(n2136), .C1(n146), .C2(n2104), .A(n892), 
        .ZN(n885) );
  AOI22_X1 U1205 ( .A1(\REGISTERS[29][13] ), .A2(n143), .B1(
        \REGISTERS[28][13] ), .B2(n140), .ZN(n892) );
  OAI221_X1 U1206 ( .B1(n116), .B2(n1816), .C1(n113), .C2(n526), .A(n899), 
        .ZN(n894) );
  AOI22_X1 U1207 ( .A1(\REGISTERS[11][13] ), .A2(n110), .B1(
        \REGISTERS[10][13] ), .B2(n107), .ZN(n899) );
  OAI221_X1 U1208 ( .B1(n128), .B2(n494), .C1(n125), .C2(n462), .A(n898), .ZN(
        n895) );
  AOI22_X1 U1209 ( .A1(\REGISTERS[7][13] ), .A2(n122), .B1(\REGISTERS[6][13] ), 
        .B2(n119), .ZN(n898) );
  OAI221_X1 U1210 ( .B1(n104), .B2(n1880), .C1(n101), .C2(n1848), .A(n900), 
        .ZN(n893) );
  AOI22_X1 U1211 ( .A1(\REGISTERS[15][13] ), .A2(n98), .B1(\REGISTERS[14][13] ), .B2(n95), .ZN(n900) );
  OAI221_X1 U1212 ( .B1(n185), .B2(n1943), .C1(n182), .C2(n1911), .A(n871), 
        .ZN(n870) );
  AOI22_X1 U1213 ( .A1(\REGISTERS[19][14] ), .A2(n179), .B1(
        \REGISTERS[18][14] ), .B2(n176), .ZN(n871) );
  OAI221_X1 U1214 ( .B1(n173), .B2(n2007), .C1(n170), .C2(n1975), .A(n872), 
        .ZN(n869) );
  AOI22_X1 U1215 ( .A1(\REGISTERS[23][14] ), .A2(n167), .B1(
        \REGISTERS[22][14] ), .B2(n164), .ZN(n872) );
  OAI221_X1 U1216 ( .B1(n161), .B2(n2071), .C1(n158), .C2(n2039), .A(n873), 
        .ZN(n868) );
  AOI22_X1 U1217 ( .A1(\REGISTERS[27][14] ), .A2(n155), .B1(
        \REGISTERS[26][14] ), .B2(n152), .ZN(n873) );
  OAI221_X1 U1218 ( .B1(n149), .B2(n2135), .C1(n146), .C2(n2103), .A(n874), 
        .ZN(n867) );
  AOI22_X1 U1219 ( .A1(\REGISTERS[29][14] ), .A2(n143), .B1(
        \REGISTERS[28][14] ), .B2(n140), .ZN(n874) );
  OAI221_X1 U1220 ( .B1(n116), .B2(n1815), .C1(n113), .C2(n525), .A(n881), 
        .ZN(n876) );
  AOI22_X1 U1221 ( .A1(\REGISTERS[11][14] ), .A2(n110), .B1(
        \REGISTERS[10][14] ), .B2(n107), .ZN(n881) );
  OAI221_X1 U1222 ( .B1(n128), .B2(n493), .C1(n125), .C2(n461), .A(n880), .ZN(
        n877) );
  AOI22_X1 U1223 ( .A1(\REGISTERS[7][14] ), .A2(n122), .B1(\REGISTERS[6][14] ), 
        .B2(n119), .ZN(n880) );
  OAI221_X1 U1224 ( .B1(n104), .B2(n1879), .C1(n101), .C2(n1847), .A(n882), 
        .ZN(n875) );
  AOI22_X1 U1225 ( .A1(\REGISTERS[15][14] ), .A2(n98), .B1(\REGISTERS[14][14] ), .B2(n95), .ZN(n882) );
  OAI221_X1 U1226 ( .B1(n185), .B2(n1942), .C1(n182), .C2(n1910), .A(n853), 
        .ZN(n852) );
  AOI22_X1 U1227 ( .A1(\REGISTERS[19][15] ), .A2(n179), .B1(
        \REGISTERS[18][15] ), .B2(n176), .ZN(n853) );
  OAI221_X1 U1228 ( .B1(n173), .B2(n2006), .C1(n170), .C2(n1974), .A(n854), 
        .ZN(n851) );
  AOI22_X1 U1229 ( .A1(\REGISTERS[23][15] ), .A2(n167), .B1(
        \REGISTERS[22][15] ), .B2(n164), .ZN(n854) );
  OAI221_X1 U1230 ( .B1(n161), .B2(n2070), .C1(n158), .C2(n2038), .A(n855), 
        .ZN(n850) );
  AOI22_X1 U1231 ( .A1(\REGISTERS[27][15] ), .A2(n155), .B1(
        \REGISTERS[26][15] ), .B2(n152), .ZN(n855) );
  OAI221_X1 U1232 ( .B1(n149), .B2(n2134), .C1(n146), .C2(n2102), .A(n856), 
        .ZN(n849) );
  AOI22_X1 U1233 ( .A1(\REGISTERS[29][15] ), .A2(n143), .B1(
        \REGISTERS[28][15] ), .B2(n140), .ZN(n856) );
  OAI221_X1 U1234 ( .B1(n116), .B2(n1814), .C1(n113), .C2(n524), .A(n863), 
        .ZN(n858) );
  AOI22_X1 U1235 ( .A1(\REGISTERS[11][15] ), .A2(n110), .B1(
        \REGISTERS[10][15] ), .B2(n107), .ZN(n863) );
  OAI221_X1 U1236 ( .B1(n128), .B2(n492), .C1(n125), .C2(n460), .A(n862), .ZN(
        n859) );
  AOI22_X1 U1237 ( .A1(\REGISTERS[7][15] ), .A2(n122), .B1(\REGISTERS[6][15] ), 
        .B2(n119), .ZN(n862) );
  OAI221_X1 U1238 ( .B1(n104), .B2(n1878), .C1(n101), .C2(n1846), .A(n864), 
        .ZN(n857) );
  AOI22_X1 U1239 ( .A1(\REGISTERS[15][15] ), .A2(n98), .B1(\REGISTERS[14][15] ), .B2(n95), .ZN(n864) );
  OAI221_X1 U1240 ( .B1(n185), .B2(n1941), .C1(n182), .C2(n1909), .A(n835), 
        .ZN(n834) );
  AOI22_X1 U1241 ( .A1(\REGISTERS[19][16] ), .A2(n179), .B1(
        \REGISTERS[18][16] ), .B2(n176), .ZN(n835) );
  OAI221_X1 U1242 ( .B1(n173), .B2(n2005), .C1(n170), .C2(n1973), .A(n836), 
        .ZN(n833) );
  AOI22_X1 U1243 ( .A1(\REGISTERS[23][16] ), .A2(n167), .B1(
        \REGISTERS[22][16] ), .B2(n164), .ZN(n836) );
  OAI221_X1 U1244 ( .B1(n161), .B2(n2069), .C1(n158), .C2(n2037), .A(n837), 
        .ZN(n832) );
  AOI22_X1 U1245 ( .A1(\REGISTERS[27][16] ), .A2(n155), .B1(
        \REGISTERS[26][16] ), .B2(n152), .ZN(n837) );
  OAI221_X1 U1246 ( .B1(n149), .B2(n2133), .C1(n146), .C2(n2101), .A(n838), 
        .ZN(n831) );
  AOI22_X1 U1247 ( .A1(\REGISTERS[29][16] ), .A2(n143), .B1(
        \REGISTERS[28][16] ), .B2(n140), .ZN(n838) );
  OAI221_X1 U1248 ( .B1(n116), .B2(n1813), .C1(n113), .C2(n523), .A(n845), 
        .ZN(n840) );
  AOI22_X1 U1249 ( .A1(\REGISTERS[11][16] ), .A2(n110), .B1(
        \REGISTERS[10][16] ), .B2(n107), .ZN(n845) );
  OAI221_X1 U1250 ( .B1(n128), .B2(n491), .C1(n125), .C2(n459), .A(n844), .ZN(
        n841) );
  AOI22_X1 U1251 ( .A1(\REGISTERS[7][16] ), .A2(n122), .B1(\REGISTERS[6][16] ), 
        .B2(n119), .ZN(n844) );
  OAI221_X1 U1252 ( .B1(n104), .B2(n1877), .C1(n101), .C2(n1845), .A(n846), 
        .ZN(n839) );
  AOI22_X1 U1253 ( .A1(\REGISTERS[15][16] ), .A2(n98), .B1(\REGISTERS[14][16] ), .B2(n95), .ZN(n846) );
  OAI221_X1 U1254 ( .B1(n185), .B2(n1940), .C1(n182), .C2(n1908), .A(n817), 
        .ZN(n816) );
  AOI22_X1 U1255 ( .A1(\REGISTERS[19][17] ), .A2(n179), .B1(
        \REGISTERS[18][17] ), .B2(n176), .ZN(n817) );
  OAI221_X1 U1256 ( .B1(n173), .B2(n2004), .C1(n170), .C2(n1972), .A(n818), 
        .ZN(n815) );
  AOI22_X1 U1257 ( .A1(\REGISTERS[23][17] ), .A2(n167), .B1(
        \REGISTERS[22][17] ), .B2(n164), .ZN(n818) );
  OAI221_X1 U1258 ( .B1(n161), .B2(n2068), .C1(n158), .C2(n2036), .A(n819), 
        .ZN(n814) );
  AOI22_X1 U1259 ( .A1(\REGISTERS[27][17] ), .A2(n155), .B1(
        \REGISTERS[26][17] ), .B2(n152), .ZN(n819) );
  OAI221_X1 U1260 ( .B1(n149), .B2(n2132), .C1(n146), .C2(n2100), .A(n820), 
        .ZN(n813) );
  AOI22_X1 U1261 ( .A1(\REGISTERS[29][17] ), .A2(n143), .B1(
        \REGISTERS[28][17] ), .B2(n140), .ZN(n820) );
  OAI221_X1 U1262 ( .B1(n116), .B2(n1812), .C1(n113), .C2(n522), .A(n827), 
        .ZN(n822) );
  AOI22_X1 U1263 ( .A1(\REGISTERS[11][17] ), .A2(n110), .B1(
        \REGISTERS[10][17] ), .B2(n107), .ZN(n827) );
  OAI221_X1 U1264 ( .B1(n128), .B2(n490), .C1(n125), .C2(n458), .A(n826), .ZN(
        n823) );
  AOI22_X1 U1265 ( .A1(\REGISTERS[7][17] ), .A2(n122), .B1(\REGISTERS[6][17] ), 
        .B2(n119), .ZN(n826) );
  OAI221_X1 U1266 ( .B1(n104), .B2(n1876), .C1(n101), .C2(n1844), .A(n828), 
        .ZN(n821) );
  AOI22_X1 U1267 ( .A1(\REGISTERS[15][17] ), .A2(n98), .B1(\REGISTERS[14][17] ), .B2(n95), .ZN(n828) );
  OAI221_X1 U1268 ( .B1(n185), .B2(n1939), .C1(n182), .C2(n1907), .A(n799), 
        .ZN(n798) );
  AOI22_X1 U1269 ( .A1(\REGISTERS[19][18] ), .A2(n179), .B1(
        \REGISTERS[18][18] ), .B2(n176), .ZN(n799) );
  OAI221_X1 U1270 ( .B1(n173), .B2(n2003), .C1(n170), .C2(n1971), .A(n800), 
        .ZN(n797) );
  AOI22_X1 U1271 ( .A1(\REGISTERS[23][18] ), .A2(n167), .B1(
        \REGISTERS[22][18] ), .B2(n164), .ZN(n800) );
  OAI221_X1 U1272 ( .B1(n161), .B2(n2067), .C1(n158), .C2(n2035), .A(n801), 
        .ZN(n796) );
  AOI22_X1 U1273 ( .A1(\REGISTERS[27][18] ), .A2(n155), .B1(
        \REGISTERS[26][18] ), .B2(n152), .ZN(n801) );
  OAI221_X1 U1274 ( .B1(n149), .B2(n2131), .C1(n146), .C2(n2099), .A(n802), 
        .ZN(n795) );
  AOI22_X1 U1275 ( .A1(\REGISTERS[29][18] ), .A2(n143), .B1(
        \REGISTERS[28][18] ), .B2(n140), .ZN(n802) );
  OAI221_X1 U1276 ( .B1(n116), .B2(n1811), .C1(n113), .C2(n521), .A(n809), 
        .ZN(n804) );
  AOI22_X1 U1277 ( .A1(\REGISTERS[11][18] ), .A2(n110), .B1(
        \REGISTERS[10][18] ), .B2(n107), .ZN(n809) );
  OAI221_X1 U1278 ( .B1(n128), .B2(n489), .C1(n125), .C2(n457), .A(n808), .ZN(
        n805) );
  AOI22_X1 U1279 ( .A1(\REGISTERS[7][18] ), .A2(n122), .B1(\REGISTERS[6][18] ), 
        .B2(n119), .ZN(n808) );
  OAI221_X1 U1280 ( .B1(n104), .B2(n1875), .C1(n101), .C2(n1843), .A(n810), 
        .ZN(n803) );
  AOI22_X1 U1281 ( .A1(\REGISTERS[15][18] ), .A2(n98), .B1(\REGISTERS[14][18] ), .B2(n95), .ZN(n810) );
  OAI221_X1 U1282 ( .B1(n185), .B2(n1938), .C1(n182), .C2(n1906), .A(n781), 
        .ZN(n780) );
  AOI22_X1 U1283 ( .A1(\REGISTERS[19][19] ), .A2(n179), .B1(
        \REGISTERS[18][19] ), .B2(n176), .ZN(n781) );
  OAI221_X1 U1284 ( .B1(n173), .B2(n2002), .C1(n170), .C2(n1970), .A(n782), 
        .ZN(n779) );
  AOI22_X1 U1285 ( .A1(\REGISTERS[23][19] ), .A2(n167), .B1(
        \REGISTERS[22][19] ), .B2(n164), .ZN(n782) );
  OAI221_X1 U1286 ( .B1(n161), .B2(n2066), .C1(n158), .C2(n2034), .A(n783), 
        .ZN(n778) );
  AOI22_X1 U1287 ( .A1(\REGISTERS[27][19] ), .A2(n155), .B1(
        \REGISTERS[26][19] ), .B2(n152), .ZN(n783) );
  OAI221_X1 U1288 ( .B1(n149), .B2(n2130), .C1(n146), .C2(n2098), .A(n784), 
        .ZN(n777) );
  AOI22_X1 U1289 ( .A1(\REGISTERS[29][19] ), .A2(n143), .B1(
        \REGISTERS[28][19] ), .B2(n140), .ZN(n784) );
  OAI221_X1 U1290 ( .B1(n116), .B2(n1810), .C1(n113), .C2(n520), .A(n791), 
        .ZN(n786) );
  AOI22_X1 U1291 ( .A1(\REGISTERS[11][19] ), .A2(n110), .B1(
        \REGISTERS[10][19] ), .B2(n107), .ZN(n791) );
  OAI221_X1 U1292 ( .B1(n128), .B2(n488), .C1(n125), .C2(n456), .A(n790), .ZN(
        n787) );
  AOI22_X1 U1293 ( .A1(\REGISTERS[7][19] ), .A2(n122), .B1(\REGISTERS[6][19] ), 
        .B2(n119), .ZN(n790) );
  OAI221_X1 U1294 ( .B1(n104), .B2(n1874), .C1(n101), .C2(n1842), .A(n792), 
        .ZN(n785) );
  AOI22_X1 U1295 ( .A1(\REGISTERS[15][19] ), .A2(n98), .B1(\REGISTERS[14][19] ), .B2(n95), .ZN(n792) );
  OAI221_X1 U1296 ( .B1(n185), .B2(n1937), .C1(n182), .C2(n1905), .A(n763), 
        .ZN(n762) );
  AOI22_X1 U1297 ( .A1(\REGISTERS[19][20] ), .A2(n179), .B1(
        \REGISTERS[18][20] ), .B2(n176), .ZN(n763) );
  OAI221_X1 U1298 ( .B1(n173), .B2(n2001), .C1(n170), .C2(n1969), .A(n764), 
        .ZN(n761) );
  AOI22_X1 U1299 ( .A1(\REGISTERS[23][20] ), .A2(n167), .B1(
        \REGISTERS[22][20] ), .B2(n164), .ZN(n764) );
  OAI221_X1 U1300 ( .B1(n161), .B2(n2065), .C1(n158), .C2(n2033), .A(n765), 
        .ZN(n760) );
  AOI22_X1 U1301 ( .A1(\REGISTERS[27][20] ), .A2(n155), .B1(
        \REGISTERS[26][20] ), .B2(n152), .ZN(n765) );
  OAI221_X1 U1302 ( .B1(n149), .B2(n2129), .C1(n146), .C2(n2097), .A(n766), 
        .ZN(n759) );
  AOI22_X1 U1303 ( .A1(\REGISTERS[29][20] ), .A2(n143), .B1(
        \REGISTERS[28][20] ), .B2(n140), .ZN(n766) );
  OAI221_X1 U1304 ( .B1(n116), .B2(n1809), .C1(n113), .C2(n519), .A(n773), 
        .ZN(n768) );
  AOI22_X1 U1305 ( .A1(\REGISTERS[11][20] ), .A2(n110), .B1(
        \REGISTERS[10][20] ), .B2(n107), .ZN(n773) );
  OAI221_X1 U1306 ( .B1(n128), .B2(n487), .C1(n125), .C2(n455), .A(n772), .ZN(
        n769) );
  AOI22_X1 U1307 ( .A1(\REGISTERS[7][20] ), .A2(n122), .B1(\REGISTERS[6][20] ), 
        .B2(n119), .ZN(n772) );
  OAI221_X1 U1308 ( .B1(n104), .B2(n1873), .C1(n101), .C2(n1841), .A(n774), 
        .ZN(n767) );
  AOI22_X1 U1309 ( .A1(\REGISTERS[15][20] ), .A2(n98), .B1(\REGISTERS[14][20] ), .B2(n95), .ZN(n774) );
  OAI221_X1 U1310 ( .B1(n185), .B2(n1936), .C1(n182), .C2(n1904), .A(n745), 
        .ZN(n744) );
  AOI22_X1 U1311 ( .A1(\REGISTERS[19][21] ), .A2(n179), .B1(
        \REGISTERS[18][21] ), .B2(n176), .ZN(n745) );
  OAI221_X1 U1312 ( .B1(n173), .B2(n2000), .C1(n170), .C2(n1968), .A(n746), 
        .ZN(n743) );
  AOI22_X1 U1313 ( .A1(\REGISTERS[23][21] ), .A2(n167), .B1(
        \REGISTERS[22][21] ), .B2(n164), .ZN(n746) );
  OAI221_X1 U1314 ( .B1(n161), .B2(n2064), .C1(n158), .C2(n2032), .A(n747), 
        .ZN(n742) );
  AOI22_X1 U1315 ( .A1(\REGISTERS[27][21] ), .A2(n155), .B1(
        \REGISTERS[26][21] ), .B2(n152), .ZN(n747) );
  OAI221_X1 U1316 ( .B1(n149), .B2(n2128), .C1(n146), .C2(n2096), .A(n748), 
        .ZN(n741) );
  AOI22_X1 U1317 ( .A1(\REGISTERS[29][21] ), .A2(n143), .B1(
        \REGISTERS[28][21] ), .B2(n140), .ZN(n748) );
  OAI221_X1 U1318 ( .B1(n116), .B2(n1808), .C1(n113), .C2(n518), .A(n755), 
        .ZN(n750) );
  AOI22_X1 U1319 ( .A1(\REGISTERS[11][21] ), .A2(n110), .B1(
        \REGISTERS[10][21] ), .B2(n107), .ZN(n755) );
  OAI221_X1 U1320 ( .B1(n128), .B2(n486), .C1(n125), .C2(n454), .A(n754), .ZN(
        n751) );
  AOI22_X1 U1321 ( .A1(\REGISTERS[7][21] ), .A2(n122), .B1(\REGISTERS[6][21] ), 
        .B2(n119), .ZN(n754) );
  OAI221_X1 U1322 ( .B1(n104), .B2(n1872), .C1(n101), .C2(n1840), .A(n756), 
        .ZN(n749) );
  AOI22_X1 U1323 ( .A1(\REGISTERS[15][21] ), .A2(n98), .B1(\REGISTERS[14][21] ), .B2(n95), .ZN(n756) );
  OAI221_X1 U1324 ( .B1(n185), .B2(n1935), .C1(n182), .C2(n1903), .A(n727), 
        .ZN(n726) );
  AOI22_X1 U1325 ( .A1(\REGISTERS[19][22] ), .A2(n179), .B1(
        \REGISTERS[18][22] ), .B2(n176), .ZN(n727) );
  OAI221_X1 U1326 ( .B1(n173), .B2(n1999), .C1(n170), .C2(n1967), .A(n728), 
        .ZN(n725) );
  AOI22_X1 U1327 ( .A1(\REGISTERS[23][22] ), .A2(n167), .B1(
        \REGISTERS[22][22] ), .B2(n164), .ZN(n728) );
  OAI221_X1 U1328 ( .B1(n161), .B2(n2063), .C1(n158), .C2(n2031), .A(n729), 
        .ZN(n724) );
  AOI22_X1 U1329 ( .A1(\REGISTERS[27][22] ), .A2(n155), .B1(
        \REGISTERS[26][22] ), .B2(n152), .ZN(n729) );
  OAI221_X1 U1330 ( .B1(n149), .B2(n2127), .C1(n146), .C2(n2095), .A(n730), 
        .ZN(n723) );
  AOI22_X1 U1331 ( .A1(\REGISTERS[29][22] ), .A2(n143), .B1(
        \REGISTERS[28][22] ), .B2(n140), .ZN(n730) );
  OAI221_X1 U1332 ( .B1(n116), .B2(n1807), .C1(n113), .C2(n517), .A(n737), 
        .ZN(n732) );
  AOI22_X1 U1333 ( .A1(\REGISTERS[11][22] ), .A2(n110), .B1(
        \REGISTERS[10][22] ), .B2(n107), .ZN(n737) );
  OAI221_X1 U1334 ( .B1(n128), .B2(n485), .C1(n125), .C2(n453), .A(n736), .ZN(
        n733) );
  AOI22_X1 U1335 ( .A1(\REGISTERS[7][22] ), .A2(n122), .B1(\REGISTERS[6][22] ), 
        .B2(n119), .ZN(n736) );
  OAI221_X1 U1336 ( .B1(n104), .B2(n1871), .C1(n101), .C2(n1839), .A(n738), 
        .ZN(n731) );
  AOI22_X1 U1337 ( .A1(\REGISTERS[15][22] ), .A2(n98), .B1(\REGISTERS[14][22] ), .B2(n95), .ZN(n738) );
  OAI221_X1 U1338 ( .B1(n185), .B2(n1934), .C1(n182), .C2(n1902), .A(n709), 
        .ZN(n708) );
  AOI22_X1 U1339 ( .A1(\REGISTERS[19][23] ), .A2(n179), .B1(
        \REGISTERS[18][23] ), .B2(n176), .ZN(n709) );
  OAI221_X1 U1340 ( .B1(n173), .B2(n1998), .C1(n170), .C2(n1966), .A(n710), 
        .ZN(n707) );
  AOI22_X1 U1341 ( .A1(\REGISTERS[23][23] ), .A2(n167), .B1(
        \REGISTERS[22][23] ), .B2(n164), .ZN(n710) );
  OAI221_X1 U1342 ( .B1(n161), .B2(n2062), .C1(n158), .C2(n2030), .A(n711), 
        .ZN(n706) );
  AOI22_X1 U1343 ( .A1(\REGISTERS[27][23] ), .A2(n155), .B1(
        \REGISTERS[26][23] ), .B2(n152), .ZN(n711) );
  OAI221_X1 U1344 ( .B1(n149), .B2(n2126), .C1(n146), .C2(n2094), .A(n712), 
        .ZN(n705) );
  AOI22_X1 U1345 ( .A1(\REGISTERS[29][23] ), .A2(n143), .B1(
        \REGISTERS[28][23] ), .B2(n140), .ZN(n712) );
  OAI221_X1 U1346 ( .B1(n116), .B2(n1806), .C1(n113), .C2(n516), .A(n719), 
        .ZN(n714) );
  AOI22_X1 U1347 ( .A1(\REGISTERS[11][23] ), .A2(n110), .B1(
        \REGISTERS[10][23] ), .B2(n107), .ZN(n719) );
  OAI221_X1 U1348 ( .B1(n128), .B2(n484), .C1(n125), .C2(n452), .A(n718), .ZN(
        n715) );
  AOI22_X1 U1349 ( .A1(\REGISTERS[7][23] ), .A2(n122), .B1(\REGISTERS[6][23] ), 
        .B2(n119), .ZN(n718) );
  OAI221_X1 U1350 ( .B1(n104), .B2(n1870), .C1(n101), .C2(n1838), .A(n720), 
        .ZN(n713) );
  AOI22_X1 U1351 ( .A1(\REGISTERS[15][23] ), .A2(n98), .B1(\REGISTERS[14][23] ), .B2(n95), .ZN(n720) );
  OAI221_X1 U1352 ( .B1(n1957), .B2(n91), .C1(n1925), .C2(n88), .A(n1747), 
        .ZN(n1746) );
  AOI22_X1 U1353 ( .A1(n85), .A2(\REGISTERS[19][0] ), .B1(n84), .B2(
        \REGISTERS[18][0] ), .ZN(n1747) );
  OAI221_X1 U1354 ( .B1(n2021), .B2(n79), .C1(n1989), .C2(n76), .A(n1752), 
        .ZN(n1745) );
  AOI22_X1 U1355 ( .A1(n73), .A2(\REGISTERS[23][0] ), .B1(n72), .B2(
        \REGISTERS[22][0] ), .ZN(n1752) );
  OAI221_X1 U1356 ( .B1(n2085), .B2(n67), .C1(n2053), .C2(n64), .A(n1756), 
        .ZN(n1744) );
  AOI22_X1 U1357 ( .A1(n61), .A2(\REGISTERS[27][0] ), .B1(n60), .B2(
        \REGISTERS[26][0] ), .ZN(n1756) );
  OAI221_X1 U1358 ( .B1(n2149), .B2(n55), .C1(n2117), .C2(n52), .A(n1759), 
        .ZN(n1743) );
  AOI22_X1 U1359 ( .A1(n49), .A2(\REGISTERS[29][0] ), .B1(n48), .B2(
        \REGISTERS[28][0] ), .ZN(n1759) );
  OAI221_X1 U1360 ( .B1(n507), .B2(n34), .C1(n475), .C2(n31), .A(n1768), .ZN(
        n1763) );
  AOI22_X1 U1361 ( .A1(n28), .A2(\REGISTERS[7][0] ), .B1(n27), .B2(
        \REGISTERS[6][0] ), .ZN(n1768) );
  OAI221_X1 U1362 ( .B1(n1829), .B2(n22), .C1(n1797), .C2(n19), .A(n1770), 
        .ZN(n1762) );
  AOI22_X1 U1363 ( .A1(n16), .A2(\REGISTERS[11][0] ), .B1(n15), .B2(
        \REGISTERS[10][0] ), .ZN(n1770) );
  OAI221_X1 U1364 ( .B1(n1956), .B2(n91), .C1(n1924), .C2(n88), .A(n1729), 
        .ZN(n1728) );
  AOI22_X1 U1365 ( .A1(n85), .A2(\REGISTERS[19][1] ), .B1(n84), .B2(
        \REGISTERS[18][1] ), .ZN(n1729) );
  OAI221_X1 U1366 ( .B1(n2020), .B2(n79), .C1(n1988), .C2(n76), .A(n1730), 
        .ZN(n1727) );
  AOI22_X1 U1367 ( .A1(n73), .A2(\REGISTERS[23][1] ), .B1(n72), .B2(
        \REGISTERS[22][1] ), .ZN(n1730) );
  OAI221_X1 U1368 ( .B1(n2084), .B2(n67), .C1(n2052), .C2(n64), .A(n1731), 
        .ZN(n1726) );
  AOI22_X1 U1369 ( .A1(n61), .A2(\REGISTERS[27][1] ), .B1(n60), .B2(
        \REGISTERS[26][1] ), .ZN(n1731) );
  OAI221_X1 U1370 ( .B1(n2148), .B2(n55), .C1(n2116), .C2(n52), .A(n1732), 
        .ZN(n1725) );
  AOI22_X1 U1371 ( .A1(n49), .A2(\REGISTERS[29][1] ), .B1(n48), .B2(
        \REGISTERS[28][1] ), .ZN(n1732) );
  OAI221_X1 U1372 ( .B1(n506), .B2(n34), .C1(n474), .C2(n31), .A(n1738), .ZN(
        n1735) );
  AOI22_X1 U1373 ( .A1(n28), .A2(\REGISTERS[7][1] ), .B1(n27), .B2(
        \REGISTERS[6][1] ), .ZN(n1738) );
  OAI221_X1 U1374 ( .B1(n1828), .B2(n22), .C1(n1796), .C2(n19), .A(n1739), 
        .ZN(n1734) );
  AOI22_X1 U1375 ( .A1(n16), .A2(\REGISTERS[11][1] ), .B1(n15), .B2(
        \REGISTERS[10][1] ), .ZN(n1739) );
  OAI221_X1 U1376 ( .B1(n1955), .B2(n91), .C1(n1923), .C2(n88), .A(n1711), 
        .ZN(n1710) );
  AOI22_X1 U1377 ( .A1(n85), .A2(\REGISTERS[19][2] ), .B1(n84), .B2(
        \REGISTERS[18][2] ), .ZN(n1711) );
  OAI221_X1 U1378 ( .B1(n2019), .B2(n79), .C1(n1987), .C2(n76), .A(n1712), 
        .ZN(n1709) );
  AOI22_X1 U1379 ( .A1(n73), .A2(\REGISTERS[23][2] ), .B1(n72), .B2(
        \REGISTERS[22][2] ), .ZN(n1712) );
  OAI221_X1 U1380 ( .B1(n2083), .B2(n67), .C1(n2051), .C2(n64), .A(n1713), 
        .ZN(n1708) );
  AOI22_X1 U1381 ( .A1(n61), .A2(\REGISTERS[27][2] ), .B1(n60), .B2(
        \REGISTERS[26][2] ), .ZN(n1713) );
  OAI221_X1 U1382 ( .B1(n2147), .B2(n55), .C1(n2115), .C2(n52), .A(n1714), 
        .ZN(n1707) );
  AOI22_X1 U1383 ( .A1(n49), .A2(\REGISTERS[29][2] ), .B1(n48), .B2(
        \REGISTERS[28][2] ), .ZN(n1714) );
  OAI221_X1 U1384 ( .B1(n505), .B2(n34), .C1(n473), .C2(n31), .A(n1720), .ZN(
        n1717) );
  AOI22_X1 U1385 ( .A1(n28), .A2(\REGISTERS[7][2] ), .B1(n27), .B2(
        \REGISTERS[6][2] ), .ZN(n1720) );
  OAI221_X1 U1386 ( .B1(n1827), .B2(n22), .C1(n1795), .C2(n19), .A(n1721), 
        .ZN(n1716) );
  AOI22_X1 U1387 ( .A1(n16), .A2(\REGISTERS[11][2] ), .B1(n15), .B2(
        \REGISTERS[10][2] ), .ZN(n1721) );
  OAI221_X1 U1388 ( .B1(n1954), .B2(n91), .C1(n1922), .C2(n88), .A(n1693), 
        .ZN(n1692) );
  AOI22_X1 U1389 ( .A1(n85), .A2(\REGISTERS[19][3] ), .B1(n84), .B2(
        \REGISTERS[18][3] ), .ZN(n1693) );
  OAI221_X1 U1390 ( .B1(n2018), .B2(n79), .C1(n1986), .C2(n76), .A(n1694), 
        .ZN(n1691) );
  AOI22_X1 U1391 ( .A1(n73), .A2(\REGISTERS[23][3] ), .B1(n72), .B2(
        \REGISTERS[22][3] ), .ZN(n1694) );
  OAI221_X1 U1392 ( .B1(n2082), .B2(n67), .C1(n2050), .C2(n64), .A(n1695), 
        .ZN(n1690) );
  AOI22_X1 U1393 ( .A1(n61), .A2(\REGISTERS[27][3] ), .B1(n60), .B2(
        \REGISTERS[26][3] ), .ZN(n1695) );
  OAI221_X1 U1394 ( .B1(n2146), .B2(n55), .C1(n2114), .C2(n52), .A(n1696), 
        .ZN(n1689) );
  AOI22_X1 U1395 ( .A1(n49), .A2(\REGISTERS[29][3] ), .B1(n48), .B2(
        \REGISTERS[28][3] ), .ZN(n1696) );
  OAI221_X1 U1396 ( .B1(n504), .B2(n34), .C1(n472), .C2(n31), .A(n1702), .ZN(
        n1699) );
  AOI22_X1 U1397 ( .A1(n28), .A2(\REGISTERS[7][3] ), .B1(n27), .B2(
        \REGISTERS[6][3] ), .ZN(n1702) );
  OAI221_X1 U1398 ( .B1(n1826), .B2(n22), .C1(n1794), .C2(n19), .A(n1703), 
        .ZN(n1698) );
  AOI22_X1 U1399 ( .A1(n16), .A2(\REGISTERS[11][3] ), .B1(n15), .B2(
        \REGISTERS[10][3] ), .ZN(n1703) );
  OAI221_X1 U1400 ( .B1(n1953), .B2(n91), .C1(n1921), .C2(n88), .A(n1675), 
        .ZN(n1674) );
  AOI22_X1 U1401 ( .A1(n85), .A2(\REGISTERS[19][4] ), .B1(n84), .B2(
        \REGISTERS[18][4] ), .ZN(n1675) );
  OAI221_X1 U1402 ( .B1(n2017), .B2(n79), .C1(n1985), .C2(n76), .A(n1676), 
        .ZN(n1673) );
  AOI22_X1 U1403 ( .A1(n73), .A2(\REGISTERS[23][4] ), .B1(n72), .B2(
        \REGISTERS[22][4] ), .ZN(n1676) );
  OAI221_X1 U1404 ( .B1(n2081), .B2(n67), .C1(n2049), .C2(n64), .A(n1677), 
        .ZN(n1672) );
  AOI22_X1 U1405 ( .A1(n61), .A2(\REGISTERS[27][4] ), .B1(n60), .B2(
        \REGISTERS[26][4] ), .ZN(n1677) );
  OAI221_X1 U1406 ( .B1(n2145), .B2(n55), .C1(n2113), .C2(n52), .A(n1678), 
        .ZN(n1671) );
  AOI22_X1 U1407 ( .A1(n49), .A2(\REGISTERS[29][4] ), .B1(n48), .B2(
        \REGISTERS[28][4] ), .ZN(n1678) );
  OAI221_X1 U1408 ( .B1(n503), .B2(n34), .C1(n471), .C2(n31), .A(n1684), .ZN(
        n1681) );
  AOI22_X1 U1409 ( .A1(n28), .A2(\REGISTERS[7][4] ), .B1(n27), .B2(
        \REGISTERS[6][4] ), .ZN(n1684) );
  OAI221_X1 U1410 ( .B1(n1825), .B2(n22), .C1(n1793), .C2(n19), .A(n1685), 
        .ZN(n1680) );
  AOI22_X1 U1411 ( .A1(n16), .A2(\REGISTERS[11][4] ), .B1(n15), .B2(
        \REGISTERS[10][4] ), .ZN(n1685) );
  OAI221_X1 U1412 ( .B1(n1952), .B2(n91), .C1(n1920), .C2(n88), .A(n1657), 
        .ZN(n1656) );
  AOI22_X1 U1413 ( .A1(n85), .A2(\REGISTERS[19][5] ), .B1(n84), .B2(
        \REGISTERS[18][5] ), .ZN(n1657) );
  OAI221_X1 U1414 ( .B1(n2016), .B2(n79), .C1(n1984), .C2(n76), .A(n1658), 
        .ZN(n1655) );
  AOI22_X1 U1415 ( .A1(n73), .A2(\REGISTERS[23][5] ), .B1(n72), .B2(
        \REGISTERS[22][5] ), .ZN(n1658) );
  OAI221_X1 U1416 ( .B1(n2080), .B2(n67), .C1(n2048), .C2(n64), .A(n1659), 
        .ZN(n1654) );
  AOI22_X1 U1417 ( .A1(n61), .A2(\REGISTERS[27][5] ), .B1(n60), .B2(
        \REGISTERS[26][5] ), .ZN(n1659) );
  OAI221_X1 U1418 ( .B1(n2144), .B2(n55), .C1(n2112), .C2(n52), .A(n1660), 
        .ZN(n1653) );
  AOI22_X1 U1419 ( .A1(n49), .A2(\REGISTERS[29][5] ), .B1(n48), .B2(
        \REGISTERS[28][5] ), .ZN(n1660) );
  OAI221_X1 U1420 ( .B1(n502), .B2(n34), .C1(n470), .C2(n31), .A(n1666), .ZN(
        n1663) );
  AOI22_X1 U1421 ( .A1(n28), .A2(\REGISTERS[7][5] ), .B1(n27), .B2(
        \REGISTERS[6][5] ), .ZN(n1666) );
  OAI221_X1 U1422 ( .B1(n1824), .B2(n22), .C1(n1792), .C2(n19), .A(n1667), 
        .ZN(n1662) );
  AOI22_X1 U1423 ( .A1(n16), .A2(\REGISTERS[11][5] ), .B1(n15), .B2(
        \REGISTERS[10][5] ), .ZN(n1667) );
  OAI221_X1 U1424 ( .B1(n1951), .B2(n91), .C1(n1919), .C2(n88), .A(n1639), 
        .ZN(n1638) );
  AOI22_X1 U1425 ( .A1(n85), .A2(\REGISTERS[19][6] ), .B1(n84), .B2(
        \REGISTERS[18][6] ), .ZN(n1639) );
  OAI221_X1 U1426 ( .B1(n2015), .B2(n79), .C1(n1983), .C2(n76), .A(n1640), 
        .ZN(n1637) );
  AOI22_X1 U1427 ( .A1(n73), .A2(\REGISTERS[23][6] ), .B1(n72), .B2(
        \REGISTERS[22][6] ), .ZN(n1640) );
  OAI221_X1 U1428 ( .B1(n2079), .B2(n67), .C1(n2047), .C2(n64), .A(n1641), 
        .ZN(n1636) );
  AOI22_X1 U1429 ( .A1(n61), .A2(\REGISTERS[27][6] ), .B1(n60), .B2(
        \REGISTERS[26][6] ), .ZN(n1641) );
  OAI221_X1 U1430 ( .B1(n2143), .B2(n55), .C1(n2111), .C2(n52), .A(n1642), 
        .ZN(n1635) );
  AOI22_X1 U1431 ( .A1(n49), .A2(\REGISTERS[29][6] ), .B1(n48), .B2(
        \REGISTERS[28][6] ), .ZN(n1642) );
  OAI221_X1 U1432 ( .B1(n501), .B2(n34), .C1(n469), .C2(n31), .A(n1648), .ZN(
        n1645) );
  AOI22_X1 U1433 ( .A1(n28), .A2(\REGISTERS[7][6] ), .B1(n27), .B2(
        \REGISTERS[6][6] ), .ZN(n1648) );
  OAI221_X1 U1434 ( .B1(n1823), .B2(n22), .C1(n1791), .C2(n19), .A(n1649), 
        .ZN(n1644) );
  AOI22_X1 U1435 ( .A1(n16), .A2(\REGISTERS[11][6] ), .B1(n15), .B2(
        \REGISTERS[10][6] ), .ZN(n1649) );
  OAI221_X1 U1436 ( .B1(n1950), .B2(n91), .C1(n1918), .C2(n88), .A(n1621), 
        .ZN(n1620) );
  AOI22_X1 U1437 ( .A1(n85), .A2(\REGISTERS[19][7] ), .B1(n84), .B2(
        \REGISTERS[18][7] ), .ZN(n1621) );
  OAI221_X1 U1438 ( .B1(n2014), .B2(n79), .C1(n1982), .C2(n76), .A(n1622), 
        .ZN(n1619) );
  AOI22_X1 U1439 ( .A1(n73), .A2(\REGISTERS[23][7] ), .B1(n72), .B2(
        \REGISTERS[22][7] ), .ZN(n1622) );
  OAI221_X1 U1440 ( .B1(n2078), .B2(n67), .C1(n2046), .C2(n64), .A(n1623), 
        .ZN(n1618) );
  AOI22_X1 U1441 ( .A1(n61), .A2(\REGISTERS[27][7] ), .B1(n60), .B2(
        \REGISTERS[26][7] ), .ZN(n1623) );
  OAI221_X1 U1442 ( .B1(n2142), .B2(n55), .C1(n2110), .C2(n52), .A(n1624), 
        .ZN(n1617) );
  AOI22_X1 U1443 ( .A1(n49), .A2(\REGISTERS[29][7] ), .B1(n48), .B2(
        \REGISTERS[28][7] ), .ZN(n1624) );
  OAI221_X1 U1444 ( .B1(n500), .B2(n34), .C1(n468), .C2(n31), .A(n1630), .ZN(
        n1627) );
  AOI22_X1 U1445 ( .A1(n28), .A2(\REGISTERS[7][7] ), .B1(n27), .B2(
        \REGISTERS[6][7] ), .ZN(n1630) );
  OAI221_X1 U1446 ( .B1(n1822), .B2(n22), .C1(n1790), .C2(n19), .A(n1631), 
        .ZN(n1626) );
  AOI22_X1 U1447 ( .A1(n16), .A2(\REGISTERS[11][7] ), .B1(n15), .B2(
        \REGISTERS[10][7] ), .ZN(n1631) );
  OAI221_X1 U1448 ( .B1(n1949), .B2(n91), .C1(n1917), .C2(n88), .A(n1603), 
        .ZN(n1602) );
  AOI22_X1 U1449 ( .A1(n85), .A2(\REGISTERS[19][8] ), .B1(n83), .B2(
        \REGISTERS[18][8] ), .ZN(n1603) );
  OAI221_X1 U1450 ( .B1(n2013), .B2(n79), .C1(n1981), .C2(n76), .A(n1604), 
        .ZN(n1601) );
  AOI22_X1 U1451 ( .A1(n73), .A2(\REGISTERS[23][8] ), .B1(n71), .B2(
        \REGISTERS[22][8] ), .ZN(n1604) );
  OAI221_X1 U1452 ( .B1(n2077), .B2(n67), .C1(n2045), .C2(n64), .A(n1605), 
        .ZN(n1600) );
  AOI22_X1 U1453 ( .A1(n61), .A2(\REGISTERS[27][8] ), .B1(n59), .B2(
        \REGISTERS[26][8] ), .ZN(n1605) );
  OAI221_X1 U1454 ( .B1(n2141), .B2(n55), .C1(n2109), .C2(n52), .A(n1606), 
        .ZN(n1599) );
  AOI22_X1 U1455 ( .A1(n49), .A2(\REGISTERS[29][8] ), .B1(n47), .B2(
        \REGISTERS[28][8] ), .ZN(n1606) );
  OAI221_X1 U1456 ( .B1(n1821), .B2(n22), .C1(n1789), .C2(n19), .A(n1613), 
        .ZN(n1608) );
  AOI22_X1 U1457 ( .A1(n16), .A2(\REGISTERS[11][8] ), .B1(n14), .B2(
        \REGISTERS[10][8] ), .ZN(n1613) );
  OAI221_X1 U1458 ( .B1(n1948), .B2(n91), .C1(n1916), .C2(n88), .A(n1585), 
        .ZN(n1584) );
  AOI22_X1 U1459 ( .A1(n85), .A2(\REGISTERS[19][9] ), .B1(n83), .B2(
        \REGISTERS[18][9] ), .ZN(n1585) );
  OAI221_X1 U1460 ( .B1(n2012), .B2(n79), .C1(n1980), .C2(n76), .A(n1586), 
        .ZN(n1583) );
  AOI22_X1 U1461 ( .A1(n73), .A2(\REGISTERS[23][9] ), .B1(n71), .B2(
        \REGISTERS[22][9] ), .ZN(n1586) );
  OAI221_X1 U1462 ( .B1(n2076), .B2(n67), .C1(n2044), .C2(n64), .A(n1587), 
        .ZN(n1582) );
  AOI22_X1 U1463 ( .A1(n61), .A2(\REGISTERS[27][9] ), .B1(n59), .B2(
        \REGISTERS[26][9] ), .ZN(n1587) );
  OAI221_X1 U1464 ( .B1(n2140), .B2(n55), .C1(n2108), .C2(n52), .A(n1588), 
        .ZN(n1581) );
  AOI22_X1 U1465 ( .A1(n49), .A2(\REGISTERS[29][9] ), .B1(n47), .B2(
        \REGISTERS[28][9] ), .ZN(n1588) );
  OAI221_X1 U1466 ( .B1(n1820), .B2(n22), .C1(n1788), .C2(n19), .A(n1595), 
        .ZN(n1590) );
  AOI22_X1 U1467 ( .A1(n16), .A2(\REGISTERS[11][9] ), .B1(n14), .B2(
        \REGISTERS[10][9] ), .ZN(n1595) );
  OAI221_X1 U1468 ( .B1(n1947), .B2(n91), .C1(n1915), .C2(n88), .A(n1567), 
        .ZN(n1566) );
  AOI22_X1 U1469 ( .A1(n85), .A2(\REGISTERS[19][10] ), .B1(n83), .B2(
        \REGISTERS[18][10] ), .ZN(n1567) );
  OAI221_X1 U1470 ( .B1(n2011), .B2(n79), .C1(n1979), .C2(n76), .A(n1568), 
        .ZN(n1565) );
  AOI22_X1 U1471 ( .A1(n73), .A2(\REGISTERS[23][10] ), .B1(n71), .B2(
        \REGISTERS[22][10] ), .ZN(n1568) );
  OAI221_X1 U1472 ( .B1(n2075), .B2(n67), .C1(n2043), .C2(n64), .A(n1569), 
        .ZN(n1564) );
  AOI22_X1 U1473 ( .A1(n61), .A2(\REGISTERS[27][10] ), .B1(n59), .B2(
        \REGISTERS[26][10] ), .ZN(n1569) );
  OAI221_X1 U1474 ( .B1(n2139), .B2(n55), .C1(n2107), .C2(n52), .A(n1570), 
        .ZN(n1563) );
  AOI22_X1 U1475 ( .A1(n49), .A2(\REGISTERS[29][10] ), .B1(n47), .B2(
        \REGISTERS[28][10] ), .ZN(n1570) );
  OAI221_X1 U1476 ( .B1(n1819), .B2(n22), .C1(n1787), .C2(n19), .A(n1577), 
        .ZN(n1572) );
  AOI22_X1 U1477 ( .A1(n16), .A2(\REGISTERS[11][10] ), .B1(n14), .B2(
        \REGISTERS[10][10] ), .ZN(n1577) );
  OAI221_X1 U1478 ( .B1(n1946), .B2(n91), .C1(n1914), .C2(n88), .A(n1549), 
        .ZN(n1548) );
  AOI22_X1 U1479 ( .A1(n85), .A2(\REGISTERS[19][11] ), .B1(n83), .B2(
        \REGISTERS[18][11] ), .ZN(n1549) );
  OAI221_X1 U1480 ( .B1(n2010), .B2(n79), .C1(n1978), .C2(n76), .A(n1550), 
        .ZN(n1547) );
  AOI22_X1 U1481 ( .A1(n73), .A2(\REGISTERS[23][11] ), .B1(n71), .B2(
        \REGISTERS[22][11] ), .ZN(n1550) );
  OAI221_X1 U1482 ( .B1(n2074), .B2(n67), .C1(n2042), .C2(n64), .A(n1551), 
        .ZN(n1546) );
  AOI22_X1 U1483 ( .A1(n61), .A2(\REGISTERS[27][11] ), .B1(n59), .B2(
        \REGISTERS[26][11] ), .ZN(n1551) );
  OAI221_X1 U1484 ( .B1(n2138), .B2(n55), .C1(n2106), .C2(n52), .A(n1552), 
        .ZN(n1545) );
  AOI22_X1 U1485 ( .A1(n49), .A2(\REGISTERS[29][11] ), .B1(n47), .B2(
        \REGISTERS[28][11] ), .ZN(n1552) );
  OAI221_X1 U1486 ( .B1(n1818), .B2(n22), .C1(n1182), .C2(n19), .A(n1559), 
        .ZN(n1554) );
  AOI22_X1 U1487 ( .A1(n16), .A2(\REGISTERS[11][11] ), .B1(n14), .B2(
        \REGISTERS[10][11] ), .ZN(n1559) );
  OAI221_X1 U1488 ( .B1(n1945), .B2(n92), .C1(n1913), .C2(n89), .A(n1531), 
        .ZN(n1530) );
  AOI22_X1 U1489 ( .A1(n86), .A2(\REGISTERS[19][12] ), .B1(n83), .B2(
        \REGISTERS[18][12] ), .ZN(n1531) );
  OAI221_X1 U1490 ( .B1(n2009), .B2(n80), .C1(n1977), .C2(n77), .A(n1532), 
        .ZN(n1529) );
  AOI22_X1 U1491 ( .A1(n74), .A2(\REGISTERS[23][12] ), .B1(n71), .B2(
        \REGISTERS[22][12] ), .ZN(n1532) );
  OAI221_X1 U1492 ( .B1(n2073), .B2(n68), .C1(n2041), .C2(n65), .A(n1533), 
        .ZN(n1528) );
  AOI22_X1 U1493 ( .A1(n62), .A2(\REGISTERS[27][12] ), .B1(n59), .B2(
        \REGISTERS[26][12] ), .ZN(n1533) );
  OAI221_X1 U1494 ( .B1(n2137), .B2(n56), .C1(n2105), .C2(n53), .A(n1534), 
        .ZN(n1527) );
  AOI22_X1 U1495 ( .A1(n50), .A2(\REGISTERS[29][12] ), .B1(n47), .B2(
        \REGISTERS[28][12] ), .ZN(n1534) );
  OAI221_X1 U1496 ( .B1(n1817), .B2(n23), .C1(n558), .C2(n20), .A(n1541), .ZN(
        n1536) );
  AOI22_X1 U1497 ( .A1(n17), .A2(\REGISTERS[11][12] ), .B1(n14), .B2(
        \REGISTERS[10][12] ), .ZN(n1541) );
  OAI221_X1 U1498 ( .B1(n1944), .B2(n92), .C1(n1912), .C2(n89), .A(n1513), 
        .ZN(n1512) );
  AOI22_X1 U1499 ( .A1(n86), .A2(\REGISTERS[19][13] ), .B1(n83), .B2(
        \REGISTERS[18][13] ), .ZN(n1513) );
  OAI221_X1 U1500 ( .B1(n2008), .B2(n80), .C1(n1976), .C2(n77), .A(n1514), 
        .ZN(n1511) );
  AOI22_X1 U1501 ( .A1(n74), .A2(\REGISTERS[23][13] ), .B1(n71), .B2(
        \REGISTERS[22][13] ), .ZN(n1514) );
  OAI221_X1 U1502 ( .B1(n2072), .B2(n68), .C1(n2040), .C2(n65), .A(n1515), 
        .ZN(n1510) );
  AOI22_X1 U1503 ( .A1(n62), .A2(\REGISTERS[27][13] ), .B1(n59), .B2(
        \REGISTERS[26][13] ), .ZN(n1515) );
  OAI221_X1 U1504 ( .B1(n2136), .B2(n56), .C1(n2104), .C2(n53), .A(n1516), 
        .ZN(n1509) );
  AOI22_X1 U1505 ( .A1(n50), .A2(\REGISTERS[29][13] ), .B1(n47), .B2(
        \REGISTERS[28][13] ), .ZN(n1516) );
  OAI221_X1 U1506 ( .B1(n1816), .B2(n23), .C1(n526), .C2(n20), .A(n1523), .ZN(
        n1518) );
  AOI22_X1 U1507 ( .A1(n17), .A2(\REGISTERS[11][13] ), .B1(n14), .B2(
        \REGISTERS[10][13] ), .ZN(n1523) );
  OAI221_X1 U1508 ( .B1(n1943), .B2(n92), .C1(n1911), .C2(n89), .A(n1495), 
        .ZN(n1494) );
  AOI22_X1 U1509 ( .A1(n86), .A2(\REGISTERS[19][14] ), .B1(n83), .B2(
        \REGISTERS[18][14] ), .ZN(n1495) );
  OAI221_X1 U1510 ( .B1(n2007), .B2(n80), .C1(n1975), .C2(n77), .A(n1496), 
        .ZN(n1493) );
  AOI22_X1 U1511 ( .A1(n74), .A2(\REGISTERS[23][14] ), .B1(n71), .B2(
        \REGISTERS[22][14] ), .ZN(n1496) );
  OAI221_X1 U1512 ( .B1(n2071), .B2(n68), .C1(n2039), .C2(n65), .A(n1497), 
        .ZN(n1492) );
  AOI22_X1 U1513 ( .A1(n62), .A2(\REGISTERS[27][14] ), .B1(n59), .B2(
        \REGISTERS[26][14] ), .ZN(n1497) );
  OAI221_X1 U1514 ( .B1(n2135), .B2(n56), .C1(n2103), .C2(n53), .A(n1498), 
        .ZN(n1491) );
  AOI22_X1 U1515 ( .A1(n50), .A2(\REGISTERS[29][14] ), .B1(n47), .B2(
        \REGISTERS[28][14] ), .ZN(n1498) );
  OAI221_X1 U1516 ( .B1(n1815), .B2(n23), .C1(n525), .C2(n20), .A(n1505), .ZN(
        n1500) );
  AOI22_X1 U1517 ( .A1(n17), .A2(\REGISTERS[11][14] ), .B1(n14), .B2(
        \REGISTERS[10][14] ), .ZN(n1505) );
  OAI221_X1 U1518 ( .B1(n1942), .B2(n92), .C1(n1910), .C2(n89), .A(n1477), 
        .ZN(n1476) );
  AOI22_X1 U1519 ( .A1(n86), .A2(\REGISTERS[19][15] ), .B1(n83), .B2(
        \REGISTERS[18][15] ), .ZN(n1477) );
  OAI221_X1 U1520 ( .B1(n2006), .B2(n80), .C1(n1974), .C2(n77), .A(n1478), 
        .ZN(n1475) );
  AOI22_X1 U1521 ( .A1(n74), .A2(\REGISTERS[23][15] ), .B1(n71), .B2(
        \REGISTERS[22][15] ), .ZN(n1478) );
  OAI221_X1 U1522 ( .B1(n2070), .B2(n68), .C1(n2038), .C2(n65), .A(n1479), 
        .ZN(n1474) );
  AOI22_X1 U1523 ( .A1(n62), .A2(\REGISTERS[27][15] ), .B1(n59), .B2(
        \REGISTERS[26][15] ), .ZN(n1479) );
  OAI221_X1 U1524 ( .B1(n2134), .B2(n56), .C1(n2102), .C2(n53), .A(n1480), 
        .ZN(n1473) );
  AOI22_X1 U1525 ( .A1(n50), .A2(\REGISTERS[29][15] ), .B1(n47), .B2(
        \REGISTERS[28][15] ), .ZN(n1480) );
  OAI221_X1 U1526 ( .B1(n1814), .B2(n23), .C1(n524), .C2(n20), .A(n1487), .ZN(
        n1482) );
  AOI22_X1 U1527 ( .A1(n17), .A2(\REGISTERS[11][15] ), .B1(n14), .B2(
        \REGISTERS[10][15] ), .ZN(n1487) );
  OAI221_X1 U1528 ( .B1(n1941), .B2(n92), .C1(n1909), .C2(n89), .A(n1459), 
        .ZN(n1458) );
  AOI22_X1 U1529 ( .A1(n86), .A2(\REGISTERS[19][16] ), .B1(n83), .B2(
        \REGISTERS[18][16] ), .ZN(n1459) );
  OAI221_X1 U1530 ( .B1(n2005), .B2(n80), .C1(n1973), .C2(n77), .A(n1460), 
        .ZN(n1457) );
  AOI22_X1 U1531 ( .A1(n74), .A2(\REGISTERS[23][16] ), .B1(n71), .B2(
        \REGISTERS[22][16] ), .ZN(n1460) );
  OAI221_X1 U1532 ( .B1(n2069), .B2(n68), .C1(n2037), .C2(n65), .A(n1461), 
        .ZN(n1456) );
  AOI22_X1 U1533 ( .A1(n62), .A2(\REGISTERS[27][16] ), .B1(n59), .B2(
        \REGISTERS[26][16] ), .ZN(n1461) );
  OAI221_X1 U1534 ( .B1(n2133), .B2(n56), .C1(n2101), .C2(n53), .A(n1462), 
        .ZN(n1455) );
  AOI22_X1 U1535 ( .A1(n50), .A2(\REGISTERS[29][16] ), .B1(n47), .B2(
        \REGISTERS[28][16] ), .ZN(n1462) );
  OAI221_X1 U1536 ( .B1(n1813), .B2(n23), .C1(n523), .C2(n20), .A(n1469), .ZN(
        n1464) );
  AOI22_X1 U1537 ( .A1(n17), .A2(\REGISTERS[11][16] ), .B1(n14), .B2(
        \REGISTERS[10][16] ), .ZN(n1469) );
  OAI221_X1 U1538 ( .B1(n1940), .B2(n92), .C1(n1908), .C2(n89), .A(n1441), 
        .ZN(n1440) );
  AOI22_X1 U1539 ( .A1(n86), .A2(\REGISTERS[19][17] ), .B1(n83), .B2(
        \REGISTERS[18][17] ), .ZN(n1441) );
  OAI221_X1 U1540 ( .B1(n2004), .B2(n80), .C1(n1972), .C2(n77), .A(n1442), 
        .ZN(n1439) );
  AOI22_X1 U1541 ( .A1(n74), .A2(\REGISTERS[23][17] ), .B1(n71), .B2(
        \REGISTERS[22][17] ), .ZN(n1442) );
  OAI221_X1 U1542 ( .B1(n2068), .B2(n68), .C1(n2036), .C2(n65), .A(n1443), 
        .ZN(n1438) );
  AOI22_X1 U1543 ( .A1(n62), .A2(\REGISTERS[27][17] ), .B1(n59), .B2(
        \REGISTERS[26][17] ), .ZN(n1443) );
  OAI221_X1 U1544 ( .B1(n2132), .B2(n56), .C1(n2100), .C2(n53), .A(n1444), 
        .ZN(n1437) );
  AOI22_X1 U1545 ( .A1(n50), .A2(\REGISTERS[29][17] ), .B1(n47), .B2(
        \REGISTERS[28][17] ), .ZN(n1444) );
  OAI221_X1 U1546 ( .B1(n1812), .B2(n23), .C1(n522), .C2(n20), .A(n1451), .ZN(
        n1446) );
  AOI22_X1 U1547 ( .A1(n17), .A2(\REGISTERS[11][17] ), .B1(n14), .B2(
        \REGISTERS[10][17] ), .ZN(n1451) );
  OAI221_X1 U1548 ( .B1(n1939), .B2(n92), .C1(n1907), .C2(n89), .A(n1423), 
        .ZN(n1422) );
  AOI22_X1 U1549 ( .A1(n86), .A2(\REGISTERS[19][18] ), .B1(n83), .B2(
        \REGISTERS[18][18] ), .ZN(n1423) );
  OAI221_X1 U1550 ( .B1(n2003), .B2(n80), .C1(n1971), .C2(n77), .A(n1424), 
        .ZN(n1421) );
  AOI22_X1 U1551 ( .A1(n74), .A2(\REGISTERS[23][18] ), .B1(n71), .B2(
        \REGISTERS[22][18] ), .ZN(n1424) );
  OAI221_X1 U1552 ( .B1(n2067), .B2(n68), .C1(n2035), .C2(n65), .A(n1425), 
        .ZN(n1420) );
  AOI22_X1 U1553 ( .A1(n62), .A2(\REGISTERS[27][18] ), .B1(n59), .B2(
        \REGISTERS[26][18] ), .ZN(n1425) );
  OAI221_X1 U1554 ( .B1(n2131), .B2(n56), .C1(n2099), .C2(n53), .A(n1426), 
        .ZN(n1419) );
  AOI22_X1 U1555 ( .A1(n50), .A2(\REGISTERS[29][18] ), .B1(n47), .B2(
        \REGISTERS[28][18] ), .ZN(n1426) );
  OAI221_X1 U1556 ( .B1(n1811), .B2(n23), .C1(n521), .C2(n20), .A(n1433), .ZN(
        n1428) );
  AOI22_X1 U1557 ( .A1(n17), .A2(\REGISTERS[11][18] ), .B1(n14), .B2(
        \REGISTERS[10][18] ), .ZN(n1433) );
  OAI221_X1 U1558 ( .B1(n1938), .B2(n92), .C1(n1906), .C2(n89), .A(n1405), 
        .ZN(n1404) );
  AOI22_X1 U1559 ( .A1(n86), .A2(\REGISTERS[19][19] ), .B1(n83), .B2(
        \REGISTERS[18][19] ), .ZN(n1405) );
  OAI221_X1 U1560 ( .B1(n2002), .B2(n80), .C1(n1970), .C2(n77), .A(n1406), 
        .ZN(n1403) );
  AOI22_X1 U1561 ( .A1(n74), .A2(\REGISTERS[23][19] ), .B1(n71), .B2(
        \REGISTERS[22][19] ), .ZN(n1406) );
  OAI221_X1 U1562 ( .B1(n2066), .B2(n68), .C1(n2034), .C2(n65), .A(n1407), 
        .ZN(n1402) );
  AOI22_X1 U1563 ( .A1(n62), .A2(\REGISTERS[27][19] ), .B1(n59), .B2(
        \REGISTERS[26][19] ), .ZN(n1407) );
  OAI221_X1 U1564 ( .B1(n2130), .B2(n56), .C1(n2098), .C2(n53), .A(n1408), 
        .ZN(n1401) );
  AOI22_X1 U1565 ( .A1(n50), .A2(\REGISTERS[29][19] ), .B1(n47), .B2(
        \REGISTERS[28][19] ), .ZN(n1408) );
  OAI221_X1 U1566 ( .B1(n1810), .B2(n23), .C1(n520), .C2(n20), .A(n1415), .ZN(
        n1410) );
  AOI22_X1 U1567 ( .A1(n17), .A2(\REGISTERS[11][19] ), .B1(n14), .B2(
        \REGISTERS[10][19] ), .ZN(n1415) );
  OAI221_X1 U1568 ( .B1(n1937), .B2(n92), .C1(n1905), .C2(n89), .A(n1387), 
        .ZN(n1386) );
  AOI22_X1 U1569 ( .A1(n86), .A2(\REGISTERS[19][20] ), .B1(n82), .B2(
        \REGISTERS[18][20] ), .ZN(n1387) );
  OAI221_X1 U1570 ( .B1(n2001), .B2(n80), .C1(n1969), .C2(n77), .A(n1388), 
        .ZN(n1385) );
  AOI22_X1 U1571 ( .A1(n74), .A2(\REGISTERS[23][20] ), .B1(n70), .B2(
        \REGISTERS[22][20] ), .ZN(n1388) );
  OAI221_X1 U1572 ( .B1(n2065), .B2(n68), .C1(n2033), .C2(n65), .A(n1389), 
        .ZN(n1384) );
  AOI22_X1 U1573 ( .A1(n62), .A2(\REGISTERS[27][20] ), .B1(n58), .B2(
        \REGISTERS[26][20] ), .ZN(n1389) );
  OAI221_X1 U1574 ( .B1(n2129), .B2(n56), .C1(n2097), .C2(n53), .A(n1390), 
        .ZN(n1383) );
  AOI22_X1 U1575 ( .A1(n50), .A2(\REGISTERS[29][20] ), .B1(n46), .B2(
        \REGISTERS[28][20] ), .ZN(n1390) );
  OAI221_X1 U1576 ( .B1(n1809), .B2(n23), .C1(n519), .C2(n20), .A(n1397), .ZN(
        n1392) );
  AOI22_X1 U1577 ( .A1(n17), .A2(\REGISTERS[11][20] ), .B1(n13), .B2(
        \REGISTERS[10][20] ), .ZN(n1397) );
  OAI221_X1 U1578 ( .B1(n1936), .B2(n92), .C1(n1904), .C2(n89), .A(n1369), 
        .ZN(n1368) );
  AOI22_X1 U1579 ( .A1(n86), .A2(\REGISTERS[19][21] ), .B1(n82), .B2(
        \REGISTERS[18][21] ), .ZN(n1369) );
  OAI221_X1 U1580 ( .B1(n2000), .B2(n80), .C1(n1968), .C2(n77), .A(n1370), 
        .ZN(n1367) );
  AOI22_X1 U1581 ( .A1(n74), .A2(\REGISTERS[23][21] ), .B1(n70), .B2(
        \REGISTERS[22][21] ), .ZN(n1370) );
  OAI221_X1 U1582 ( .B1(n2064), .B2(n68), .C1(n2032), .C2(n65), .A(n1371), 
        .ZN(n1366) );
  AOI22_X1 U1583 ( .A1(n62), .A2(\REGISTERS[27][21] ), .B1(n58), .B2(
        \REGISTERS[26][21] ), .ZN(n1371) );
  OAI221_X1 U1584 ( .B1(n2128), .B2(n56), .C1(n2096), .C2(n53), .A(n1372), 
        .ZN(n1365) );
  AOI22_X1 U1585 ( .A1(n50), .A2(\REGISTERS[29][21] ), .B1(n46), .B2(
        \REGISTERS[28][21] ), .ZN(n1372) );
  OAI221_X1 U1586 ( .B1(n1808), .B2(n23), .C1(n518), .C2(n20), .A(n1379), .ZN(
        n1374) );
  AOI22_X1 U1587 ( .A1(n17), .A2(\REGISTERS[11][21] ), .B1(n13), .B2(
        \REGISTERS[10][21] ), .ZN(n1379) );
  OAI221_X1 U1588 ( .B1(n1935), .B2(n92), .C1(n1903), .C2(n89), .A(n1351), 
        .ZN(n1350) );
  AOI22_X1 U1589 ( .A1(n86), .A2(\REGISTERS[19][22] ), .B1(n82), .B2(
        \REGISTERS[18][22] ), .ZN(n1351) );
  OAI221_X1 U1590 ( .B1(n1999), .B2(n80), .C1(n1967), .C2(n77), .A(n1352), 
        .ZN(n1349) );
  AOI22_X1 U1591 ( .A1(n74), .A2(\REGISTERS[23][22] ), .B1(n70), .B2(
        \REGISTERS[22][22] ), .ZN(n1352) );
  OAI221_X1 U1592 ( .B1(n2063), .B2(n68), .C1(n2031), .C2(n65), .A(n1353), 
        .ZN(n1348) );
  AOI22_X1 U1593 ( .A1(n62), .A2(\REGISTERS[27][22] ), .B1(n58), .B2(
        \REGISTERS[26][22] ), .ZN(n1353) );
  OAI221_X1 U1594 ( .B1(n2127), .B2(n56), .C1(n2095), .C2(n53), .A(n1354), 
        .ZN(n1347) );
  AOI22_X1 U1595 ( .A1(n50), .A2(\REGISTERS[29][22] ), .B1(n46), .B2(
        \REGISTERS[28][22] ), .ZN(n1354) );
  OAI221_X1 U1596 ( .B1(n1807), .B2(n23), .C1(n517), .C2(n20), .A(n1361), .ZN(
        n1356) );
  AOI22_X1 U1597 ( .A1(n17), .A2(\REGISTERS[11][22] ), .B1(n13), .B2(
        \REGISTERS[10][22] ), .ZN(n1361) );
  OAI221_X1 U1598 ( .B1(n1934), .B2(n92), .C1(n1902), .C2(n89), .A(n1333), 
        .ZN(n1332) );
  AOI22_X1 U1599 ( .A1(n86), .A2(\REGISTERS[19][23] ), .B1(n82), .B2(
        \REGISTERS[18][23] ), .ZN(n1333) );
  OAI221_X1 U1600 ( .B1(n1998), .B2(n80), .C1(n1966), .C2(n77), .A(n1334), 
        .ZN(n1331) );
  AOI22_X1 U1601 ( .A1(n74), .A2(\REGISTERS[23][23] ), .B1(n70), .B2(
        \REGISTERS[22][23] ), .ZN(n1334) );
  OAI221_X1 U1602 ( .B1(n2062), .B2(n68), .C1(n2030), .C2(n65), .A(n1335), 
        .ZN(n1330) );
  AOI22_X1 U1603 ( .A1(n62), .A2(\REGISTERS[27][23] ), .B1(n58), .B2(
        \REGISTERS[26][23] ), .ZN(n1335) );
  OAI221_X1 U1604 ( .B1(n2126), .B2(n56), .C1(n2094), .C2(n53), .A(n1336), 
        .ZN(n1329) );
  AOI22_X1 U1605 ( .A1(n50), .A2(\REGISTERS[29][23] ), .B1(n46), .B2(
        \REGISTERS[28][23] ), .ZN(n1336) );
  OAI221_X1 U1606 ( .B1(n1806), .B2(n23), .C1(n516), .C2(n20), .A(n1343), .ZN(
        n1338) );
  AOI22_X1 U1607 ( .A1(n17), .A2(\REGISTERS[11][23] ), .B1(n13), .B2(
        \REGISTERS[10][23] ), .ZN(n1343) );
  OAI221_X1 U1608 ( .B1(n2061), .B2(n69), .C1(n2029), .C2(n66), .A(n1317), 
        .ZN(n1312) );
  AOI22_X1 U1609 ( .A1(n63), .A2(\REGISTERS[27][24] ), .B1(n58), .B2(
        \REGISTERS[26][24] ), .ZN(n1317) );
  OAI221_X1 U1610 ( .B1(n2125), .B2(n57), .C1(n2093), .C2(n54), .A(n1318), 
        .ZN(n1311) );
  AOI22_X1 U1611 ( .A1(n51), .A2(\REGISTERS[29][24] ), .B1(n46), .B2(
        \REGISTERS[28][24] ), .ZN(n1318) );
  OAI221_X1 U1612 ( .B1(n1805), .B2(n24), .C1(n515), .C2(n21), .A(n1325), .ZN(
        n1320) );
  AOI22_X1 U1613 ( .A1(n18), .A2(\REGISTERS[11][24] ), .B1(n13), .B2(
        \REGISTERS[10][24] ), .ZN(n1325) );
  OAI221_X1 U1614 ( .B1(n2060), .B2(n69), .C1(n2028), .C2(n66), .A(n1299), 
        .ZN(n1294) );
  AOI22_X1 U1615 ( .A1(n63), .A2(\REGISTERS[27][25] ), .B1(n58), .B2(
        \REGISTERS[26][25] ), .ZN(n1299) );
  OAI221_X1 U1616 ( .B1(n2124), .B2(n57), .C1(n2092), .C2(n54), .A(n1300), 
        .ZN(n1293) );
  AOI22_X1 U1617 ( .A1(n51), .A2(\REGISTERS[29][25] ), .B1(n46), .B2(
        \REGISTERS[28][25] ), .ZN(n1300) );
  OAI221_X1 U1618 ( .B1(n1804), .B2(n24), .C1(n514), .C2(n21), .A(n1307), .ZN(
        n1302) );
  AOI22_X1 U1619 ( .A1(n18), .A2(\REGISTERS[11][25] ), .B1(n13), .B2(
        \REGISTERS[10][25] ), .ZN(n1307) );
  OAI221_X1 U1620 ( .B1(n2059), .B2(n69), .C1(n2027), .C2(n66), .A(n1281), 
        .ZN(n1276) );
  AOI22_X1 U1621 ( .A1(n63), .A2(\REGISTERS[27][26] ), .B1(n58), .B2(
        \REGISTERS[26][26] ), .ZN(n1281) );
  OAI221_X1 U1622 ( .B1(n2123), .B2(n57), .C1(n2091), .C2(n54), .A(n1282), 
        .ZN(n1275) );
  AOI22_X1 U1623 ( .A1(n51), .A2(\REGISTERS[29][26] ), .B1(n46), .B2(
        \REGISTERS[28][26] ), .ZN(n1282) );
  OAI221_X1 U1624 ( .B1(n1803), .B2(n24), .C1(n513), .C2(n21), .A(n1289), .ZN(
        n1284) );
  AOI22_X1 U1625 ( .A1(n18), .A2(\REGISTERS[11][26] ), .B1(n13), .B2(
        \REGISTERS[10][26] ), .ZN(n1289) );
  OAI221_X1 U1626 ( .B1(n2058), .B2(n69), .C1(n2026), .C2(n66), .A(n1263), 
        .ZN(n1258) );
  AOI22_X1 U1627 ( .A1(n63), .A2(\REGISTERS[27][27] ), .B1(n58), .B2(
        \REGISTERS[26][27] ), .ZN(n1263) );
  OAI221_X1 U1628 ( .B1(n2122), .B2(n57), .C1(n2090), .C2(n54), .A(n1264), 
        .ZN(n1257) );
  AOI22_X1 U1629 ( .A1(n51), .A2(\REGISTERS[29][27] ), .B1(n46), .B2(
        \REGISTERS[28][27] ), .ZN(n1264) );
  OAI221_X1 U1630 ( .B1(n1802), .B2(n24), .C1(n512), .C2(n21), .A(n1271), .ZN(
        n1266) );
  AOI22_X1 U1631 ( .A1(n18), .A2(\REGISTERS[11][27] ), .B1(n13), .B2(
        \REGISTERS[10][27] ), .ZN(n1271) );
  OAI221_X1 U1632 ( .B1(n2057), .B2(n69), .C1(n2025), .C2(n66), .A(n1245), 
        .ZN(n1240) );
  AOI22_X1 U1633 ( .A1(n63), .A2(\REGISTERS[27][28] ), .B1(n58), .B2(
        \REGISTERS[26][28] ), .ZN(n1245) );
  OAI221_X1 U1634 ( .B1(n2121), .B2(n57), .C1(n2089), .C2(n54), .A(n1246), 
        .ZN(n1239) );
  AOI22_X1 U1635 ( .A1(n51), .A2(\REGISTERS[29][28] ), .B1(n46), .B2(
        \REGISTERS[28][28] ), .ZN(n1246) );
  OAI221_X1 U1636 ( .B1(n1801), .B2(n24), .C1(n511), .C2(n21), .A(n1253), .ZN(
        n1248) );
  AOI22_X1 U1637 ( .A1(n18), .A2(\REGISTERS[11][28] ), .B1(n13), .B2(
        \REGISTERS[10][28] ), .ZN(n1253) );
  OAI221_X1 U1638 ( .B1(n2056), .B2(n69), .C1(n2024), .C2(n66), .A(n1227), 
        .ZN(n1222) );
  AOI22_X1 U1639 ( .A1(n63), .A2(\REGISTERS[27][29] ), .B1(n58), .B2(
        \REGISTERS[26][29] ), .ZN(n1227) );
  OAI221_X1 U1640 ( .B1(n2120), .B2(n57), .C1(n2088), .C2(n54), .A(n1228), 
        .ZN(n1221) );
  AOI22_X1 U1641 ( .A1(n51), .A2(\REGISTERS[29][29] ), .B1(n46), .B2(
        \REGISTERS[28][29] ), .ZN(n1228) );
  OAI221_X1 U1642 ( .B1(n1800), .B2(n24), .C1(n510), .C2(n21), .A(n1235), .ZN(
        n1230) );
  AOI22_X1 U1643 ( .A1(n18), .A2(\REGISTERS[11][29] ), .B1(n13), .B2(
        \REGISTERS[10][29] ), .ZN(n1235) );
  OAI221_X1 U1644 ( .B1(n2055), .B2(n69), .C1(n2023), .C2(n66), .A(n1209), 
        .ZN(n1204) );
  AOI22_X1 U1645 ( .A1(n63), .A2(\REGISTERS[27][30] ), .B1(n58), .B2(
        \REGISTERS[26][30] ), .ZN(n1209) );
  OAI221_X1 U1646 ( .B1(n2119), .B2(n57), .C1(n2087), .C2(n54), .A(n1210), 
        .ZN(n1203) );
  AOI22_X1 U1647 ( .A1(n51), .A2(\REGISTERS[29][30] ), .B1(n46), .B2(
        \REGISTERS[28][30] ), .ZN(n1210) );
  OAI221_X1 U1648 ( .B1(n1799), .B2(n24), .C1(n509), .C2(n21), .A(n1217), .ZN(
        n1212) );
  AOI22_X1 U1649 ( .A1(n18), .A2(\REGISTERS[11][30] ), .B1(n13), .B2(
        \REGISTERS[10][30] ), .ZN(n1217) );
  OAI221_X1 U1650 ( .B1(n2054), .B2(n69), .C1(n2022), .C2(n66), .A(n1169), 
        .ZN(n1154) );
  AOI22_X1 U1651 ( .A1(n63), .A2(\REGISTERS[27][31] ), .B1(n58), .B2(
        \REGISTERS[26][31] ), .ZN(n1169) );
  OAI221_X1 U1652 ( .B1(n2118), .B2(n57), .C1(n2086), .C2(n54), .A(n1174), 
        .ZN(n1153) );
  AOI22_X1 U1653 ( .A1(n51), .A2(\REGISTERS[29][31] ), .B1(n46), .B2(
        \REGISTERS[28][31] ), .ZN(n1174) );
  OAI221_X1 U1654 ( .B1(n1798), .B2(n24), .C1(n508), .C2(n21), .A(n1193), .ZN(
        n1178) );
  AOI22_X1 U1655 ( .A1(n18), .A2(\REGISTERS[11][31] ), .B1(n13), .B2(
        \REGISTERS[10][31] ), .ZN(n1193) );
  AOI22_X1 U1656 ( .A1(\REGISTERS[3][24] ), .A2(n135), .B1(\REGISTERS[2][24] ), 
        .B2(n132), .ZN(n699) );
  AOI22_X1 U1657 ( .A1(\REGISTERS[3][25] ), .A2(n135), .B1(\REGISTERS[2][25] ), 
        .B2(n132), .ZN(n681) );
  AOI22_X1 U1658 ( .A1(\REGISTERS[3][26] ), .A2(n135), .B1(\REGISTERS[2][26] ), 
        .B2(n132), .ZN(n663) );
  AOI22_X1 U1659 ( .A1(\REGISTERS[3][27] ), .A2(n135), .B1(\REGISTERS[2][27] ), 
        .B2(n132), .ZN(n645) );
  AOI22_X1 U1660 ( .A1(\REGISTERS[3][28] ), .A2(n135), .B1(\REGISTERS[2][28] ), 
        .B2(n132), .ZN(n627) );
  AOI22_X1 U1661 ( .A1(\REGISTERS[3][29] ), .A2(n135), .B1(\REGISTERS[2][29] ), 
        .B2(n132), .ZN(n609) );
  AOI22_X1 U1662 ( .A1(\REGISTERS[3][30] ), .A2(n135), .B1(\REGISTERS[2][30] ), 
        .B2(n132), .ZN(n591) );
  AOI22_X1 U1663 ( .A1(\REGISTERS[3][31] ), .A2(n135), .B1(\REGISTERS[2][31] ), 
        .B2(n132), .ZN(n559) );
  AOI22_X1 U1664 ( .A1(\REGISTERS[3][0] ), .A2(n133), .B1(\REGISTERS[2][0] ), 
        .B2(n130), .ZN(n1141) );
  AOI22_X1 U1665 ( .A1(\REGISTERS[3][1] ), .A2(n133), .B1(\REGISTERS[2][1] ), 
        .B2(n130), .ZN(n1113) );
  AOI22_X1 U1666 ( .A1(\REGISTERS[3][2] ), .A2(n133), .B1(\REGISTERS[2][2] ), 
        .B2(n130), .ZN(n1095) );
  AOI22_X1 U1667 ( .A1(\REGISTERS[3][3] ), .A2(n133), .B1(\REGISTERS[2][3] ), 
        .B2(n130), .ZN(n1077) );
  AOI22_X1 U1668 ( .A1(\REGISTERS[3][4] ), .A2(n133), .B1(\REGISTERS[2][4] ), 
        .B2(n130), .ZN(n1059) );
  AOI22_X1 U1669 ( .A1(\REGISTERS[3][5] ), .A2(n133), .B1(\REGISTERS[2][5] ), 
        .B2(n130), .ZN(n1041) );
  AOI22_X1 U1670 ( .A1(\REGISTERS[3][6] ), .A2(n133), .B1(\REGISTERS[2][6] ), 
        .B2(n130), .ZN(n1023) );
  AOI22_X1 U1671 ( .A1(\REGISTERS[3][7] ), .A2(n133), .B1(\REGISTERS[2][7] ), 
        .B2(n130), .ZN(n1005) );
  AOI22_X1 U1672 ( .A1(\REGISTERS[3][8] ), .A2(n133), .B1(\REGISTERS[2][8] ), 
        .B2(n130), .ZN(n987) );
  AOI22_X1 U1673 ( .A1(\REGISTERS[3][9] ), .A2(n133), .B1(\REGISTERS[2][9] ), 
        .B2(n130), .ZN(n969) );
  AOI22_X1 U1674 ( .A1(\REGISTERS[3][10] ), .A2(n133), .B1(\REGISTERS[2][10] ), 
        .B2(n130), .ZN(n951) );
  AOI22_X1 U1675 ( .A1(\REGISTERS[3][11] ), .A2(n133), .B1(\REGISTERS[2][11] ), 
        .B2(n130), .ZN(n933) );
  AOI22_X1 U1676 ( .A1(\REGISTERS[3][12] ), .A2(n134), .B1(\REGISTERS[2][12] ), 
        .B2(n131), .ZN(n915) );
  AOI22_X1 U1677 ( .A1(\REGISTERS[3][13] ), .A2(n134), .B1(\REGISTERS[2][13] ), 
        .B2(n131), .ZN(n897) );
  AOI22_X1 U1678 ( .A1(\REGISTERS[3][14] ), .A2(n134), .B1(\REGISTERS[2][14] ), 
        .B2(n131), .ZN(n879) );
  AOI22_X1 U1679 ( .A1(\REGISTERS[3][15] ), .A2(n134), .B1(\REGISTERS[2][15] ), 
        .B2(n131), .ZN(n861) );
  AOI22_X1 U1680 ( .A1(\REGISTERS[3][16] ), .A2(n134), .B1(\REGISTERS[2][16] ), 
        .B2(n131), .ZN(n843) );
  AOI22_X1 U1681 ( .A1(\REGISTERS[3][17] ), .A2(n134), .B1(\REGISTERS[2][17] ), 
        .B2(n131), .ZN(n825) );
  AOI22_X1 U1682 ( .A1(\REGISTERS[3][18] ), .A2(n134), .B1(\REGISTERS[2][18] ), 
        .B2(n131), .ZN(n807) );
  AOI22_X1 U1683 ( .A1(\REGISTERS[3][19] ), .A2(n134), .B1(\REGISTERS[2][19] ), 
        .B2(n131), .ZN(n789) );
  AOI22_X1 U1684 ( .A1(\REGISTERS[3][20] ), .A2(n134), .B1(\REGISTERS[2][20] ), 
        .B2(n131), .ZN(n771) );
  AOI22_X1 U1685 ( .A1(\REGISTERS[3][21] ), .A2(n134), .B1(\REGISTERS[2][21] ), 
        .B2(n131), .ZN(n753) );
  AOI22_X1 U1686 ( .A1(\REGISTERS[3][22] ), .A2(n134), .B1(\REGISTERS[2][22] ), 
        .B2(n131), .ZN(n735) );
  AOI22_X1 U1687 ( .A1(\REGISTERS[3][23] ), .A2(n134), .B1(\REGISTERS[2][23] ), 
        .B2(n131), .ZN(n717) );
  OAI21_X1 U1688 ( .B1(n419), .B2(n45), .A(n1323), .ZN(n1322) );
  AOI22_X1 U1689 ( .A1(n42), .A2(\REGISTERS[3][24] ), .B1(n37), .B2(
        \REGISTERS[2][24] ), .ZN(n1323) );
  OAI21_X1 U1690 ( .B1(n418), .B2(n45), .A(n1305), .ZN(n1304) );
  AOI22_X1 U1691 ( .A1(n42), .A2(\REGISTERS[3][25] ), .B1(n37), .B2(
        \REGISTERS[2][25] ), .ZN(n1305) );
  OAI21_X1 U1692 ( .B1(n417), .B2(n45), .A(n1287), .ZN(n1286) );
  AOI22_X1 U1693 ( .A1(n42), .A2(\REGISTERS[3][26] ), .B1(n37), .B2(
        \REGISTERS[2][26] ), .ZN(n1287) );
  OAI21_X1 U1694 ( .B1(n416), .B2(n45), .A(n1269), .ZN(n1268) );
  AOI22_X1 U1695 ( .A1(n42), .A2(\REGISTERS[3][27] ), .B1(n37), .B2(
        \REGISTERS[2][27] ), .ZN(n1269) );
  OAI21_X1 U1696 ( .B1(n415), .B2(n45), .A(n1251), .ZN(n1250) );
  AOI22_X1 U1697 ( .A1(n42), .A2(\REGISTERS[3][28] ), .B1(n37), .B2(
        \REGISTERS[2][28] ), .ZN(n1251) );
  OAI21_X1 U1698 ( .B1(n414), .B2(n45), .A(n1233), .ZN(n1232) );
  AOI22_X1 U1699 ( .A1(n42), .A2(\REGISTERS[3][29] ), .B1(n37), .B2(
        \REGISTERS[2][29] ), .ZN(n1233) );
  OAI21_X1 U1700 ( .B1(n413), .B2(n45), .A(n1215), .ZN(n1214) );
  AOI22_X1 U1701 ( .A1(n42), .A2(\REGISTERS[3][30] ), .B1(n37), .B2(
        \REGISTERS[2][30] ), .ZN(n1215) );
  OAI21_X1 U1702 ( .B1(n412), .B2(n45), .A(n1183), .ZN(n1180) );
  AOI22_X1 U1703 ( .A1(n42), .A2(\REGISTERS[3][31] ), .B1(n37), .B2(
        \REGISTERS[2][31] ), .ZN(n1183) );
  OAI21_X1 U1704 ( .B1(n443), .B2(n43), .A(n1765), .ZN(n1764) );
  AOI22_X1 U1705 ( .A1(n40), .A2(\REGISTERS[3][0] ), .B1(n39), .B2(
        \REGISTERS[2][0] ), .ZN(n1765) );
  OAI21_X1 U1706 ( .B1(n442), .B2(n43), .A(n1737), .ZN(n1736) );
  AOI22_X1 U1707 ( .A1(n40), .A2(\REGISTERS[3][1] ), .B1(n39), .B2(
        \REGISTERS[2][1] ), .ZN(n1737) );
  OAI21_X1 U1708 ( .B1(n441), .B2(n43), .A(n1719), .ZN(n1718) );
  AOI22_X1 U1709 ( .A1(n40), .A2(\REGISTERS[3][2] ), .B1(n39), .B2(
        \REGISTERS[2][2] ), .ZN(n1719) );
  OAI21_X1 U1710 ( .B1(n440), .B2(n43), .A(n1701), .ZN(n1700) );
  AOI22_X1 U1711 ( .A1(n40), .A2(\REGISTERS[3][3] ), .B1(n39), .B2(
        \REGISTERS[2][3] ), .ZN(n1701) );
  OAI21_X1 U1712 ( .B1(n439), .B2(n43), .A(n1683), .ZN(n1682) );
  AOI22_X1 U1713 ( .A1(n40), .A2(\REGISTERS[3][4] ), .B1(n39), .B2(
        \REGISTERS[2][4] ), .ZN(n1683) );
  OAI21_X1 U1714 ( .B1(n438), .B2(n43), .A(n1665), .ZN(n1664) );
  AOI22_X1 U1715 ( .A1(n40), .A2(\REGISTERS[3][5] ), .B1(n39), .B2(
        \REGISTERS[2][5] ), .ZN(n1665) );
  OAI21_X1 U1716 ( .B1(n437), .B2(n43), .A(n1647), .ZN(n1646) );
  AOI22_X1 U1717 ( .A1(n40), .A2(\REGISTERS[3][6] ), .B1(n39), .B2(
        \REGISTERS[2][6] ), .ZN(n1647) );
  OAI21_X1 U1718 ( .B1(n436), .B2(n43), .A(n1629), .ZN(n1628) );
  AOI22_X1 U1719 ( .A1(n40), .A2(\REGISTERS[3][7] ), .B1(n39), .B2(
        \REGISTERS[2][7] ), .ZN(n1629) );
  OAI21_X1 U1720 ( .B1(n435), .B2(n43), .A(n1611), .ZN(n1610) );
  AOI22_X1 U1721 ( .A1(n40), .A2(\REGISTERS[3][8] ), .B1(n38), .B2(
        \REGISTERS[2][8] ), .ZN(n1611) );
  OAI21_X1 U1722 ( .B1(n434), .B2(n43), .A(n1593), .ZN(n1592) );
  AOI22_X1 U1723 ( .A1(n40), .A2(\REGISTERS[3][9] ), .B1(n38), .B2(
        \REGISTERS[2][9] ), .ZN(n1593) );
  OAI21_X1 U1724 ( .B1(n433), .B2(n43), .A(n1575), .ZN(n1574) );
  AOI22_X1 U1725 ( .A1(n40), .A2(\REGISTERS[3][10] ), .B1(n38), .B2(
        \REGISTERS[2][10] ), .ZN(n1575) );
  OAI21_X1 U1726 ( .B1(n432), .B2(n43), .A(n1557), .ZN(n1556) );
  AOI22_X1 U1727 ( .A1(n40), .A2(\REGISTERS[3][11] ), .B1(n38), .B2(
        \REGISTERS[2][11] ), .ZN(n1557) );
  OAI21_X1 U1728 ( .B1(n431), .B2(n44), .A(n1539), .ZN(n1538) );
  AOI22_X1 U1729 ( .A1(n41), .A2(\REGISTERS[3][12] ), .B1(n38), .B2(
        \REGISTERS[2][12] ), .ZN(n1539) );
  OAI21_X1 U1730 ( .B1(n430), .B2(n44), .A(n1521), .ZN(n1520) );
  AOI22_X1 U1731 ( .A1(n41), .A2(\REGISTERS[3][13] ), .B1(n38), .B2(
        \REGISTERS[2][13] ), .ZN(n1521) );
  OAI21_X1 U1732 ( .B1(n429), .B2(n44), .A(n1503), .ZN(n1502) );
  AOI22_X1 U1733 ( .A1(n41), .A2(\REGISTERS[3][14] ), .B1(n38), .B2(
        \REGISTERS[2][14] ), .ZN(n1503) );
  OAI21_X1 U1734 ( .B1(n428), .B2(n44), .A(n1485), .ZN(n1484) );
  AOI22_X1 U1735 ( .A1(n41), .A2(\REGISTERS[3][15] ), .B1(n38), .B2(
        \REGISTERS[2][15] ), .ZN(n1485) );
  OAI21_X1 U1736 ( .B1(n427), .B2(n44), .A(n1467), .ZN(n1466) );
  AOI22_X1 U1737 ( .A1(n41), .A2(\REGISTERS[3][16] ), .B1(n38), .B2(
        \REGISTERS[2][16] ), .ZN(n1467) );
  OAI21_X1 U1738 ( .B1(n426), .B2(n44), .A(n1449), .ZN(n1448) );
  AOI22_X1 U1739 ( .A1(n41), .A2(\REGISTERS[3][17] ), .B1(n38), .B2(
        \REGISTERS[2][17] ), .ZN(n1449) );
  OAI21_X1 U1740 ( .B1(n425), .B2(n44), .A(n1431), .ZN(n1430) );
  AOI22_X1 U1741 ( .A1(n41), .A2(\REGISTERS[3][18] ), .B1(n38), .B2(
        \REGISTERS[2][18] ), .ZN(n1431) );
  OAI21_X1 U1742 ( .B1(n424), .B2(n44), .A(n1413), .ZN(n1412) );
  AOI22_X1 U1743 ( .A1(n41), .A2(\REGISTERS[3][19] ), .B1(n38), .B2(
        \REGISTERS[2][19] ), .ZN(n1413) );
  OAI21_X1 U1744 ( .B1(n423), .B2(n44), .A(n1395), .ZN(n1394) );
  AOI22_X1 U1745 ( .A1(n41), .A2(\REGISTERS[3][20] ), .B1(n37), .B2(
        \REGISTERS[2][20] ), .ZN(n1395) );
  OAI21_X1 U1746 ( .B1(n422), .B2(n44), .A(n1377), .ZN(n1376) );
  AOI22_X1 U1747 ( .A1(n41), .A2(\REGISTERS[3][21] ), .B1(n37), .B2(
        \REGISTERS[2][21] ), .ZN(n1377) );
  OAI21_X1 U1748 ( .B1(n421), .B2(n44), .A(n1359), .ZN(n1358) );
  AOI22_X1 U1749 ( .A1(n41), .A2(\REGISTERS[3][22] ), .B1(n37), .B2(
        \REGISTERS[2][22] ), .ZN(n1359) );
  OAI21_X1 U1750 ( .B1(n420), .B2(n44), .A(n1341), .ZN(n1340) );
  AOI22_X1 U1751 ( .A1(n41), .A2(\REGISTERS[3][23] ), .B1(n37), .B2(
        \REGISTERS[2][23] ), .ZN(n1341) );
  INV_X1 U1752 ( .A(ADD_WR[2]), .ZN(n409) );
  INV_X1 U1753 ( .A(ADD_WR[0]), .ZN(n411) );
  INV_X1 U1754 ( .A(ADD_WR[1]), .ZN(n410) );
  INV_X1 U1755 ( .A(ADD_WR[3]), .ZN(n408) );
  INV_X1 U1756 ( .A(ADD_WR[4]), .ZN(n407) );
  OR2_X1 U1757 ( .A1(RE), .A2(n391), .ZN(N307) );
  INV_X1 U1758 ( .A(\REGISTERS[17][0] ), .ZN(n1957) );
  INV_X1 U1759 ( .A(\REGISTERS[21][0] ), .ZN(n2021) );
  INV_X1 U1760 ( .A(\REGISTERS[25][0] ), .ZN(n2085) );
  INV_X1 U1761 ( .A(\REGISTERS[31][0] ), .ZN(n2149) );
  INV_X1 U1762 ( .A(\REGISTERS[5][0] ), .ZN(n507) );
  INV_X1 U1763 ( .A(\REGISTERS[9][0] ), .ZN(n1829) );
  INV_X1 U1764 ( .A(\REGISTERS[13][0] ), .ZN(n1893) );
  INV_X1 U1765 ( .A(\REGISTERS[17][1] ), .ZN(n1956) );
  INV_X1 U1766 ( .A(\REGISTERS[21][1] ), .ZN(n2020) );
  INV_X1 U1767 ( .A(\REGISTERS[25][1] ), .ZN(n2084) );
  INV_X1 U1768 ( .A(\REGISTERS[31][1] ), .ZN(n2148) );
  INV_X1 U1769 ( .A(\REGISTERS[5][1] ), .ZN(n506) );
  INV_X1 U1770 ( .A(\REGISTERS[9][1] ), .ZN(n1828) );
  INV_X1 U1771 ( .A(\REGISTERS[13][1] ), .ZN(n1892) );
  INV_X1 U1772 ( .A(\REGISTERS[17][2] ), .ZN(n1955) );
  INV_X1 U1773 ( .A(\REGISTERS[21][2] ), .ZN(n2019) );
  INV_X1 U1774 ( .A(\REGISTERS[25][2] ), .ZN(n2083) );
  INV_X1 U1775 ( .A(\REGISTERS[31][2] ), .ZN(n2147) );
  INV_X1 U1776 ( .A(\REGISTERS[5][2] ), .ZN(n505) );
  INV_X1 U1777 ( .A(\REGISTERS[9][2] ), .ZN(n1827) );
  INV_X1 U1778 ( .A(\REGISTERS[13][2] ), .ZN(n1891) );
  INV_X1 U1779 ( .A(\REGISTERS[17][3] ), .ZN(n1954) );
  INV_X1 U1780 ( .A(\REGISTERS[21][3] ), .ZN(n2018) );
  INV_X1 U1781 ( .A(\REGISTERS[25][3] ), .ZN(n2082) );
  INV_X1 U1782 ( .A(\REGISTERS[31][3] ), .ZN(n2146) );
  INV_X1 U1783 ( .A(\REGISTERS[5][3] ), .ZN(n504) );
  INV_X1 U1784 ( .A(\REGISTERS[9][3] ), .ZN(n1826) );
  INV_X1 U1785 ( .A(\REGISTERS[13][3] ), .ZN(n1890) );
  INV_X1 U1786 ( .A(\REGISTERS[17][4] ), .ZN(n1953) );
  INV_X1 U1787 ( .A(\REGISTERS[21][4] ), .ZN(n2017) );
  INV_X1 U1788 ( .A(\REGISTERS[25][4] ), .ZN(n2081) );
  INV_X1 U1789 ( .A(\REGISTERS[31][4] ), .ZN(n2145) );
  INV_X1 U1790 ( .A(\REGISTERS[5][4] ), .ZN(n503) );
  INV_X1 U1791 ( .A(\REGISTERS[9][4] ), .ZN(n1825) );
  INV_X1 U1792 ( .A(\REGISTERS[13][4] ), .ZN(n1889) );
  INV_X1 U1793 ( .A(\REGISTERS[17][5] ), .ZN(n1952) );
  INV_X1 U1794 ( .A(\REGISTERS[21][5] ), .ZN(n2016) );
  INV_X1 U1795 ( .A(\REGISTERS[25][5] ), .ZN(n2080) );
  INV_X1 U1796 ( .A(\REGISTERS[31][5] ), .ZN(n2144) );
  INV_X1 U1797 ( .A(\REGISTERS[5][5] ), .ZN(n502) );
  INV_X1 U1798 ( .A(\REGISTERS[9][5] ), .ZN(n1824) );
  INV_X1 U1799 ( .A(\REGISTERS[13][5] ), .ZN(n1888) );
  INV_X1 U1800 ( .A(\REGISTERS[17][6] ), .ZN(n1951) );
  INV_X1 U1801 ( .A(\REGISTERS[21][6] ), .ZN(n2015) );
  INV_X1 U1802 ( .A(\REGISTERS[25][6] ), .ZN(n2079) );
  INV_X1 U1803 ( .A(\REGISTERS[31][6] ), .ZN(n2143) );
  INV_X1 U1804 ( .A(\REGISTERS[5][6] ), .ZN(n501) );
  INV_X1 U1805 ( .A(\REGISTERS[9][6] ), .ZN(n1823) );
  INV_X1 U1806 ( .A(\REGISTERS[13][6] ), .ZN(n1887) );
  INV_X1 U1807 ( .A(\REGISTERS[17][7] ), .ZN(n1950) );
  INV_X1 U1808 ( .A(\REGISTERS[21][7] ), .ZN(n2014) );
  INV_X1 U1809 ( .A(\REGISTERS[25][7] ), .ZN(n2078) );
  INV_X1 U1810 ( .A(\REGISTERS[31][7] ), .ZN(n2142) );
  INV_X1 U1811 ( .A(\REGISTERS[5][7] ), .ZN(n500) );
  INV_X1 U1812 ( .A(\REGISTERS[9][7] ), .ZN(n1822) );
  INV_X1 U1813 ( .A(\REGISTERS[13][7] ), .ZN(n1886) );
  INV_X1 U1814 ( .A(\REGISTERS[17][8] ), .ZN(n1949) );
  INV_X1 U1815 ( .A(\REGISTERS[21][8] ), .ZN(n2013) );
  INV_X1 U1816 ( .A(\REGISTERS[25][8] ), .ZN(n2077) );
  INV_X1 U1817 ( .A(\REGISTERS[31][8] ), .ZN(n2141) );
  INV_X1 U1818 ( .A(\REGISTERS[5][8] ), .ZN(n499) );
  INV_X1 U1819 ( .A(\REGISTERS[9][8] ), .ZN(n1821) );
  INV_X1 U1820 ( .A(\REGISTERS[13][8] ), .ZN(n1885) );
  INV_X1 U1821 ( .A(\REGISTERS[17][9] ), .ZN(n1948) );
  INV_X1 U1822 ( .A(\REGISTERS[21][9] ), .ZN(n2012) );
  INV_X1 U1823 ( .A(\REGISTERS[25][9] ), .ZN(n2076) );
  INV_X1 U1824 ( .A(\REGISTERS[31][9] ), .ZN(n2140) );
  INV_X1 U1825 ( .A(\REGISTERS[5][9] ), .ZN(n498) );
  INV_X1 U1826 ( .A(\REGISTERS[9][9] ), .ZN(n1820) );
  INV_X1 U1827 ( .A(\REGISTERS[13][9] ), .ZN(n1884) );
  INV_X1 U1828 ( .A(\REGISTERS[17][10] ), .ZN(n1947) );
  INV_X1 U1829 ( .A(\REGISTERS[21][10] ), .ZN(n2011) );
  INV_X1 U1830 ( .A(\REGISTERS[25][10] ), .ZN(n2075) );
  INV_X1 U1831 ( .A(\REGISTERS[31][10] ), .ZN(n2139) );
  INV_X1 U1832 ( .A(\REGISTERS[5][10] ), .ZN(n497) );
  INV_X1 U1833 ( .A(\REGISTERS[9][10] ), .ZN(n1819) );
  INV_X1 U1834 ( .A(\REGISTERS[13][10] ), .ZN(n1883) );
  INV_X1 U1835 ( .A(\REGISTERS[17][11] ), .ZN(n1946) );
  INV_X1 U1836 ( .A(\REGISTERS[21][11] ), .ZN(n2010) );
  INV_X1 U1837 ( .A(\REGISTERS[25][11] ), .ZN(n2074) );
  INV_X1 U1838 ( .A(\REGISTERS[31][11] ), .ZN(n2138) );
  INV_X1 U1839 ( .A(\REGISTERS[5][11] ), .ZN(n496) );
  INV_X1 U1840 ( .A(\REGISTERS[9][11] ), .ZN(n1818) );
  INV_X1 U1841 ( .A(\REGISTERS[13][11] ), .ZN(n1882) );
  INV_X1 U1842 ( .A(\REGISTERS[17][12] ), .ZN(n1945) );
  INV_X1 U1843 ( .A(\REGISTERS[21][12] ), .ZN(n2009) );
  INV_X1 U1844 ( .A(\REGISTERS[25][12] ), .ZN(n2073) );
  INV_X1 U1845 ( .A(\REGISTERS[31][12] ), .ZN(n2137) );
  INV_X1 U1846 ( .A(\REGISTERS[5][12] ), .ZN(n495) );
  INV_X1 U1847 ( .A(\REGISTERS[9][12] ), .ZN(n1817) );
  INV_X1 U1848 ( .A(\REGISTERS[13][12] ), .ZN(n1881) );
  INV_X1 U1849 ( .A(\REGISTERS[17][13] ), .ZN(n1944) );
  INV_X1 U1850 ( .A(\REGISTERS[21][13] ), .ZN(n2008) );
  INV_X1 U1851 ( .A(\REGISTERS[25][13] ), .ZN(n2072) );
  INV_X1 U1852 ( .A(\REGISTERS[31][13] ), .ZN(n2136) );
  INV_X1 U1853 ( .A(\REGISTERS[5][13] ), .ZN(n494) );
  INV_X1 U1854 ( .A(\REGISTERS[9][13] ), .ZN(n1816) );
  INV_X1 U1855 ( .A(\REGISTERS[13][13] ), .ZN(n1880) );
  INV_X1 U1856 ( .A(\REGISTERS[17][14] ), .ZN(n1943) );
  INV_X1 U1857 ( .A(\REGISTERS[21][14] ), .ZN(n2007) );
  INV_X1 U1858 ( .A(\REGISTERS[25][14] ), .ZN(n2071) );
  INV_X1 U1859 ( .A(\REGISTERS[31][14] ), .ZN(n2135) );
  INV_X1 U1860 ( .A(\REGISTERS[5][14] ), .ZN(n493) );
  INV_X1 U1861 ( .A(\REGISTERS[9][14] ), .ZN(n1815) );
  INV_X1 U1862 ( .A(\REGISTERS[13][14] ), .ZN(n1879) );
  INV_X1 U1863 ( .A(\REGISTERS[17][15] ), .ZN(n1942) );
  INV_X1 U1864 ( .A(\REGISTERS[21][15] ), .ZN(n2006) );
  INV_X1 U1865 ( .A(\REGISTERS[25][15] ), .ZN(n2070) );
  INV_X1 U1866 ( .A(\REGISTERS[31][15] ), .ZN(n2134) );
  INV_X1 U1867 ( .A(\REGISTERS[5][15] ), .ZN(n492) );
  INV_X1 U1868 ( .A(\REGISTERS[9][15] ), .ZN(n1814) );
  INV_X1 U1869 ( .A(\REGISTERS[13][15] ), .ZN(n1878) );
  INV_X1 U1870 ( .A(\REGISTERS[17][16] ), .ZN(n1941) );
  INV_X1 U1871 ( .A(\REGISTERS[21][16] ), .ZN(n2005) );
  INV_X1 U1872 ( .A(\REGISTERS[25][16] ), .ZN(n2069) );
  INV_X1 U1873 ( .A(\REGISTERS[31][16] ), .ZN(n2133) );
  INV_X1 U1874 ( .A(\REGISTERS[5][16] ), .ZN(n491) );
  INV_X1 U1875 ( .A(\REGISTERS[9][16] ), .ZN(n1813) );
  INV_X1 U1876 ( .A(\REGISTERS[13][16] ), .ZN(n1877) );
  INV_X1 U1877 ( .A(\REGISTERS[17][17] ), .ZN(n1940) );
  INV_X1 U1878 ( .A(\REGISTERS[21][17] ), .ZN(n2004) );
  INV_X1 U1879 ( .A(\REGISTERS[25][17] ), .ZN(n2068) );
  INV_X1 U1880 ( .A(\REGISTERS[31][17] ), .ZN(n2132) );
  INV_X1 U1881 ( .A(\REGISTERS[5][17] ), .ZN(n490) );
  INV_X1 U1882 ( .A(\REGISTERS[9][17] ), .ZN(n1812) );
  INV_X1 U1883 ( .A(\REGISTERS[13][17] ), .ZN(n1876) );
  INV_X1 U1884 ( .A(\REGISTERS[17][18] ), .ZN(n1939) );
  INV_X1 U1885 ( .A(\REGISTERS[21][18] ), .ZN(n2003) );
  INV_X1 U1886 ( .A(\REGISTERS[25][18] ), .ZN(n2067) );
  INV_X1 U1887 ( .A(\REGISTERS[31][18] ), .ZN(n2131) );
  INV_X1 U1888 ( .A(\REGISTERS[5][18] ), .ZN(n489) );
  INV_X1 U1889 ( .A(\REGISTERS[9][18] ), .ZN(n1811) );
  INV_X1 U1890 ( .A(\REGISTERS[13][18] ), .ZN(n1875) );
  INV_X1 U1891 ( .A(\REGISTERS[17][19] ), .ZN(n1938) );
  INV_X1 U1892 ( .A(\REGISTERS[21][19] ), .ZN(n2002) );
  INV_X1 U1893 ( .A(\REGISTERS[25][19] ), .ZN(n2066) );
  INV_X1 U1894 ( .A(\REGISTERS[31][19] ), .ZN(n2130) );
  INV_X1 U1895 ( .A(\REGISTERS[5][19] ), .ZN(n488) );
  INV_X1 U1896 ( .A(\REGISTERS[9][19] ), .ZN(n1810) );
  INV_X1 U1897 ( .A(\REGISTERS[13][19] ), .ZN(n1874) );
  INV_X1 U1898 ( .A(\REGISTERS[17][20] ), .ZN(n1937) );
  INV_X1 U1899 ( .A(\REGISTERS[21][20] ), .ZN(n2001) );
  INV_X1 U1900 ( .A(\REGISTERS[25][20] ), .ZN(n2065) );
  INV_X1 U1901 ( .A(\REGISTERS[31][20] ), .ZN(n2129) );
  INV_X1 U1902 ( .A(\REGISTERS[5][20] ), .ZN(n487) );
  INV_X1 U1903 ( .A(\REGISTERS[9][20] ), .ZN(n1809) );
  INV_X1 U1904 ( .A(\REGISTERS[13][20] ), .ZN(n1873) );
  INV_X1 U1917 ( .A(\REGISTERS[17][21] ), .ZN(n1936) );
  INV_X1 U1918 ( .A(\REGISTERS[21][21] ), .ZN(n2000) );
  INV_X1 U1919 ( .A(\REGISTERS[25][21] ), .ZN(n2064) );
  INV_X1 U1920 ( .A(\REGISTERS[31][21] ), .ZN(n2128) );
  INV_X1 U1921 ( .A(\REGISTERS[5][21] ), .ZN(n486) );
  INV_X1 U1922 ( .A(\REGISTERS[9][21] ), .ZN(n1808) );
  INV_X1 U1923 ( .A(\REGISTERS[13][21] ), .ZN(n1872) );
  INV_X1 U1924 ( .A(\REGISTERS[17][22] ), .ZN(n1935) );
  INV_X1 U1925 ( .A(\REGISTERS[21][22] ), .ZN(n1999) );
  INV_X1 U1926 ( .A(\REGISTERS[25][22] ), .ZN(n2063) );
  INV_X1 U1927 ( .A(\REGISTERS[31][22] ), .ZN(n2127) );
  INV_X1 U1928 ( .A(\REGISTERS[5][22] ), .ZN(n485) );
  INV_X1 U1929 ( .A(\REGISTERS[9][22] ), .ZN(n1807) );
  INV_X1 U1930 ( .A(\REGISTERS[13][22] ), .ZN(n1871) );
  INV_X1 U1931 ( .A(\REGISTERS[17][23] ), .ZN(n1934) );
  INV_X1 U1932 ( .A(\REGISTERS[21][23] ), .ZN(n1998) );
  INV_X1 U1933 ( .A(\REGISTERS[25][23] ), .ZN(n2062) );
  INV_X1 U1934 ( .A(\REGISTERS[31][23] ), .ZN(n2126) );
  INV_X1 U1935 ( .A(\REGISTERS[5][23] ), .ZN(n484) );
  INV_X1 U1936 ( .A(\REGISTERS[9][23] ), .ZN(n1806) );
  INV_X1 U1937 ( .A(\REGISTERS[13][23] ), .ZN(n1870) );
  INV_X1 U1938 ( .A(\REGISTERS[17][24] ), .ZN(n1933) );
  INV_X1 U1939 ( .A(\REGISTERS[21][24] ), .ZN(n1997) );
  INV_X1 U1940 ( .A(\REGISTERS[25][24] ), .ZN(n2061) );
  INV_X1 U1941 ( .A(\REGISTERS[31][24] ), .ZN(n2125) );
  INV_X1 U1942 ( .A(\REGISTERS[5][24] ), .ZN(n483) );
  INV_X1 U1943 ( .A(\REGISTERS[9][24] ), .ZN(n1805) );
  INV_X1 U1944 ( .A(\REGISTERS[13][24] ), .ZN(n1869) );
  INV_X1 U1945 ( .A(\REGISTERS[17][25] ), .ZN(n1932) );
  INV_X1 U1946 ( .A(\REGISTERS[21][25] ), .ZN(n1996) );
  INV_X1 U1947 ( .A(\REGISTERS[25][25] ), .ZN(n2060) );
  INV_X1 U1948 ( .A(\REGISTERS[31][25] ), .ZN(n2124) );
  INV_X1 U1949 ( .A(\REGISTERS[5][25] ), .ZN(n482) );
  INV_X1 U1950 ( .A(\REGISTERS[9][25] ), .ZN(n1804) );
  INV_X1 U1951 ( .A(\REGISTERS[13][25] ), .ZN(n1868) );
  INV_X1 U1952 ( .A(\REGISTERS[17][26] ), .ZN(n1931) );
  INV_X1 U1953 ( .A(\REGISTERS[21][26] ), .ZN(n1995) );
  INV_X1 U1954 ( .A(\REGISTERS[25][26] ), .ZN(n2059) );
  INV_X1 U1955 ( .A(\REGISTERS[31][26] ), .ZN(n2123) );
  INV_X1 U1956 ( .A(\REGISTERS[5][26] ), .ZN(n481) );
  INV_X1 U1957 ( .A(\REGISTERS[9][26] ), .ZN(n1803) );
  INV_X1 U1958 ( .A(\REGISTERS[13][26] ), .ZN(n1867) );
  INV_X1 U1959 ( .A(\REGISTERS[17][27] ), .ZN(n1930) );
  INV_X1 U1960 ( .A(\REGISTERS[21][27] ), .ZN(n1994) );
  INV_X1 U1961 ( .A(\REGISTERS[25][27] ), .ZN(n2058) );
  INV_X1 U1962 ( .A(\REGISTERS[31][27] ), .ZN(n2122) );
  INV_X1 U1963 ( .A(\REGISTERS[5][27] ), .ZN(n480) );
  INV_X1 U1964 ( .A(\REGISTERS[9][27] ), .ZN(n1802) );
  INV_X1 U1965 ( .A(\REGISTERS[13][27] ), .ZN(n1866) );
  INV_X1 U1966 ( .A(\REGISTERS[17][28] ), .ZN(n1929) );
  INV_X1 U1967 ( .A(\REGISTERS[21][28] ), .ZN(n1993) );
  INV_X1 U1968 ( .A(\REGISTERS[25][28] ), .ZN(n2057) );
  INV_X1 U1969 ( .A(\REGISTERS[31][28] ), .ZN(n2121) );
  INV_X1 U1970 ( .A(\REGISTERS[5][28] ), .ZN(n479) );
  INV_X1 U1971 ( .A(\REGISTERS[9][28] ), .ZN(n1801) );
  INV_X1 U1972 ( .A(\REGISTERS[13][28] ), .ZN(n1865) );
  INV_X1 U1973 ( .A(\REGISTERS[17][29] ), .ZN(n1928) );
  INV_X1 U1974 ( .A(\REGISTERS[21][29] ), .ZN(n1992) );
  INV_X1 U1975 ( .A(\REGISTERS[25][29] ), .ZN(n2056) );
  INV_X1 U1976 ( .A(\REGISTERS[31][29] ), .ZN(n2120) );
  INV_X1 U1977 ( .A(\REGISTERS[5][29] ), .ZN(n478) );
  INV_X1 U1978 ( .A(\REGISTERS[9][29] ), .ZN(n1800) );
  INV_X1 U1979 ( .A(\REGISTERS[13][29] ), .ZN(n1864) );
  INV_X1 U1980 ( .A(\REGISTERS[17][30] ), .ZN(n1927) );
  INV_X1 U1981 ( .A(\REGISTERS[21][30] ), .ZN(n1991) );
  INV_X1 U1982 ( .A(\REGISTERS[25][30] ), .ZN(n2055) );
  INV_X1 U1983 ( .A(\REGISTERS[31][30] ), .ZN(n2119) );
  INV_X1 U1984 ( .A(\REGISTERS[5][30] ), .ZN(n477) );
  INV_X1 U1985 ( .A(\REGISTERS[9][30] ), .ZN(n1799) );
  INV_X1 U1986 ( .A(\REGISTERS[13][30] ), .ZN(n1863) );
  INV_X1 U1987 ( .A(\REGISTERS[17][31] ), .ZN(n1926) );
  INV_X1 U1988 ( .A(\REGISTERS[21][31] ), .ZN(n1990) );
  INV_X1 U1989 ( .A(\REGISTERS[25][31] ), .ZN(n2054) );
  INV_X1 U1990 ( .A(\REGISTERS[31][31] ), .ZN(n2118) );
  INV_X1 U1991 ( .A(\REGISTERS[5][31] ), .ZN(n476) );
  INV_X1 U1992 ( .A(\REGISTERS[9][31] ), .ZN(n1798) );
  INV_X1 U1993 ( .A(\REGISTERS[13][31] ), .ZN(n1862) );
  INV_X1 U1994 ( .A(\REGISTERS[1][0] ), .ZN(n443) );
  INV_X1 U1995 ( .A(\REGISTERS[1][1] ), .ZN(n442) );
  INV_X1 U1996 ( .A(\REGISTERS[1][2] ), .ZN(n441) );
  INV_X1 U1997 ( .A(\REGISTERS[1][3] ), .ZN(n440) );
  INV_X1 U1998 ( .A(\REGISTERS[1][4] ), .ZN(n439) );
  INV_X1 U1999 ( .A(\REGISTERS[1][5] ), .ZN(n438) );
  INV_X1 U2000 ( .A(\REGISTERS[1][6] ), .ZN(n437) );
  INV_X1 U2001 ( .A(\REGISTERS[1][7] ), .ZN(n436) );
  INV_X1 U2002 ( .A(\REGISTERS[1][8] ), .ZN(n435) );
  INV_X1 U2003 ( .A(\REGISTERS[1][9] ), .ZN(n434) );
  INV_X1 U2004 ( .A(\REGISTERS[1][10] ), .ZN(n433) );
  INV_X1 U2005 ( .A(\REGISTERS[1][11] ), .ZN(n432) );
  INV_X1 U2006 ( .A(\REGISTERS[1][12] ), .ZN(n431) );
  INV_X1 U2007 ( .A(\REGISTERS[1][13] ), .ZN(n430) );
  INV_X1 U2008 ( .A(\REGISTERS[1][14] ), .ZN(n429) );
  INV_X1 U2009 ( .A(\REGISTERS[1][15] ), .ZN(n428) );
  INV_X1 U2010 ( .A(\REGISTERS[1][16] ), .ZN(n427) );
  INV_X1 U2011 ( .A(\REGISTERS[1][17] ), .ZN(n426) );
  INV_X1 U2012 ( .A(\REGISTERS[1][18] ), .ZN(n425) );
  INV_X1 U2013 ( .A(\REGISTERS[1][19] ), .ZN(n424) );
  INV_X1 U2014 ( .A(\REGISTERS[1][20] ), .ZN(n423) );
  INV_X1 U2015 ( .A(\REGISTERS[1][21] ), .ZN(n422) );
  INV_X1 U2016 ( .A(\REGISTERS[1][22] ), .ZN(n421) );
  INV_X1 U2017 ( .A(\REGISTERS[1][23] ), .ZN(n420) );
  INV_X1 U2018 ( .A(\REGISTERS[1][24] ), .ZN(n419) );
  INV_X1 U2019 ( .A(\REGISTERS[1][25] ), .ZN(n418) );
  INV_X1 U2020 ( .A(\REGISTERS[1][26] ), .ZN(n417) );
  INV_X1 U2021 ( .A(\REGISTERS[1][27] ), .ZN(n416) );
  INV_X1 U2022 ( .A(\REGISTERS[1][28] ), .ZN(n415) );
  INV_X1 U2023 ( .A(\REGISTERS[1][29] ), .ZN(n414) );
  INV_X1 U2024 ( .A(\REGISTERS[1][30] ), .ZN(n413) );
  INV_X1 U2025 ( .A(\REGISTERS[1][31] ), .ZN(n412) );
  INV_X1 U2026 ( .A(\REGISTERS[16][0] ), .ZN(n1925) );
  INV_X1 U2027 ( .A(\REGISTERS[20][0] ), .ZN(n1989) );
  INV_X1 U2028 ( .A(\REGISTERS[24][0] ), .ZN(n2053) );
  INV_X1 U2029 ( .A(\REGISTERS[30][0] ), .ZN(n2117) );
  INV_X1 U2030 ( .A(\REGISTERS[4][0] ), .ZN(n475) );
  INV_X1 U2031 ( .A(\REGISTERS[8][0] ), .ZN(n1797) );
  INV_X1 U2032 ( .A(\REGISTERS[12][0] ), .ZN(n1861) );
  INV_X1 U2033 ( .A(\REGISTERS[16][1] ), .ZN(n1924) );
  INV_X1 U2034 ( .A(\REGISTERS[20][1] ), .ZN(n1988) );
  INV_X1 U2035 ( .A(\REGISTERS[24][1] ), .ZN(n2052) );
  INV_X1 U2036 ( .A(\REGISTERS[30][1] ), .ZN(n2116) );
  INV_X1 U2037 ( .A(\REGISTERS[4][1] ), .ZN(n474) );
  INV_X1 U2038 ( .A(\REGISTERS[8][1] ), .ZN(n1796) );
  INV_X1 U2039 ( .A(\REGISTERS[12][1] ), .ZN(n1860) );
  INV_X1 U2040 ( .A(\REGISTERS[16][2] ), .ZN(n1923) );
  INV_X1 U2041 ( .A(\REGISTERS[20][2] ), .ZN(n1987) );
  INV_X1 U2042 ( .A(\REGISTERS[24][2] ), .ZN(n2051) );
  INV_X1 U2043 ( .A(\REGISTERS[30][2] ), .ZN(n2115) );
  INV_X1 U2044 ( .A(\REGISTERS[4][2] ), .ZN(n473) );
  INV_X1 U2045 ( .A(\REGISTERS[8][2] ), .ZN(n1795) );
  INV_X1 U2046 ( .A(\REGISTERS[12][2] ), .ZN(n1859) );
  INV_X1 U2047 ( .A(\REGISTERS[16][3] ), .ZN(n1922) );
  INV_X1 U2048 ( .A(\REGISTERS[20][3] ), .ZN(n1986) );
  INV_X1 U2049 ( .A(\REGISTERS[24][3] ), .ZN(n2050) );
  INV_X1 U2050 ( .A(\REGISTERS[30][3] ), .ZN(n2114) );
  INV_X1 U2051 ( .A(\REGISTERS[4][3] ), .ZN(n472) );
  INV_X1 U2052 ( .A(\REGISTERS[8][3] ), .ZN(n1794) );
  INV_X1 U2053 ( .A(\REGISTERS[12][3] ), .ZN(n1858) );
  INV_X1 U2054 ( .A(\REGISTERS[16][4] ), .ZN(n1921) );
  INV_X1 U2055 ( .A(\REGISTERS[20][4] ), .ZN(n1985) );
  INV_X1 U2056 ( .A(\REGISTERS[24][4] ), .ZN(n2049) );
  INV_X1 U2057 ( .A(\REGISTERS[30][4] ), .ZN(n2113) );
  INV_X1 U2058 ( .A(\REGISTERS[4][4] ), .ZN(n471) );
  INV_X1 U2059 ( .A(\REGISTERS[8][4] ), .ZN(n1793) );
  INV_X1 U2060 ( .A(\REGISTERS[12][4] ), .ZN(n1857) );
  INV_X1 U2061 ( .A(\REGISTERS[16][5] ), .ZN(n1920) );
  INV_X1 U2062 ( .A(\REGISTERS[20][5] ), .ZN(n1984) );
  INV_X1 U2063 ( .A(\REGISTERS[24][5] ), .ZN(n2048) );
  INV_X1 U2064 ( .A(\REGISTERS[30][5] ), .ZN(n2112) );
  INV_X1 U2065 ( .A(\REGISTERS[4][5] ), .ZN(n470) );
  INV_X1 U2066 ( .A(\REGISTERS[8][5] ), .ZN(n1792) );
  INV_X1 U2067 ( .A(\REGISTERS[12][5] ), .ZN(n1856) );
  INV_X1 U2068 ( .A(\REGISTERS[16][6] ), .ZN(n1919) );
  INV_X1 U2069 ( .A(\REGISTERS[20][6] ), .ZN(n1983) );
  INV_X1 U2070 ( .A(\REGISTERS[24][6] ), .ZN(n2047) );
  INV_X1 U2071 ( .A(\REGISTERS[30][6] ), .ZN(n2111) );
  INV_X1 U2072 ( .A(\REGISTERS[4][6] ), .ZN(n469) );
  INV_X1 U2073 ( .A(\REGISTERS[8][6] ), .ZN(n1791) );
  INV_X1 U2074 ( .A(\REGISTERS[12][6] ), .ZN(n1855) );
  INV_X1 U2075 ( .A(\REGISTERS[16][7] ), .ZN(n1918) );
  INV_X1 U2076 ( .A(\REGISTERS[20][7] ), .ZN(n1982) );
  INV_X1 U2077 ( .A(\REGISTERS[24][7] ), .ZN(n2046) );
  INV_X1 U2078 ( .A(\REGISTERS[30][7] ), .ZN(n2110) );
  INV_X1 U2079 ( .A(\REGISTERS[4][7] ), .ZN(n468) );
  INV_X1 U2080 ( .A(\REGISTERS[8][7] ), .ZN(n1790) );
  INV_X1 U2081 ( .A(\REGISTERS[12][7] ), .ZN(n1854) );
  INV_X1 U2082 ( .A(\REGISTERS[16][8] ), .ZN(n1917) );
  INV_X1 U2083 ( .A(\REGISTERS[20][8] ), .ZN(n1981) );
  INV_X1 U2084 ( .A(\REGISTERS[24][8] ), .ZN(n2045) );
  INV_X1 U2085 ( .A(\REGISTERS[30][8] ), .ZN(n2109) );
  INV_X1 U2086 ( .A(\REGISTERS[4][8] ), .ZN(n467) );
  INV_X1 U2087 ( .A(\REGISTERS[8][8] ), .ZN(n1789) );
  INV_X1 U2088 ( .A(\REGISTERS[12][8] ), .ZN(n1853) );
  INV_X1 U2089 ( .A(\REGISTERS[16][9] ), .ZN(n1916) );
  INV_X1 U2090 ( .A(\REGISTERS[20][9] ), .ZN(n1980) );
  INV_X1 U2091 ( .A(\REGISTERS[24][9] ), .ZN(n2044) );
  INV_X1 U2092 ( .A(\REGISTERS[30][9] ), .ZN(n2108) );
  INV_X1 U2093 ( .A(\REGISTERS[4][9] ), .ZN(n466) );
  INV_X1 U2094 ( .A(\REGISTERS[8][9] ), .ZN(n1788) );
  INV_X1 U2095 ( .A(\REGISTERS[12][9] ), .ZN(n1852) );
  INV_X1 U2096 ( .A(\REGISTERS[16][10] ), .ZN(n1915) );
  INV_X1 U2097 ( .A(\REGISTERS[20][10] ), .ZN(n1979) );
  INV_X1 U2098 ( .A(\REGISTERS[24][10] ), .ZN(n2043) );
  INV_X1 U2099 ( .A(\REGISTERS[30][10] ), .ZN(n2107) );
  INV_X1 U2100 ( .A(\REGISTERS[4][10] ), .ZN(n465) );
  INV_X1 U2101 ( .A(\REGISTERS[8][10] ), .ZN(n1787) );
  INV_X1 U2102 ( .A(\REGISTERS[12][10] ), .ZN(n1851) );
  INV_X1 U2103 ( .A(\REGISTERS[16][11] ), .ZN(n1914) );
  INV_X1 U2104 ( .A(\REGISTERS[20][11] ), .ZN(n1978) );
  INV_X1 U2105 ( .A(\REGISTERS[24][11] ), .ZN(n2042) );
  INV_X1 U2106 ( .A(\REGISTERS[30][11] ), .ZN(n2106) );
  INV_X1 U2107 ( .A(\REGISTERS[4][11] ), .ZN(n464) );
  INV_X1 U2108 ( .A(\REGISTERS[8][11] ), .ZN(n1182) );
  INV_X1 U2109 ( .A(\REGISTERS[12][11] ), .ZN(n1850) );
  INV_X1 U2110 ( .A(\REGISTERS[16][12] ), .ZN(n1913) );
  INV_X1 U2111 ( .A(\REGISTERS[20][12] ), .ZN(n1977) );
  INV_X1 U2112 ( .A(\REGISTERS[24][12] ), .ZN(n2041) );
  INV_X1 U2113 ( .A(\REGISTERS[30][12] ), .ZN(n2105) );
  INV_X1 U2114 ( .A(\REGISTERS[4][12] ), .ZN(n463) );
  INV_X1 U2115 ( .A(\REGISTERS[8][12] ), .ZN(n558) );
  INV_X1 U2116 ( .A(\REGISTERS[12][12] ), .ZN(n1849) );
  INV_X1 U2117 ( .A(\REGISTERS[16][13] ), .ZN(n1912) );
  INV_X1 U2118 ( .A(\REGISTERS[20][13] ), .ZN(n1976) );
  INV_X1 U2119 ( .A(\REGISTERS[24][13] ), .ZN(n2040) );
  INV_X1 U2120 ( .A(\REGISTERS[30][13] ), .ZN(n2104) );
  INV_X1 U2121 ( .A(\REGISTERS[4][13] ), .ZN(n462) );
  INV_X1 U2122 ( .A(\REGISTERS[8][13] ), .ZN(n526) );
  INV_X1 U2123 ( .A(\REGISTERS[12][13] ), .ZN(n1848) );
  INV_X1 U2124 ( .A(\REGISTERS[16][14] ), .ZN(n1911) );
  INV_X1 U2125 ( .A(\REGISTERS[20][14] ), .ZN(n1975) );
  INV_X1 U2126 ( .A(\REGISTERS[24][14] ), .ZN(n2039) );
  INV_X1 U2127 ( .A(\REGISTERS[30][14] ), .ZN(n2103) );
  INV_X1 U2128 ( .A(\REGISTERS[4][14] ), .ZN(n461) );
  INV_X1 U2129 ( .A(\REGISTERS[8][14] ), .ZN(n525) );
  INV_X1 U2130 ( .A(\REGISTERS[12][14] ), .ZN(n1847) );
  INV_X1 U2131 ( .A(\REGISTERS[16][15] ), .ZN(n1910) );
  INV_X1 U2132 ( .A(\REGISTERS[20][15] ), .ZN(n1974) );
  INV_X1 U2133 ( .A(\REGISTERS[24][15] ), .ZN(n2038) );
  INV_X1 U2134 ( .A(\REGISTERS[30][15] ), .ZN(n2102) );
  INV_X1 U2135 ( .A(\REGISTERS[4][15] ), .ZN(n460) );
  INV_X1 U2136 ( .A(\REGISTERS[8][15] ), .ZN(n524) );
  INV_X1 U2137 ( .A(\REGISTERS[12][15] ), .ZN(n1846) );
  INV_X1 U2138 ( .A(\REGISTERS[16][16] ), .ZN(n1909) );
  INV_X1 U2139 ( .A(\REGISTERS[20][16] ), .ZN(n1973) );
  INV_X1 U2140 ( .A(\REGISTERS[24][16] ), .ZN(n2037) );
  INV_X1 U2141 ( .A(\REGISTERS[30][16] ), .ZN(n2101) );
  INV_X1 U2142 ( .A(\REGISTERS[4][16] ), .ZN(n459) );
  INV_X1 U2143 ( .A(\REGISTERS[8][16] ), .ZN(n523) );
  INV_X1 U2144 ( .A(\REGISTERS[12][16] ), .ZN(n1845) );
  INV_X1 U2145 ( .A(\REGISTERS[16][17] ), .ZN(n1908) );
  INV_X1 U2146 ( .A(\REGISTERS[20][17] ), .ZN(n1972) );
  INV_X1 U2147 ( .A(\REGISTERS[24][17] ), .ZN(n2036) );
  INV_X1 U2148 ( .A(\REGISTERS[30][17] ), .ZN(n2100) );
  INV_X1 U2149 ( .A(\REGISTERS[4][17] ), .ZN(n458) );
  INV_X1 U2150 ( .A(\REGISTERS[8][17] ), .ZN(n522) );
  INV_X1 U2151 ( .A(\REGISTERS[12][17] ), .ZN(n1844) );
  INV_X1 U2152 ( .A(\REGISTERS[16][18] ), .ZN(n1907) );
  INV_X1 U2153 ( .A(\REGISTERS[20][18] ), .ZN(n1971) );
  INV_X1 U2154 ( .A(\REGISTERS[24][18] ), .ZN(n2035) );
  INV_X1 U2155 ( .A(\REGISTERS[30][18] ), .ZN(n2099) );
  INV_X1 U2156 ( .A(\REGISTERS[4][18] ), .ZN(n457) );
  INV_X1 U2157 ( .A(\REGISTERS[8][18] ), .ZN(n521) );
  INV_X1 U2158 ( .A(\REGISTERS[12][18] ), .ZN(n1843) );
  INV_X1 U2159 ( .A(\REGISTERS[16][19] ), .ZN(n1906) );
  INV_X1 U2160 ( .A(\REGISTERS[20][19] ), .ZN(n1970) );
  INV_X1 U2161 ( .A(\REGISTERS[24][19] ), .ZN(n2034) );
  INV_X1 U2162 ( .A(\REGISTERS[30][19] ), .ZN(n2098) );
  INV_X1 U2163 ( .A(\REGISTERS[4][19] ), .ZN(n456) );
  INV_X1 U2164 ( .A(\REGISTERS[8][19] ), .ZN(n520) );
  INV_X1 U2165 ( .A(\REGISTERS[12][19] ), .ZN(n1842) );
  INV_X1 U2166 ( .A(\REGISTERS[16][20] ), .ZN(n1905) );
  INV_X1 U2167 ( .A(\REGISTERS[20][20] ), .ZN(n1969) );
  INV_X1 U2168 ( .A(\REGISTERS[24][20] ), .ZN(n2033) );
  INV_X1 U2169 ( .A(\REGISTERS[30][20] ), .ZN(n2097) );
  INV_X1 U2170 ( .A(\REGISTERS[4][20] ), .ZN(n455) );
  INV_X1 U2171 ( .A(\REGISTERS[8][20] ), .ZN(n519) );
  INV_X1 U2172 ( .A(\REGISTERS[12][20] ), .ZN(n1841) );
  INV_X1 U2173 ( .A(\REGISTERS[16][21] ), .ZN(n1904) );
  INV_X1 U2174 ( .A(\REGISTERS[20][21] ), .ZN(n1968) );
  INV_X1 U2175 ( .A(\REGISTERS[24][21] ), .ZN(n2032) );
  INV_X1 U2176 ( .A(\REGISTERS[30][21] ), .ZN(n2096) );
  INV_X1 U2177 ( .A(\REGISTERS[4][21] ), .ZN(n454) );
  INV_X1 U2178 ( .A(\REGISTERS[8][21] ), .ZN(n518) );
  INV_X1 U2179 ( .A(\REGISTERS[12][21] ), .ZN(n1840) );
  INV_X1 U2180 ( .A(\REGISTERS[16][22] ), .ZN(n1903) );
  INV_X1 U2181 ( .A(\REGISTERS[20][22] ), .ZN(n1967) );
  INV_X1 U2182 ( .A(\REGISTERS[24][22] ), .ZN(n2031) );
  INV_X1 U2183 ( .A(\REGISTERS[30][22] ), .ZN(n2095) );
  INV_X1 U2184 ( .A(\REGISTERS[4][22] ), .ZN(n453) );
  INV_X1 U2185 ( .A(\REGISTERS[8][22] ), .ZN(n517) );
  INV_X1 U2186 ( .A(\REGISTERS[12][22] ), .ZN(n1839) );
  INV_X1 U2187 ( .A(\REGISTERS[16][23] ), .ZN(n1902) );
  INV_X1 U2188 ( .A(\REGISTERS[20][23] ), .ZN(n1966) );
  INV_X1 U2189 ( .A(\REGISTERS[24][23] ), .ZN(n2030) );
  INV_X1 U2190 ( .A(\REGISTERS[30][23] ), .ZN(n2094) );
  INV_X1 U2191 ( .A(\REGISTERS[4][23] ), .ZN(n452) );
  INV_X1 U2192 ( .A(\REGISTERS[8][23] ), .ZN(n516) );
  INV_X1 U2193 ( .A(\REGISTERS[12][23] ), .ZN(n1838) );
  INV_X1 U2194 ( .A(\REGISTERS[16][24] ), .ZN(n1901) );
  INV_X1 U2195 ( .A(\REGISTERS[20][24] ), .ZN(n1965) );
  INV_X1 U2196 ( .A(\REGISTERS[24][24] ), .ZN(n2029) );
  INV_X1 U2197 ( .A(\REGISTERS[30][24] ), .ZN(n2093) );
  INV_X1 U2198 ( .A(\REGISTERS[4][24] ), .ZN(n451) );
  INV_X1 U2199 ( .A(\REGISTERS[8][24] ), .ZN(n515) );
  INV_X1 U2200 ( .A(\REGISTERS[12][24] ), .ZN(n1837) );
  INV_X1 U2201 ( .A(\REGISTERS[16][25] ), .ZN(n1900) );
  INV_X1 U2202 ( .A(\REGISTERS[20][25] ), .ZN(n1964) );
  INV_X1 U2203 ( .A(\REGISTERS[24][25] ), .ZN(n2028) );
  INV_X1 U2204 ( .A(\REGISTERS[30][25] ), .ZN(n2092) );
  INV_X1 U2205 ( .A(\REGISTERS[4][25] ), .ZN(n450) );
  INV_X1 U2206 ( .A(\REGISTERS[8][25] ), .ZN(n514) );
  INV_X1 U2207 ( .A(\REGISTERS[12][25] ), .ZN(n1836) );
  INV_X1 U2208 ( .A(\REGISTERS[16][26] ), .ZN(n1899) );
  INV_X1 U2209 ( .A(\REGISTERS[20][26] ), .ZN(n1963) );
  INV_X1 U2210 ( .A(\REGISTERS[24][26] ), .ZN(n2027) );
  INV_X1 U2211 ( .A(\REGISTERS[30][26] ), .ZN(n2091) );
  INV_X1 U2212 ( .A(\REGISTERS[4][26] ), .ZN(n449) );
  INV_X1 U2213 ( .A(\REGISTERS[8][26] ), .ZN(n513) );
  INV_X1 U2214 ( .A(\REGISTERS[12][26] ), .ZN(n1835) );
  INV_X1 U2215 ( .A(\REGISTERS[16][27] ), .ZN(n1898) );
  INV_X1 U2216 ( .A(\REGISTERS[20][27] ), .ZN(n1962) );
  INV_X1 U2217 ( .A(\REGISTERS[24][27] ), .ZN(n2026) );
  INV_X1 U2218 ( .A(\REGISTERS[30][27] ), .ZN(n2090) );
  INV_X1 U2219 ( .A(\REGISTERS[4][27] ), .ZN(n448) );
  INV_X1 U2220 ( .A(\REGISTERS[8][27] ), .ZN(n512) );
  INV_X1 U2221 ( .A(\REGISTERS[12][27] ), .ZN(n1834) );
  INV_X1 U2222 ( .A(\REGISTERS[16][28] ), .ZN(n1897) );
  INV_X1 U2223 ( .A(\REGISTERS[20][28] ), .ZN(n1961) );
  INV_X1 U2224 ( .A(\REGISTERS[24][28] ), .ZN(n2025) );
  INV_X1 U2225 ( .A(\REGISTERS[30][28] ), .ZN(n2089) );
  INV_X1 U2226 ( .A(\REGISTERS[4][28] ), .ZN(n447) );
  INV_X1 U2227 ( .A(\REGISTERS[8][28] ), .ZN(n511) );
  INV_X1 U2228 ( .A(\REGISTERS[12][28] ), .ZN(n1833) );
  INV_X1 U2229 ( .A(\REGISTERS[16][29] ), .ZN(n1896) );
  INV_X1 U2230 ( .A(\REGISTERS[20][29] ), .ZN(n1960) );
  INV_X1 U2231 ( .A(\REGISTERS[24][29] ), .ZN(n2024) );
  INV_X1 U2232 ( .A(\REGISTERS[30][29] ), .ZN(n2088) );
  INV_X1 U2233 ( .A(\REGISTERS[4][29] ), .ZN(n446) );
  INV_X1 U2234 ( .A(\REGISTERS[8][29] ), .ZN(n510) );
  INV_X1 U2235 ( .A(\REGISTERS[12][29] ), .ZN(n1832) );
  INV_X1 U2236 ( .A(\REGISTERS[16][30] ), .ZN(n1895) );
  INV_X1 U2237 ( .A(\REGISTERS[20][30] ), .ZN(n1959) );
  INV_X1 U2238 ( .A(\REGISTERS[24][30] ), .ZN(n2023) );
  INV_X1 U2239 ( .A(\REGISTERS[30][30] ), .ZN(n2087) );
  INV_X1 U2240 ( .A(\REGISTERS[4][30] ), .ZN(n445) );
  INV_X1 U2241 ( .A(\REGISTERS[8][30] ), .ZN(n509) );
  INV_X1 U2242 ( .A(\REGISTERS[12][30] ), .ZN(n1831) );
  INV_X1 U2243 ( .A(\REGISTERS[16][31] ), .ZN(n1894) );
  INV_X1 U2244 ( .A(\REGISTERS[20][31] ), .ZN(n1958) );
  INV_X1 U2245 ( .A(\REGISTERS[24][31] ), .ZN(n2022) );
  INV_X1 U2246 ( .A(\REGISTERS[30][31] ), .ZN(n2086) );
  INV_X1 U2247 ( .A(\REGISTERS[4][31] ), .ZN(n444) );
  INV_X1 U2248 ( .A(\REGISTERS[8][31] ), .ZN(n508) );
  INV_X1 U2249 ( .A(\REGISTERS[12][31] ), .ZN(n1830) );
  AND2_X1 U2250 ( .A1(DATAIN[0]), .A2(n406), .ZN(N244) );
  AND2_X1 U2251 ( .A1(DATAIN[1]), .A2(n406), .ZN(N245) );
  AND2_X1 U2252 ( .A1(DATAIN[2]), .A2(n405), .ZN(N246) );
  AND2_X1 U2253 ( .A1(DATAIN[3]), .A2(n405), .ZN(N247) );
  AND2_X1 U2254 ( .A1(DATAIN[4]), .A2(n405), .ZN(N248) );
  AND2_X1 U2255 ( .A1(DATAIN[5]), .A2(n405), .ZN(N249) );
  AND2_X1 U2256 ( .A1(DATAIN[6]), .A2(n405), .ZN(N250) );
  AND2_X1 U2257 ( .A1(DATAIN[7]), .A2(n405), .ZN(N251) );
  AND2_X1 U2258 ( .A1(DATAIN[8]), .A2(n405), .ZN(N252) );
  AND2_X1 U2259 ( .A1(DATAIN[9]), .A2(n402), .ZN(N253) );
  AND2_X1 U2260 ( .A1(DATAIN[10]), .A2(n404), .ZN(N254) );
  AND2_X1 U2261 ( .A1(DATAIN[11]), .A2(n404), .ZN(N255) );
  AND2_X1 U2262 ( .A1(DATAIN[12]), .A2(n404), .ZN(N256) );
  AND2_X1 U2263 ( .A1(DATAIN[13]), .A2(n404), .ZN(N257) );
  AND2_X1 U2264 ( .A1(DATAIN[14]), .A2(n404), .ZN(N258) );
  AND2_X1 U2265 ( .A1(DATAIN[15]), .A2(n404), .ZN(N259) );
  AND2_X1 U2266 ( .A1(DATAIN[16]), .A2(n404), .ZN(N260) );
  AND2_X1 U2267 ( .A1(DATAIN[17]), .A2(n403), .ZN(N261) );
  AND2_X1 U2268 ( .A1(DATAIN[18]), .A2(n403), .ZN(N262) );
  AND2_X1 U2269 ( .A1(DATAIN[19]), .A2(n403), .ZN(N263) );
  AND2_X1 U2270 ( .A1(DATAIN[20]), .A2(n403), .ZN(N264) );
  AND2_X1 U2271 ( .A1(DATAIN[21]), .A2(n403), .ZN(N265) );
  AND2_X1 U2272 ( .A1(DATAIN[22]), .A2(n403), .ZN(N266) );
  AND2_X1 U2273 ( .A1(DATAIN[23]), .A2(n403), .ZN(N267) );
  AND2_X1 U2274 ( .A1(DATAIN[24]), .A2(n402), .ZN(N268) );
  AND2_X1 U2275 ( .A1(DATAIN[25]), .A2(n402), .ZN(N269) );
  AND2_X1 U2276 ( .A1(DATAIN[26]), .A2(n402), .ZN(N270) );
  AND2_X1 U2277 ( .A1(DATAIN[27]), .A2(n402), .ZN(N271) );
  AND2_X1 U2278 ( .A1(DATAIN[28]), .A2(n402), .ZN(N272) );
  AND2_X1 U2279 ( .A1(DATAIN[29]), .A2(n402), .ZN(N273) );
  AND2_X1 U2280 ( .A1(DATAIN[30]), .A2(n401), .ZN(N274) );
  AND2_X1 U2281 ( .A1(DATAIN[31]), .A2(n401), .ZN(N275) );
  CLKBUF_X1 U2282 ( .A(N307), .Z(n187) );
  CLKBUF_X1 U2283 ( .A(N307), .Z(n188) );
  CLKBUF_X1 U2284 ( .A(N307), .Z(n189) );
  CLKBUF_X1 U2285 ( .A(N307), .Z(n190) );
  CLKBUF_X1 U2286 ( .A(N307), .Z(n191) );
  CLKBUF_X1 U2287 ( .A(N307), .Z(n192) );
endmodule


module sign_extender ( d_in, rst, d_ext );
  input [31:0] d_in;
  output [31:0] d_ext;
  input rst;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n1, n2, n3, n4, n5, n6, n7,
         n30;
  assign d_ext[25] = d_ext[31];
  assign d_ext[26] = d_ext[31];
  assign d_ext[27] = d_ext[31];
  assign d_ext[28] = d_ext[31];
  assign d_ext[29] = d_ext[31];
  assign d_ext[30] = d_ext[31];

  OAI33_X1 U56 ( .A1(n5), .A2(d_in[28]), .A3(d_in[27]), .B1(n7), .B2(n27), 
        .B3(n30), .ZN(n26) );
  NAND3_X1 U2 ( .A1(n1), .A2(n10), .A3(n9), .ZN(n11) );
  NOR2_X1 U3 ( .A1(n10), .A2(n2), .ZN(n13) );
  INV_X1 U4 ( .A(rst), .ZN(n2) );
  AOI21_X1 U5 ( .B1(d_in[29]), .B2(d_in[26]), .A(d_in[31]), .ZN(n27) );
  OAI22_X1 U6 ( .A1(n6), .A2(n5), .B1(d_in[28]), .B2(d_in[26]), .ZN(n25) );
  INV_X1 U7 ( .A(d_in[28]), .ZN(n7) );
  NOR2_X1 U8 ( .A1(n8), .A2(n2), .ZN(d_ext[31]) );
  AOI22_X1 U9 ( .A1(n9), .A2(n10), .B1(d_in[25]), .B2(n4), .ZN(n8) );
  INV_X1 U10 ( .A(n10), .ZN(n4) );
  AOI21_X1 U11 ( .B1(n30), .B2(d_in[26]), .A(d_in[31]), .ZN(n28) );
  INV_X1 U12 ( .A(d_in[30]), .ZN(n5) );
  INV_X1 U13 ( .A(d_in[27]), .ZN(n30) );
  AND2_X1 U14 ( .A1(d_in[15]), .A2(n22), .ZN(n9) );
  OAI221_X1 U15 ( .B1(d_in[29]), .B2(n23), .C1(d_in[30]), .C2(n3), .A(n24), 
        .ZN(n22) );
  AND3_X1 U16 ( .A1(n28), .A2(d_in[28]), .A3(d_in[30]), .ZN(n23) );
  AOI21_X1 U17 ( .B1(n25), .B2(n3), .A(n26), .ZN(n24) );
  NAND2_X1 U18 ( .A1(n11), .A2(n21), .ZN(d_ext[16]) );
  NAND2_X1 U19 ( .A1(d_in[16]), .A2(n13), .ZN(n21) );
  NAND2_X1 U20 ( .A1(n11), .A2(n20), .ZN(d_ext[17]) );
  NAND2_X1 U21 ( .A1(d_in[17]), .A2(n13), .ZN(n20) );
  NAND2_X1 U22 ( .A1(n11), .A2(n19), .ZN(d_ext[18]) );
  NAND2_X1 U23 ( .A1(d_in[18]), .A2(n13), .ZN(n19) );
  NAND2_X1 U24 ( .A1(n11), .A2(n18), .ZN(d_ext[19]) );
  NAND2_X1 U25 ( .A1(d_in[19]), .A2(n13), .ZN(n18) );
  NAND2_X1 U26 ( .A1(n11), .A2(n17), .ZN(d_ext[20]) );
  NAND2_X1 U27 ( .A1(d_in[20]), .A2(n13), .ZN(n17) );
  NAND2_X1 U28 ( .A1(n11), .A2(n16), .ZN(d_ext[21]) );
  NAND2_X1 U29 ( .A1(d_in[21]), .A2(n13), .ZN(n16) );
  NAND2_X1 U30 ( .A1(n11), .A2(n15), .ZN(d_ext[22]) );
  NAND2_X1 U31 ( .A1(d_in[22]), .A2(n13), .ZN(n15) );
  NAND2_X1 U32 ( .A1(n11), .A2(n14), .ZN(d_ext[23]) );
  NAND2_X1 U33 ( .A1(d_in[23]), .A2(n13), .ZN(n14) );
  NAND2_X1 U34 ( .A1(n11), .A2(n12), .ZN(d_ext[24]) );
  NAND2_X1 U35 ( .A1(d_in[24]), .A2(n13), .ZN(n12) );
  NAND4_X1 U36 ( .A1(d_in[27]), .A2(n7), .A3(n29), .A4(n6), .ZN(n10) );
  NOR2_X1 U37 ( .A1(d_in[31]), .A2(d_in[30]), .ZN(n29) );
  INV_X1 U38 ( .A(d_in[29]), .ZN(n6) );
  INV_X1 U39 ( .A(d_in[31]), .ZN(n3) );
  AND2_X1 U40 ( .A1(d_in[5]), .A2(n1), .ZN(d_ext[5]) );
  AND2_X1 U41 ( .A1(d_in[0]), .A2(n1), .ZN(d_ext[0]) );
  AND2_X1 U42 ( .A1(d_in[1]), .A2(n1), .ZN(d_ext[1]) );
  AND2_X1 U43 ( .A1(d_in[2]), .A2(n1), .ZN(d_ext[2]) );
  AND2_X1 U44 ( .A1(d_in[3]), .A2(n1), .ZN(d_ext[3]) );
  AND2_X1 U45 ( .A1(d_in[4]), .A2(n1), .ZN(d_ext[4]) );
  AND2_X1 U46 ( .A1(d_in[6]), .A2(n1), .ZN(d_ext[6]) );
  AND2_X1 U47 ( .A1(d_in[7]), .A2(n1), .ZN(d_ext[7]) );
  AND2_X1 U48 ( .A1(d_in[8]), .A2(n1), .ZN(d_ext[8]) );
  AND2_X1 U49 ( .A1(d_in[10]), .A2(n1), .ZN(d_ext[10]) );
  AND2_X1 U50 ( .A1(d_in[13]), .A2(n1), .ZN(d_ext[13]) );
  AND2_X1 U51 ( .A1(d_in[14]), .A2(n1), .ZN(d_ext[14]) );
  AND2_X1 U52 ( .A1(n1), .A2(d_in[9]), .ZN(d_ext[9]) );
  AND2_X1 U53 ( .A1(n1), .A2(d_in[15]), .ZN(d_ext[15]) );
  AND2_X1 U54 ( .A1(d_in[11]), .A2(n1), .ZN(d_ext[11]) );
  AND2_X1 U55 ( .A1(d_in[12]), .A2(n1), .ZN(d_ext[12]) );
  INV_X1 U57 ( .A(n2), .ZN(n1) );
endmodule


module ID_EX ( CLK, RST, NPC_IN, NPC_L_IN, A_IN, B_IN, IMM_IN, RS1_IN, RS2_IN, 
        RD_IN, OPCODE_IN, IR_IN, PR_IN, NPC_OUT, NPC_L_OUT, A_OUT, B_OUT, 
        IMM_OUT, RS1_OUT, RS2_OUT, RD_OUT, OPCODE_OUT, IR_OUT, PR_OUT );
  input [31:0] NPC_IN;
  input [31:0] NPC_L_IN;
  input [31:0] A_IN;
  input [31:0] B_IN;
  input [31:0] IMM_IN;
  input [4:0] RS1_IN;
  input [4:0] RS2_IN;
  input [4:0] RD_IN;
  input [5:0] OPCODE_IN;
  input [15:0] IR_IN;
  output [31:0] NPC_OUT;
  output [31:0] NPC_L_OUT;
  output [31:0] A_OUT;
  output [31:0] B_OUT;
  output [31:0] IMM_OUT;
  output [4:0] RS1_OUT;
  output [4:0] RS2_OUT;
  output [4:0] RD_OUT;
  output [5:0] OPCODE_OUT;
  output [15:0] IR_OUT;
  input CLK, RST, PR_IN;
  output PR_OUT;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23;

  DFFR_X1 PR_OUT_reg ( .D(PR_IN), .CK(CLK), .RN(n7), .Q(PR_OUT) );
  DFFR_X1 \A_OUT_reg[31]  ( .D(A_IN[31]), .CK(CLK), .RN(n7), .Q(A_OUT[31]) );
  DFFR_X1 \A_OUT_reg[30]  ( .D(A_IN[30]), .CK(CLK), .RN(n7), .Q(A_OUT[30]) );
  DFFR_X1 \A_OUT_reg[29]  ( .D(A_IN[29]), .CK(CLK), .RN(n7), .Q(A_OUT[29]) );
  DFFR_X1 \A_OUT_reg[28]  ( .D(A_IN[28]), .CK(CLK), .RN(n7), .Q(A_OUT[28]) );
  DFFR_X1 \A_OUT_reg[27]  ( .D(A_IN[27]), .CK(CLK), .RN(n7), .Q(A_OUT[27]) );
  DFFR_X1 \A_OUT_reg[26]  ( .D(A_IN[26]), .CK(CLK), .RN(n7), .Q(A_OUT[26]) );
  DFFR_X1 \A_OUT_reg[25]  ( .D(A_IN[25]), .CK(CLK), .RN(n7), .Q(A_OUT[25]) );
  DFFR_X1 \A_OUT_reg[24]  ( .D(A_IN[24]), .CK(CLK), .RN(n7), .Q(A_OUT[24]) );
  DFFR_X1 \A_OUT_reg[23]  ( .D(A_IN[23]), .CK(CLK), .RN(n7), .Q(A_OUT[23]) );
  DFFR_X1 \A_OUT_reg[22]  ( .D(A_IN[22]), .CK(CLK), .RN(n7), .Q(A_OUT[22]) );
  DFFR_X1 \A_OUT_reg[21]  ( .D(A_IN[21]), .CK(CLK), .RN(n7), .Q(A_OUT[21]) );
  DFFR_X1 \A_OUT_reg[20]  ( .D(A_IN[20]), .CK(CLK), .RN(n8), .Q(A_OUT[20]) );
  DFFR_X1 \A_OUT_reg[19]  ( .D(A_IN[19]), .CK(CLK), .RN(n8), .Q(A_OUT[19]) );
  DFFR_X1 \A_OUT_reg[18]  ( .D(A_IN[18]), .CK(CLK), .RN(n8), .Q(A_OUT[18]) );
  DFFR_X1 \A_OUT_reg[17]  ( .D(A_IN[17]), .CK(CLK), .RN(n8), .Q(A_OUT[17]) );
  DFFR_X1 \A_OUT_reg[16]  ( .D(A_IN[16]), .CK(CLK), .RN(n8), .Q(A_OUT[16]) );
  DFFR_X1 \A_OUT_reg[15]  ( .D(A_IN[15]), .CK(CLK), .RN(n8), .Q(A_OUT[15]) );
  DFFR_X1 \A_OUT_reg[14]  ( .D(A_IN[14]), .CK(CLK), .RN(n8), .Q(A_OUT[14]) );
  DFFR_X1 \A_OUT_reg[13]  ( .D(A_IN[13]), .CK(CLK), .RN(n8), .Q(A_OUT[13]) );
  DFFR_X1 \A_OUT_reg[12]  ( .D(A_IN[12]), .CK(CLK), .RN(n8), .Q(A_OUT[12]) );
  DFFR_X1 \A_OUT_reg[11]  ( .D(A_IN[11]), .CK(CLK), .RN(n8), .Q(A_OUT[11]) );
  DFFR_X1 \A_OUT_reg[10]  ( .D(A_IN[10]), .CK(CLK), .RN(n8), .Q(A_OUT[10]) );
  DFFR_X1 \A_OUT_reg[9]  ( .D(A_IN[9]), .CK(CLK), .RN(n8), .Q(A_OUT[9]) );
  DFFR_X1 \A_OUT_reg[8]  ( .D(A_IN[8]), .CK(CLK), .RN(n9), .Q(A_OUT[8]) );
  DFFR_X1 \A_OUT_reg[7]  ( .D(A_IN[7]), .CK(CLK), .RN(n9), .Q(A_OUT[7]) );
  DFFR_X1 \A_OUT_reg[6]  ( .D(A_IN[6]), .CK(CLK), .RN(n9), .Q(A_OUT[6]) );
  DFFR_X1 \A_OUT_reg[5]  ( .D(A_IN[5]), .CK(CLK), .RN(n9), .Q(A_OUT[5]) );
  DFFR_X1 \A_OUT_reg[4]  ( .D(A_IN[4]), .CK(CLK), .RN(n9), .Q(A_OUT[4]) );
  DFFR_X1 \A_OUT_reg[3]  ( .D(A_IN[3]), .CK(CLK), .RN(n9), .Q(A_OUT[3]) );
  DFFR_X1 \A_OUT_reg[2]  ( .D(A_IN[2]), .CK(CLK), .RN(n9), .Q(A_OUT[2]) );
  DFFR_X1 \A_OUT_reg[1]  ( .D(A_IN[1]), .CK(CLK), .RN(n9), .Q(A_OUT[1]) );
  DFFR_X1 \A_OUT_reg[0]  ( .D(A_IN[0]), .CK(CLK), .RN(n9), .Q(A_OUT[0]) );
  DFFR_X1 \B_OUT_reg[31]  ( .D(B_IN[31]), .CK(CLK), .RN(n9), .Q(B_OUT[31]) );
  DFFR_X1 \B_OUT_reg[30]  ( .D(B_IN[30]), .CK(CLK), .RN(n9), .Q(B_OUT[30]) );
  DFFR_X1 \B_OUT_reg[29]  ( .D(B_IN[29]), .CK(CLK), .RN(n9), .Q(B_OUT[29]) );
  DFFR_X1 \B_OUT_reg[28]  ( .D(B_IN[28]), .CK(CLK), .RN(n10), .Q(B_OUT[28]) );
  DFFR_X1 \B_OUT_reg[27]  ( .D(B_IN[27]), .CK(CLK), .RN(n10), .Q(B_OUT[27]) );
  DFFR_X1 \B_OUT_reg[26]  ( .D(B_IN[26]), .CK(CLK), .RN(n10), .Q(B_OUT[26]) );
  DFFR_X1 \B_OUT_reg[25]  ( .D(B_IN[25]), .CK(CLK), .RN(n10), .Q(B_OUT[25]) );
  DFFR_X1 \B_OUT_reg[24]  ( .D(B_IN[24]), .CK(CLK), .RN(n10), .Q(B_OUT[24]) );
  DFFR_X1 \B_OUT_reg[23]  ( .D(B_IN[23]), .CK(CLK), .RN(n10), .Q(B_OUT[23]) );
  DFFR_X1 \B_OUT_reg[22]  ( .D(B_IN[22]), .CK(CLK), .RN(n10), .Q(B_OUT[22]) );
  DFFR_X1 \B_OUT_reg[21]  ( .D(B_IN[21]), .CK(CLK), .RN(n10), .Q(B_OUT[21]) );
  DFFR_X1 \B_OUT_reg[20]  ( .D(B_IN[20]), .CK(CLK), .RN(n10), .Q(B_OUT[20]) );
  DFFR_X1 \B_OUT_reg[19]  ( .D(B_IN[19]), .CK(CLK), .RN(n10), .Q(B_OUT[19]) );
  DFFR_X1 \B_OUT_reg[18]  ( .D(B_IN[18]), .CK(CLK), .RN(n10), .Q(B_OUT[18]) );
  DFFR_X1 \B_OUT_reg[17]  ( .D(B_IN[17]), .CK(CLK), .RN(n10), .Q(B_OUT[17]) );
  DFFR_X1 \B_OUT_reg[16]  ( .D(B_IN[16]), .CK(CLK), .RN(n11), .Q(B_OUT[16]) );
  DFFR_X1 \B_OUT_reg[15]  ( .D(B_IN[15]), .CK(CLK), .RN(n11), .Q(B_OUT[15]) );
  DFFR_X1 \B_OUT_reg[14]  ( .D(B_IN[14]), .CK(CLK), .RN(n11), .Q(B_OUT[14]) );
  DFFR_X1 \B_OUT_reg[13]  ( .D(B_IN[13]), .CK(CLK), .RN(n11), .Q(B_OUT[13]) );
  DFFR_X1 \B_OUT_reg[12]  ( .D(B_IN[12]), .CK(CLK), .RN(n11), .Q(B_OUT[12]) );
  DFFR_X1 \B_OUT_reg[11]  ( .D(B_IN[11]), .CK(CLK), .RN(n11), .Q(B_OUT[11]) );
  DFFR_X1 \B_OUT_reg[10]  ( .D(B_IN[10]), .CK(CLK), .RN(n11), .Q(B_OUT[10]) );
  DFFR_X1 \B_OUT_reg[9]  ( .D(B_IN[9]), .CK(CLK), .RN(n11), .Q(B_OUT[9]) );
  DFFR_X1 \B_OUT_reg[8]  ( .D(B_IN[8]), .CK(CLK), .RN(n11), .Q(B_OUT[8]) );
  DFFR_X1 \B_OUT_reg[7]  ( .D(B_IN[7]), .CK(CLK), .RN(n11), .Q(B_OUT[7]) );
  DFFR_X1 \B_OUT_reg[6]  ( .D(B_IN[6]), .CK(CLK), .RN(n11), .Q(B_OUT[6]) );
  DFFR_X1 \B_OUT_reg[5]  ( .D(B_IN[5]), .CK(CLK), .RN(n11), .Q(B_OUT[5]) );
  DFFR_X1 \B_OUT_reg[4]  ( .D(B_IN[4]), .CK(CLK), .RN(n12), .Q(B_OUT[4]) );
  DFFR_X1 \B_OUT_reg[3]  ( .D(B_IN[3]), .CK(CLK), .RN(n12), .Q(B_OUT[3]) );
  DFFR_X1 \B_OUT_reg[2]  ( .D(B_IN[2]), .CK(CLK), .RN(n12), .Q(B_OUT[2]) );
  DFFR_X1 \B_OUT_reg[1]  ( .D(B_IN[1]), .CK(CLK), .RN(n12), .Q(B_OUT[1]) );
  DFFR_X1 \B_OUT_reg[0]  ( .D(B_IN[0]), .CK(CLK), .RN(n12), .Q(B_OUT[0]) );
  DFFR_X1 \IMM_OUT_reg[31]  ( .D(IMM_IN[31]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[31]) );
  DFFR_X1 \IMM_OUT_reg[30]  ( .D(IMM_IN[30]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[30]) );
  DFFR_X1 \IMM_OUT_reg[29]  ( .D(IMM_IN[29]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[29]) );
  DFFR_X1 \IMM_OUT_reg[28]  ( .D(IMM_IN[28]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[28]) );
  DFFR_X1 \IMM_OUT_reg[27]  ( .D(IMM_IN[27]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[27]) );
  DFFR_X1 \IMM_OUT_reg[26]  ( .D(IMM_IN[26]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[26]) );
  DFFR_X1 \IMM_OUT_reg[25]  ( .D(IMM_IN[25]), .CK(CLK), .RN(n12), .Q(
        IMM_OUT[25]) );
  DFFR_X1 \IMM_OUT_reg[24]  ( .D(IMM_IN[24]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[24]) );
  DFFR_X1 \IMM_OUT_reg[23]  ( .D(IMM_IN[23]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[23]) );
  DFFR_X1 \IMM_OUT_reg[22]  ( .D(IMM_IN[22]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[22]) );
  DFFR_X1 \IMM_OUT_reg[21]  ( .D(IMM_IN[21]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[21]) );
  DFFR_X1 \IMM_OUT_reg[20]  ( .D(IMM_IN[20]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[20]) );
  DFFR_X1 \IMM_OUT_reg[19]  ( .D(IMM_IN[19]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[19]) );
  DFFR_X1 \IMM_OUT_reg[18]  ( .D(IMM_IN[18]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[18]) );
  DFFR_X1 \IMM_OUT_reg[17]  ( .D(IMM_IN[17]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[17]) );
  DFFR_X1 \IMM_OUT_reg[16]  ( .D(IMM_IN[16]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[16]) );
  DFFR_X1 \IMM_OUT_reg[15]  ( .D(IMM_IN[15]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[15]) );
  DFFR_X1 \IMM_OUT_reg[14]  ( .D(IMM_IN[14]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[14]) );
  DFFR_X1 \IMM_OUT_reg[13]  ( .D(IMM_IN[13]), .CK(CLK), .RN(n13), .Q(
        IMM_OUT[13]) );
  DFFR_X1 \IMM_OUT_reg[12]  ( .D(IMM_IN[12]), .CK(CLK), .RN(n14), .Q(
        IMM_OUT[12]) );
  DFFR_X1 \IMM_OUT_reg[11]  ( .D(IMM_IN[11]), .CK(CLK), .RN(n14), .Q(
        IMM_OUT[11]) );
  DFFR_X1 \IMM_OUT_reg[10]  ( .D(IMM_IN[10]), .CK(CLK), .RN(n14), .Q(
        IMM_OUT[10]) );
  DFFR_X1 \IMM_OUT_reg[9]  ( .D(IMM_IN[9]), .CK(CLK), .RN(n14), .Q(IMM_OUT[9])
         );
  DFFR_X1 \IMM_OUT_reg[8]  ( .D(IMM_IN[8]), .CK(CLK), .RN(n14), .Q(IMM_OUT[8])
         );
  DFFR_X1 \IMM_OUT_reg[7]  ( .D(IMM_IN[7]), .CK(CLK), .RN(n14), .Q(IMM_OUT[7])
         );
  DFFR_X1 \IMM_OUT_reg[6]  ( .D(IMM_IN[6]), .CK(CLK), .RN(n14), .Q(IMM_OUT[6])
         );
  DFFR_X1 \IMM_OUT_reg[5]  ( .D(IMM_IN[5]), .CK(CLK), .RN(n14), .Q(IMM_OUT[5])
         );
  DFFR_X1 \IMM_OUT_reg[4]  ( .D(IMM_IN[4]), .CK(CLK), .RN(n14), .Q(IMM_OUT[4])
         );
  DFFR_X1 \IMM_OUT_reg[3]  ( .D(IMM_IN[3]), .CK(CLK), .RN(n14), .Q(IMM_OUT[3])
         );
  DFFR_X1 \IMM_OUT_reg[2]  ( .D(IMM_IN[2]), .CK(CLK), .RN(n14), .Q(IMM_OUT[2])
         );
  DFFR_X1 \IMM_OUT_reg[1]  ( .D(IMM_IN[1]), .CK(CLK), .RN(n14), .Q(IMM_OUT[1])
         );
  DFFR_X1 \IMM_OUT_reg[0]  ( .D(IMM_IN[0]), .CK(CLK), .RN(n15), .Q(IMM_OUT[0])
         );
  DFFR_X1 \NPC_OUT_reg[31]  ( .D(NPC_IN[31]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[31]) );
  DFFR_X1 \NPC_OUT_reg[30]  ( .D(NPC_IN[30]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[30]) );
  DFFR_X1 \NPC_OUT_reg[29]  ( .D(NPC_IN[29]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[29]) );
  DFFR_X1 \NPC_OUT_reg[28]  ( .D(NPC_IN[28]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[28]) );
  DFFR_X1 \NPC_OUT_reg[27]  ( .D(NPC_IN[27]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[27]) );
  DFFR_X1 \NPC_OUT_reg[26]  ( .D(NPC_IN[26]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[26]) );
  DFFR_X1 \NPC_OUT_reg[25]  ( .D(NPC_IN[25]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[25]) );
  DFFR_X1 \NPC_OUT_reg[24]  ( .D(NPC_IN[24]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[24]) );
  DFFR_X1 \NPC_OUT_reg[23]  ( .D(NPC_IN[23]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[23]) );
  DFFR_X1 \NPC_OUT_reg[22]  ( .D(NPC_IN[22]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[22]) );
  DFFR_X1 \NPC_OUT_reg[21]  ( .D(NPC_IN[21]), .CK(CLK), .RN(n15), .Q(
        NPC_OUT[21]) );
  DFFR_X1 \NPC_OUT_reg[20]  ( .D(NPC_IN[20]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[20]) );
  DFFR_X1 \NPC_OUT_reg[19]  ( .D(NPC_IN[19]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[19]) );
  DFFR_X1 \NPC_OUT_reg[18]  ( .D(NPC_IN[18]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[18]) );
  DFFR_X1 \NPC_OUT_reg[17]  ( .D(NPC_IN[17]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[17]) );
  DFFR_X1 \NPC_OUT_reg[16]  ( .D(NPC_IN[16]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[16]) );
  DFFR_X1 \NPC_OUT_reg[15]  ( .D(NPC_IN[15]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[15]) );
  DFFR_X1 \NPC_OUT_reg[14]  ( .D(NPC_IN[14]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[14]) );
  DFFR_X1 \NPC_OUT_reg[13]  ( .D(NPC_IN[13]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[13]) );
  DFFR_X1 \NPC_OUT_reg[12]  ( .D(NPC_IN[12]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[12]) );
  DFFR_X1 \NPC_OUT_reg[11]  ( .D(NPC_IN[11]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[11]) );
  DFFR_X1 \NPC_OUT_reg[10]  ( .D(NPC_IN[10]), .CK(CLK), .RN(n16), .Q(
        NPC_OUT[10]) );
  DFFR_X1 \NPC_OUT_reg[9]  ( .D(NPC_IN[9]), .CK(CLK), .RN(n16), .Q(NPC_OUT[9])
         );
  DFFR_X1 \NPC_OUT_reg[8]  ( .D(NPC_IN[8]), .CK(CLK), .RN(n17), .Q(NPC_OUT[8])
         );
  DFFR_X1 \NPC_OUT_reg[7]  ( .D(NPC_IN[7]), .CK(CLK), .RN(n17), .Q(NPC_OUT[7])
         );
  DFFR_X1 \NPC_OUT_reg[6]  ( .D(NPC_IN[6]), .CK(CLK), .RN(n17), .Q(NPC_OUT[6])
         );
  DFFR_X1 \NPC_OUT_reg[5]  ( .D(NPC_IN[5]), .CK(CLK), .RN(n17), .Q(NPC_OUT[5])
         );
  DFFR_X1 \NPC_OUT_reg[4]  ( .D(NPC_IN[4]), .CK(CLK), .RN(n17), .Q(NPC_OUT[4])
         );
  DFFR_X1 \NPC_OUT_reg[3]  ( .D(NPC_IN[3]), .CK(CLK), .RN(n17), .Q(NPC_OUT[3])
         );
  DFFR_X1 \NPC_OUT_reg[2]  ( .D(NPC_IN[2]), .CK(CLK), .RN(n17), .Q(NPC_OUT[2])
         );
  DFFR_X1 \NPC_OUT_reg[1]  ( .D(NPC_IN[1]), .CK(CLK), .RN(n17), .Q(NPC_OUT[1])
         );
  DFFR_X1 \NPC_OUT_reg[0]  ( .D(NPC_IN[0]), .CK(CLK), .RN(n17), .Q(NPC_OUT[0])
         );
  DFFR_X1 \NPC_L_OUT_reg[31]  ( .D(NPC_L_IN[31]), .CK(CLK), .RN(n17), .Q(
        NPC_L_OUT[31]) );
  DFFR_X1 \NPC_L_OUT_reg[30]  ( .D(NPC_L_IN[30]), .CK(CLK), .RN(n17), .Q(
        NPC_L_OUT[30]) );
  DFFR_X1 \NPC_L_OUT_reg[29]  ( .D(NPC_L_IN[29]), .CK(CLK), .RN(n17), .Q(
        NPC_L_OUT[29]) );
  DFFR_X1 \NPC_L_OUT_reg[28]  ( .D(NPC_L_IN[28]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[28]) );
  DFFR_X1 \NPC_L_OUT_reg[27]  ( .D(NPC_L_IN[27]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[27]) );
  DFFR_X1 \NPC_L_OUT_reg[26]  ( .D(NPC_L_IN[26]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[26]) );
  DFFR_X1 \NPC_L_OUT_reg[25]  ( .D(NPC_L_IN[25]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[25]) );
  DFFR_X1 \NPC_L_OUT_reg[24]  ( .D(NPC_L_IN[24]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[24]) );
  DFFR_X1 \NPC_L_OUT_reg[23]  ( .D(NPC_L_IN[23]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[23]) );
  DFFR_X1 \NPC_L_OUT_reg[22]  ( .D(NPC_L_IN[22]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[22]) );
  DFFR_X1 \NPC_L_OUT_reg[21]  ( .D(NPC_L_IN[21]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[21]) );
  DFFR_X1 \NPC_L_OUT_reg[20]  ( .D(NPC_L_IN[20]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[20]) );
  DFFR_X1 \NPC_L_OUT_reg[19]  ( .D(NPC_L_IN[19]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[19]) );
  DFFR_X1 \NPC_L_OUT_reg[18]  ( .D(NPC_L_IN[18]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[18]) );
  DFFR_X1 \NPC_L_OUT_reg[17]  ( .D(NPC_L_IN[17]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[17]) );
  DFFR_X1 \NPC_L_OUT_reg[16]  ( .D(NPC_L_IN[16]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[16]) );
  DFFR_X1 \NPC_L_OUT_reg[15]  ( .D(NPC_L_IN[15]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[15]) );
  DFFR_X1 \NPC_L_OUT_reg[14]  ( .D(NPC_L_IN[14]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[14]) );
  DFFR_X1 \NPC_L_OUT_reg[13]  ( .D(NPC_L_IN[13]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[13]) );
  DFFR_X1 \NPC_L_OUT_reg[12]  ( .D(NPC_L_IN[12]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[12]) );
  DFFR_X1 \NPC_L_OUT_reg[11]  ( .D(NPC_L_IN[11]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[11]) );
  DFFR_X1 \NPC_L_OUT_reg[10]  ( .D(NPC_L_IN[10]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[10]) );
  DFFR_X1 \NPC_L_OUT_reg[9]  ( .D(NPC_L_IN[9]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[9]) );
  DFFR_X1 \NPC_L_OUT_reg[8]  ( .D(NPC_L_IN[8]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[8]) );
  DFFR_X1 \NPC_L_OUT_reg[7]  ( .D(NPC_L_IN[7]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[7]) );
  DFFR_X1 \NPC_L_OUT_reg[6]  ( .D(NPC_L_IN[6]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[6]) );
  DFFR_X1 \NPC_L_OUT_reg[5]  ( .D(NPC_L_IN[5]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[5]) );
  DFFR_X1 \NPC_L_OUT_reg[4]  ( .D(NPC_L_IN[4]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[4]) );
  DFFR_X1 \NPC_L_OUT_reg[3]  ( .D(NPC_L_IN[3]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[3]) );
  DFFR_X1 \NPC_L_OUT_reg[2]  ( .D(NPC_L_IN[2]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[2]) );
  DFFR_X1 \NPC_L_OUT_reg[1]  ( .D(NPC_L_IN[1]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[1]) );
  DFFR_X1 \NPC_L_OUT_reg[0]  ( .D(NPC_L_IN[0]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[0]) );
  DFFR_X1 \RS1_OUT_reg[4]  ( .D(RS1_IN[4]), .CK(CLK), .RN(n20), .Q(RS1_OUT[4])
         );
  DFFR_X1 \RS1_OUT_reg[3]  ( .D(RS1_IN[3]), .CK(CLK), .RN(n20), .Q(RS1_OUT[3])
         );
  DFFR_X1 \RS1_OUT_reg[2]  ( .D(RS1_IN[2]), .CK(CLK), .RN(n20), .Q(RS1_OUT[2])
         );
  DFFR_X1 \RS1_OUT_reg[1]  ( .D(RS1_IN[1]), .CK(CLK), .RN(n20), .Q(RS1_OUT[1])
         );
  DFFR_X1 \RS1_OUT_reg[0]  ( .D(RS1_IN[0]), .CK(CLK), .RN(n20), .Q(RS1_OUT[0])
         );
  DFFR_X1 \RS2_OUT_reg[4]  ( .D(RS2_IN[4]), .CK(CLK), .RN(n20), .Q(RS2_OUT[4])
         );
  DFFR_X1 \RS2_OUT_reg[3]  ( .D(RS2_IN[3]), .CK(CLK), .RN(n20), .Q(RS2_OUT[3])
         );
  DFFR_X1 \RS2_OUT_reg[2]  ( .D(RS2_IN[2]), .CK(CLK), .RN(n21), .Q(RS2_OUT[2])
         );
  DFFR_X1 \RS2_OUT_reg[1]  ( .D(RS2_IN[1]), .CK(CLK), .RN(n21), .Q(RS2_OUT[1])
         );
  DFFR_X1 \RS2_OUT_reg[0]  ( .D(RS2_IN[0]), .CK(CLK), .RN(n21), .Q(RS2_OUT[0])
         );
  DFFR_X1 \RD_OUT_reg[4]  ( .D(RD_IN[4]), .CK(CLK), .RN(n21), .Q(RD_OUT[4]) );
  DFFR_X1 \RD_OUT_reg[3]  ( .D(RD_IN[3]), .CK(CLK), .RN(n21), .Q(RD_OUT[3]) );
  DFFR_X1 \RD_OUT_reg[2]  ( .D(RD_IN[2]), .CK(CLK), .RN(n21), .Q(RD_OUT[2]) );
  DFFR_X1 \RD_OUT_reg[1]  ( .D(RD_IN[1]), .CK(CLK), .RN(n21), .Q(RD_OUT[1]) );
  DFFR_X1 \RD_OUT_reg[0]  ( .D(RD_IN[0]), .CK(CLK), .RN(n21), .Q(RD_OUT[0]) );
  DFFR_X1 \OPCODE_OUT_reg[5]  ( .D(OPCODE_IN[5]), .CK(CLK), .RN(n21), .Q(
        OPCODE_OUT[5]) );
  DFFR_X1 \OPCODE_OUT_reg[4]  ( .D(OPCODE_IN[4]), .CK(CLK), .RN(n21), .Q(
        OPCODE_OUT[4]) );
  DFFR_X1 \OPCODE_OUT_reg[3]  ( .D(OPCODE_IN[3]), .CK(CLK), .RN(n21), .Q(
        OPCODE_OUT[3]) );
  DFFR_X1 \OPCODE_OUT_reg[2]  ( .D(OPCODE_IN[2]), .CK(CLK), .RN(n21), .QN(n2)
         );
  DFFR_X1 \OPCODE_OUT_reg[1]  ( .D(OPCODE_IN[1]), .CK(CLK), .RN(n22), .Q(
        OPCODE_OUT[1]) );
  DFFR_X1 \OPCODE_OUT_reg[0]  ( .D(OPCODE_IN[0]), .CK(CLK), .RN(n22), .Q(
        OPCODE_OUT[0]) );
  DFFR_X1 \IR_OUT_reg[15]  ( .D(IR_IN[15]), .CK(CLK), .RN(n22), .Q(IR_OUT[15])
         );
  DFFR_X1 \IR_OUT_reg[14]  ( .D(IR_IN[14]), .CK(CLK), .RN(n22), .Q(IR_OUT[14])
         );
  DFFR_X1 \IR_OUT_reg[13]  ( .D(IR_IN[13]), .CK(CLK), .RN(n22), .Q(IR_OUT[13])
         );
  DFFR_X1 \IR_OUT_reg[12]  ( .D(IR_IN[12]), .CK(CLK), .RN(n22), .Q(IR_OUT[12])
         );
  DFFR_X1 \IR_OUT_reg[11]  ( .D(IR_IN[11]), .CK(CLK), .RN(n22), .Q(IR_OUT[11])
         );
  DFFR_X1 \IR_OUT_reg[10]  ( .D(IR_IN[10]), .CK(CLK), .RN(n22), .Q(IR_OUT[10])
         );
  DFFR_X1 \IR_OUT_reg[9]  ( .D(IR_IN[9]), .CK(CLK), .RN(n22), .Q(IR_OUT[9]) );
  DFFR_X1 \IR_OUT_reg[8]  ( .D(IR_IN[8]), .CK(CLK), .RN(n22), .Q(IR_OUT[8]) );
  DFFR_X1 \IR_OUT_reg[7]  ( .D(IR_IN[7]), .CK(CLK), .RN(n22), .Q(IR_OUT[7]) );
  DFFR_X1 \IR_OUT_reg[6]  ( .D(IR_IN[6]), .CK(CLK), .RN(n22), .Q(IR_OUT[6]) );
  DFFR_X1 \IR_OUT_reg[5]  ( .D(IR_IN[5]), .CK(CLK), .RN(n23), .Q(IR_OUT[5]) );
  DFFR_X1 \IR_OUT_reg[4]  ( .D(IR_IN[4]), .CK(CLK), .RN(n23), .Q(IR_OUT[4]) );
  DFFR_X1 \IR_OUT_reg[3]  ( .D(IR_IN[3]), .CK(CLK), .RN(n23), .Q(IR_OUT[3]) );
  DFFR_X1 \IR_OUT_reg[2]  ( .D(IR_IN[2]), .CK(CLK), .RN(n23), .Q(IR_OUT[2]) );
  DFFR_X1 \IR_OUT_reg[1]  ( .D(IR_IN[1]), .CK(CLK), .RN(n23), .Q(IR_OUT[1]) );
  DFFR_X1 \IR_OUT_reg[0]  ( .D(IR_IN[0]), .CK(CLK), .RN(n23), .Q(IR_OUT[0]) );
  INV_X1 U3 ( .A(n2), .ZN(OPCODE_OUT[2]) );
  BUF_X1 U4 ( .A(RST), .Z(n5) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n6) );
  CLKBUF_X1 U7 ( .A(n4), .Z(n7) );
  CLKBUF_X1 U8 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n4), .Z(n9) );
  CLKBUF_X1 U10 ( .A(n4), .Z(n10) );
  CLKBUF_X1 U11 ( .A(n4), .Z(n11) );
  CLKBUF_X1 U12 ( .A(n4), .Z(n12) );
  CLKBUF_X1 U13 ( .A(n5), .Z(n13) );
  CLKBUF_X1 U14 ( .A(n5), .Z(n14) );
  CLKBUF_X1 U15 ( .A(n5), .Z(n15) );
  CLKBUF_X1 U16 ( .A(n5), .Z(n16) );
  CLKBUF_X1 U17 ( .A(n5), .Z(n17) );
  CLKBUF_X1 U18 ( .A(n5), .Z(n18) );
  CLKBUF_X1 U19 ( .A(n6), .Z(n19) );
  CLKBUF_X1 U20 ( .A(n6), .Z(n20) );
  CLKBUF_X1 U21 ( .A(n6), .Z(n21) );
  CLKBUF_X1 U22 ( .A(n6), .Z(n22) );
  CLKBUF_X1 U23 ( .A(n6), .Z(n23) );
endmodule


module MUX21_GENERIC_N32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U2 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U3 ( .A(SEL), .Z(n3) );
  MUX2_X1 U4 ( .A(B[0]), .B(A[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(B[1]), .B(A[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(B[2]), .B(A[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U7 ( .A(B[3]), .B(A[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U8 ( .A(B[4]), .B(A[4]), .S(n1), .Z(Y[4]) );
  MUX2_X1 U9 ( .A(B[5]), .B(A[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(B[6]), .B(A[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(B[7]), .B(A[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(B[8]), .B(A[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(B[9]), .B(A[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(B[10]), .B(A[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(B[11]), .B(A[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(B[12]), .B(A[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(B[13]), .B(A[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(B[14]), .B(A[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(B[15]), .B(A[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(B[16]), .B(A[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(B[17]), .B(A[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(B[18]), .B(A[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(B[19]), .B(A[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(B[20]), .B(A[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(B[21]), .B(A[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(B[22]), .B(A[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(B[23]), .B(A[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(B[24]), .B(A[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(B[25]), .B(A[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(B[26]), .B(A[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(B[27]), .B(A[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(B[28]), .B(A[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(B[29]), .B(A[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(B[30]), .B(A[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(B[31]), .B(A[31]), .S(n3), .Z(Y[31]) );
endmodule


module MUX21_GENERIC_N32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  MUX2_X1 U2 ( .A(B[4]), .B(A[4]), .S(n1), .Z(Y[4]) );
  CLKBUF_X1 U3 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U4 ( .A(SEL), .Z(n3) );
  MUX2_X1 U5 ( .A(B[0]), .B(A[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(B[1]), .B(A[1]), .S(n1), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(B[2]), .B(A[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U8 ( .A(B[3]), .B(A[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U9 ( .A(B[5]), .B(A[5]), .S(n1), .Z(Y[5]) );
  MUX2_X1 U10 ( .A(B[6]), .B(A[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U11 ( .A(B[7]), .B(A[7]), .S(n1), .Z(Y[7]) );
  MUX2_X1 U12 ( .A(B[8]), .B(A[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U13 ( .A(B[9]), .B(A[9]), .S(n1), .Z(Y[9]) );
  MUX2_X1 U14 ( .A(B[10]), .B(A[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U15 ( .A(B[11]), .B(A[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U16 ( .A(B[12]), .B(A[12]), .S(n2), .Z(Y[12]) );
  MUX2_X1 U17 ( .A(B[13]), .B(A[13]), .S(n2), .Z(Y[13]) );
  MUX2_X1 U18 ( .A(B[14]), .B(A[14]), .S(n2), .Z(Y[14]) );
  MUX2_X1 U19 ( .A(B[15]), .B(A[15]), .S(n2), .Z(Y[15]) );
  MUX2_X1 U20 ( .A(B[16]), .B(A[16]), .S(n2), .Z(Y[16]) );
  MUX2_X1 U21 ( .A(B[17]), .B(A[17]), .S(n2), .Z(Y[17]) );
  MUX2_X1 U22 ( .A(B[18]), .B(A[18]), .S(n2), .Z(Y[18]) );
  MUX2_X1 U23 ( .A(B[19]), .B(A[19]), .S(n2), .Z(Y[19]) );
  MUX2_X1 U24 ( .A(B[20]), .B(A[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(B[21]), .B(A[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(B[22]), .B(A[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(B[23]), .B(A[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(B[24]), .B(A[24]), .S(n3), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(B[25]), .B(A[25]), .S(n3), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(B[26]), .B(A[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(B[27]), .B(A[27]), .S(n3), .Z(Y[27]) );
  MUX2_X1 U32 ( .A(B[28]), .B(A[28]), .S(n3), .Z(Y[28]) );
  MUX2_X1 U33 ( .A(B[29]), .B(A[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U34 ( .A(B[30]), .B(A[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U35 ( .A(B[31]), .B(A[31]), .S(n3), .Z(Y[31]) );
endmodule


module FWD_CAM_0 ( RST, DATA_IN_1, DATA_IN_2, DATA_IN_3, MATCH_1, MATCH_2, 
        MATCH_3 );
  input [5:0] DATA_IN_1;
  input [5:0] DATA_IN_2;
  input [5:0] DATA_IN_3;
  input RST;
  output MATCH_1, MATCH_2, MATCH_3;
  wire   net35857, net28092, net28091, net28089, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37;

  AND2_X1 U3 ( .A1(n29), .A2(RST), .ZN(MATCH_2) );
  AND2_X1 U4 ( .A1(DATA_IN_1[3]), .A2(DATA_IN_1[4]), .ZN(n1) );
  AND2_X1 U5 ( .A1(DATA_IN_2[3]), .A2(DATA_IN_2[4]), .ZN(n2) );
  AOI22_X1 U6 ( .A1(n5), .A2(n4), .B1(n6), .B2(n8), .ZN(n3) );
  OAI21_X1 U7 ( .B1(n3), .B2(DATA_IN_3[5]), .A(net28091), .ZN(net28089) );
  CLKBUF_X1 U8 ( .A(DATA_IN_3[3]), .Z(n8) );
  AND2_X1 U9 ( .A1(DATA_IN_3[4]), .A2(n8), .ZN(net35857) );
  OAI211_X1 U10 ( .C1(DATA_IN_3[0]), .C2(DATA_IN_3[4]), .A(DATA_IN_3[1]), .B(
        DATA_IN_3[2]), .ZN(n6) );
  AND2_X1 U11 ( .A1(DATA_IN_3[4]), .A2(DATA_IN_3[2]), .ZN(n4) );
  NAND2_X1 U12 ( .A1(n9), .A2(n10), .ZN(n5) );
  NAND2_X1 U13 ( .A1(n7), .A2(DATA_IN_3[1]), .ZN(n10) );
  INV_X1 U14 ( .A(DATA_IN_3[3]), .ZN(n7) );
  OR2_X1 U15 ( .A1(DATA_IN_3[0]), .A2(DATA_IN_3[1]), .ZN(n9) );
  XOR2_X1 U16 ( .A(DATA_IN_3[1]), .B(DATA_IN_3[2]), .Z(net28092) );
  OR2_X1 U17 ( .A1(DATA_IN_1[1]), .A2(DATA_IN_1[0]), .ZN(n16) );
  AND2_X1 U18 ( .A1(net28089), .A2(RST), .ZN(MATCH_3) );
  NAND2_X1 U19 ( .A1(net28092), .A2(net35857), .ZN(net28091) );
  NAND2_X1 U20 ( .A1(n26), .A2(n2), .ZN(n27) );
  NAND2_X1 U21 ( .A1(DATA_IN_2[1]), .A2(n12), .ZN(n13) );
  NAND2_X1 U22 ( .A1(n11), .A2(DATA_IN_2[2]), .ZN(n14) );
  NAND2_X1 U23 ( .A1(n13), .A2(n14), .ZN(n26) );
  INV_X1 U24 ( .A(DATA_IN_2[1]), .ZN(n11) );
  INV_X1 U25 ( .A(DATA_IN_2[2]), .ZN(n12) );
  AND2_X1 U26 ( .A1(DATA_IN_1[4]), .A2(DATA_IN_1[2]), .ZN(n33) );
  NAND2_X1 U27 ( .A1(n30), .A2(DATA_IN_1[1]), .ZN(n17) );
  NAND2_X1 U28 ( .A1(n16), .A2(n17), .ZN(n32) );
  INV_X1 U29 ( .A(DATA_IN_1[1]), .ZN(n15) );
  NAND2_X1 U30 ( .A1(n34), .A2(n1), .ZN(n35) );
  AND2_X1 U31 ( .A1(DATA_IN_2[4]), .A2(DATA_IN_2[2]), .ZN(n25) );
  NAND2_X1 U32 ( .A1(DATA_IN_1[1]), .A2(n18), .ZN(n19) );
  NAND2_X1 U33 ( .A1(n15), .A2(DATA_IN_1[2]), .ZN(n20) );
  NAND2_X1 U34 ( .A1(n19), .A2(n20), .ZN(n34) );
  INV_X1 U35 ( .A(DATA_IN_1[2]), .ZN(n18) );
  INV_X1 U36 ( .A(DATA_IN_2[0]), .ZN(n22) );
  INV_X1 U37 ( .A(DATA_IN_2[3]), .ZN(n21) );
  MUX2_X1 U38 ( .A(n22), .B(n21), .S(DATA_IN_2[1]), .Z(n24) );
  OAI211_X1 U39 ( .C1(DATA_IN_2[0]), .C2(DATA_IN_2[4]), .A(DATA_IN_2[1]), .B(
        DATA_IN_2[2]), .ZN(n23) );
  AOI22_X1 U40 ( .A1(n24), .A2(n25), .B1(n23), .B2(DATA_IN_2[3]), .ZN(n28) );
  OAI21_X1 U41 ( .B1(n28), .B2(DATA_IN_2[5]), .A(n27), .ZN(n29) );
  INV_X1 U42 ( .A(DATA_IN_1[3]), .ZN(n30) );
  OAI211_X1 U43 ( .C1(DATA_IN_1[0]), .C2(DATA_IN_1[4]), .A(DATA_IN_1[1]), .B(
        DATA_IN_1[2]), .ZN(n31) );
  AOI22_X1 U44 ( .A1(n33), .A2(n32), .B1(DATA_IN_1[3]), .B2(n31), .ZN(n36) );
  OAI21_X1 U45 ( .B1(n36), .B2(DATA_IN_1[5]), .A(n35), .ZN(n37) );
  AND2_X1 U46 ( .A1(n37), .A2(RST), .ZN(MATCH_1) );
endmodule


module FWD_UNIT ( Rst, Rs1, Rs2, Rd_M, Rd_W, ICODE, ICODE_M, ICODE_W, SEL_A, 
        SEL_B );
  input [4:0] Rs1;
  input [4:0] Rs2;
  input [4:0] Rd_M;
  input [4:0] Rd_W;
  input [5:0] ICODE;
  input [5:0] ICODE_M;
  input [5:0] ICODE_W;
  output [1:0] SEL_A;
  output [1:0] SEL_B;
  input Rst;
  wire   match_op, match_op_M, match_op_W, net28103, net28106, net28110,
         net28111, net28112, net28113, net28115, net28123, net28125, net28127,
         net28128, net28129, net28130, net28133, net28136, net28142, net28165,
         net28166, net28167, net28170, net29934, net35871, net37653, net35872,
         net28154, net28152, net28150, net28148, net28137, net28135, net28117,
         net28105, net28169, net28168, net28138, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54;

  FWD_CAM_0 CAM ( .RST(Rst), .DATA_IN_1(ICODE), .DATA_IN_2(ICODE_M), 
        .DATA_IN_3(ICODE_W), .MATCH_1(match_op), .MATCH_2(match_op_M), 
        .MATCH_3(match_op_W) );
  OR2_X1 U2 ( .A1(n23), .A2(net35871), .ZN(n1) );
  AND2_X1 U3 ( .A1(net28166), .A2(net28165), .ZN(n2) );
  AND2_X1 U4 ( .A1(n46), .A2(n45), .ZN(n3) );
  OR2_X1 U5 ( .A1(n1), .A2(n47), .ZN(n4) );
  NOR2_X1 U6 ( .A1(n6), .A2(net28138), .ZN(SEL_B[1]) );
  NAND4_X1 U7 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(net28138) );
  XOR2_X1 U8 ( .A(n14), .B(Rd_W[2]), .Z(n13) );
  INV_X1 U9 ( .A(Rs2[2]), .ZN(n14) );
  XOR2_X1 U10 ( .A(n15), .B(Rd_W[3]), .Z(n12) );
  INV_X1 U11 ( .A(Rs2[3]), .ZN(n15) );
  XOR2_X1 U12 ( .A(n16), .B(Rd_W[1]), .Z(n11) );
  INV_X1 U13 ( .A(Rs2[1]), .ZN(n16) );
  XOR2_X1 U14 ( .A(n16), .B(Rd_M[1]), .Z(net28166) );
  XOR2_X1 U15 ( .A(n17), .B(Rd_W[4]), .Z(n10) );
  INV_X1 U16 ( .A(Rs2[4]), .ZN(n17) );
  NAND3_X1 U17 ( .A1(n5), .A2(n8), .A3(n19), .ZN(n6) );
  AND2_X1 U18 ( .A1(net28105), .A2(n7), .ZN(n19) );
  XOR2_X1 U19 ( .A(n9), .B(Rd_W[0]), .Z(n7) );
  INV_X1 U20 ( .A(Rs2[0]), .ZN(n9) );
  XOR2_X1 U21 ( .A(n9), .B(Rd_M[0]), .Z(net28165) );
  NOR3_X1 U22 ( .A1(net35872), .A2(n18), .A3(net28106), .ZN(n8) );
  INV_X1 U23 ( .A(Rst), .ZN(n18) );
  NOR4_X1 U24 ( .A1(net28129), .A2(net28130), .A3(net35871), .A4(n18), .ZN(
        net28127) );
  NOR4_X1 U25 ( .A1(net28168), .A2(net28169), .A3(net28170), .A4(n18), .ZN(
        net28167) );
  OR2_X1 U26 ( .A1(match_op_W), .A2(net28142), .ZN(n5) );
  XOR2_X1 U27 ( .A(Rs1[2]), .B(Rd_W[2]), .Z(net28111) );
  NOR3_X1 U28 ( .A1(Rd_W[2]), .A2(Rd_W[1]), .A3(Rd_W[0]), .ZN(net28148) );
  XOR2_X1 U29 ( .A(net28137), .B(Rd_W[2]), .Z(net28150) );
  XOR2_X1 U30 ( .A(Rd_M[2]), .B(Rs2[2]), .Z(net28169) );
  INV_X1 U31 ( .A(Rd_W[3]), .ZN(net28115) );
  XOR2_X1 U32 ( .A(Rd_W[3]), .B(Rd_M[3]), .Z(net28154) );
  XOR2_X1 U33 ( .A(Rd_M[3]), .B(Rs2[3]), .Z(net28168) );
  XNOR2_X1 U34 ( .A(Rd_W[1]), .B(Rs1[1]), .ZN(net28113) );
  XOR2_X1 U35 ( .A(Rd_W[1]), .B(Rd_M[1]), .Z(net28152) );
  NAND3_X1 U36 ( .A1(n21), .A2(net28150), .A3(n20), .ZN(net28105) );
  XOR2_X1 U37 ( .A(net28135), .B(Rd_W[0]), .Z(n20) );
  INV_X1 U38 ( .A(Rd_M[0]), .ZN(net28135) );
  XOR2_X1 U39 ( .A(net28135), .B(Rs1[0]), .Z(net28123) );
  INV_X1 U40 ( .A(Rd_M[2]), .ZN(net28137) );
  NOR3_X1 U41 ( .A1(net28152), .A2(net28154), .A3(n22), .ZN(n21) );
  XOR2_X1 U42 ( .A(Rd_W[4]), .B(Rd_M[4]), .Z(n22) );
  XOR2_X1 U43 ( .A(Rs1[0]), .B(Rd_W[0]), .Z(net28110) );
  AND3_X1 U44 ( .A1(net28115), .A2(net28117), .A3(net28148), .ZN(net35872) );
  OR2_X1 U45 ( .A1(net28103), .A2(net35872), .ZN(net37653) );
  INV_X1 U46 ( .A(Rd_W[4]), .ZN(net28117) );
  XOR2_X1 U47 ( .A(net28117), .B(Rs1[4]), .Z(net28112) );
  NAND3_X1 U48 ( .A1(n26), .A2(net28127), .A3(n3), .ZN(n44) );
  INV_X1 U49 ( .A(n23), .ZN(n46) );
  NOR3_X1 U50 ( .A1(n53), .A2(net37653), .A3(n54), .ZN(SEL_A[1]) );
  XOR2_X1 U51 ( .A(Rd_M[2]), .B(Rs1[2]), .Z(n23) );
  OAI21_X1 U52 ( .B1(match_op_M), .B2(n34), .A(n33), .ZN(n24) );
  NOR2_X1 U53 ( .A1(n48), .A2(n4), .ZN(n54) );
  CLKBUF_X1 U54 ( .A(ICODE_W[0]), .Z(n25) );
  OR2_X1 U55 ( .A1(net28128), .A2(match_op), .ZN(n26) );
  NAND3_X1 U56 ( .A1(net28128), .A2(net28167), .A3(n2), .ZN(n39) );
  NOR4_X2 U57 ( .A1(n31), .A2(n30), .A3(ICODE_M[4]), .A4(ICODE_M[5]), .ZN(n34)
         );
  CLKBUF_X1 U58 ( .A(ICODE_W[1]), .Z(n27) );
  OAI21_X1 U59 ( .B1(match_op_M), .B2(n34), .A(n33), .ZN(n28) );
  OAI21_X1 U60 ( .B1(n34), .B2(match_op_M), .A(n33), .ZN(n48) );
  XNOR2_X1 U61 ( .A(Rd_M[1]), .B(Rs1[1]), .ZN(net28125) );
  OR3_X1 U62 ( .A1(ICODE_M[1]), .A2(ICODE_M[2]), .A3(ICODE_M[0]), .ZN(n31) );
  XNOR2_X1 U63 ( .A(net28133), .B(Rs1[4]), .ZN(net35871) );
  OR2_X1 U64 ( .A1(match_op), .A2(net28128), .ZN(n51) );
  OR2_X1 U65 ( .A1(net28142), .A2(match_op_W), .ZN(net29934) );
  CLKBUF_X1 U66 ( .A(ICODE_W[3]), .Z(n29) );
  CLKBUF_X1 U67 ( .A(ICODE_M[3]), .Z(n30) );
  INV_X1 U68 ( .A(Rd_M[4]), .ZN(net28133) );
  INV_X1 U69 ( .A(Rd_M[3]), .ZN(net28136) );
  NOR3_X1 U70 ( .A1(Rd_M[2]), .A2(Rd_M[0]), .A3(Rd_M[1]), .ZN(n32) );
  NAND3_X1 U71 ( .A1(net28133), .A2(net28136), .A3(n32), .ZN(n33) );
  INV_X1 U72 ( .A(ICODE[0]), .ZN(n38) );
  INV_X1 U73 ( .A(ICODE[1]), .ZN(n37) );
  INV_X1 U74 ( .A(ICODE[2]), .ZN(n36) );
  NOR3_X1 U75 ( .A1(ICODE[5]), .A2(ICODE[4]), .A3(ICODE[3]), .ZN(n35) );
  NAND4_X1 U76 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(net28106) );
  INV_X1 U77 ( .A(net28106), .ZN(net28128) );
  XOR2_X1 U78 ( .A(Rd_M[4]), .B(Rs2[4]), .Z(net28170) );
  NOR2_X1 U79 ( .A1(n28), .A2(n39), .ZN(SEL_B[0]) );
  INV_X1 U80 ( .A(ICODE_W[2]), .ZN(n42) );
  INV_X1 U81 ( .A(n27), .ZN(n41) );
  INV_X1 U82 ( .A(n25), .ZN(n40) );
  NAND3_X1 U83 ( .A1(n42), .A2(n41), .A3(n40), .ZN(n43) );
  NOR4_X1 U84 ( .A1(n43), .A2(n29), .A3(ICODE_W[4]), .A4(ICODE_W[5]), .ZN(
        net28142) );
  XOR2_X1 U85 ( .A(net28136), .B(Rs1[3]), .Z(n45) );
  INV_X1 U86 ( .A(net28123), .ZN(net28129) );
  INV_X1 U87 ( .A(net28125), .ZN(net28130) );
  NOR2_X1 U88 ( .A1(n44), .A2(n24), .ZN(SEL_A[0]) );
  NAND3_X1 U89 ( .A1(net28123), .A2(n45), .A3(net28125), .ZN(n47) );
  XOR2_X1 U90 ( .A(net28115), .B(Rs1[3]), .Z(n49) );
  NAND4_X1 U91 ( .A1(Rst), .A2(net28112), .A3(net28113), .A4(n49), .ZN(n50) );
  NOR3_X1 U92 ( .A1(n50), .A2(net28110), .A3(net28111), .ZN(n52) );
  OAI211_X1 U93 ( .C1(net28105), .C2(net28106), .A(n51), .B(n52), .ZN(n53) );
  INV_X1 U94 ( .A(net29934), .ZN(net28103) );
endmodule


module mux_3to1_N32_0 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n18, n19, n20,
         n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67;

  CLKBUF_X3 U1 ( .A(n65), .Z(n33) );
  OR3_X2 U2 ( .A1(n28), .A2(n29), .A3(n30), .ZN(Y[2]) );
  INV_X2 U3 ( .A(n59), .ZN(Y[24]) );
  NAND3_X2 U4 ( .A1(n14), .A2(n15), .A3(n16), .ZN(Y[26]) );
  BUF_X2 U5 ( .A(n65), .Z(n32) );
  OR3_X1 U6 ( .A1(n18), .A2(n19), .A3(n20), .ZN(Y[4]) );
  INV_X1 U7 ( .A(n51), .ZN(Y[16]) );
  INV_X1 U8 ( .A(n52), .ZN(Y[17]) );
  INV_X1 U9 ( .A(n53), .ZN(Y[18]) );
  INV_X1 U10 ( .A(n50), .ZN(Y[15]) );
  INV_X1 U11 ( .A(n58), .ZN(Y[23]) );
  NAND3_X1 U12 ( .A1(n7), .A2(n8), .A3(n9), .ZN(Y[3]) );
  BUF_X1 U13 ( .A(n31), .Z(n34) );
  BUF_X2 U14 ( .A(n33), .Z(n22) );
  OR3_X2 U15 ( .A1(n4), .A2(n5), .A3(n6), .ZN(Y[1]) );
  BUF_X2 U16 ( .A(n31), .Z(n21) );
  AND2_X1 U17 ( .A1(B[1]), .A2(n66), .ZN(n4) );
  AND2_X1 U18 ( .A1(A[1]), .A2(n31), .ZN(n5) );
  AND2_X1 U19 ( .A1(C[1]), .A2(n32), .ZN(n6) );
  BUF_X2 U20 ( .A(n66), .Z(n37) );
  INV_X1 U21 ( .A(n45), .ZN(Y[10]) );
  NAND2_X1 U22 ( .A1(B[3]), .A2(n36), .ZN(n7) );
  NAND2_X1 U23 ( .A1(A[3]), .A2(n21), .ZN(n8) );
  NAND2_X1 U24 ( .A1(C[3]), .A2(n33), .ZN(n9) );
  INV_X2 U25 ( .A(n44), .ZN(Y[9]) );
  NAND3_X1 U26 ( .A1(n10), .A2(n11), .A3(n12), .ZN(Y[5]) );
  NAND2_X1 U27 ( .A1(B[5]), .A2(n37), .ZN(n10) );
  NAND2_X1 U28 ( .A1(A[5]), .A2(n31), .ZN(n11) );
  NAND2_X1 U29 ( .A1(C[5]), .A2(n33), .ZN(n12) );
  INV_X2 U30 ( .A(n55), .ZN(Y[20]) );
  CLKBUF_X1 U31 ( .A(n31), .Z(n35) );
  INV_X1 U32 ( .A(n48), .ZN(Y[13]) );
  NAND2_X1 U33 ( .A1(B[26]), .A2(n37), .ZN(n14) );
  NAND2_X1 U34 ( .A1(A[26]), .A2(n21), .ZN(n15) );
  NAND2_X1 U35 ( .A1(C[26]), .A2(n32), .ZN(n16) );
  INV_X1 U36 ( .A(n47), .ZN(Y[12]) );
  INV_X1 U37 ( .A(n60), .ZN(Y[25]) );
  INV_X1 U38 ( .A(n56), .ZN(Y[21]) );
  AND2_X1 U39 ( .A1(B[4]), .A2(n66), .ZN(n18) );
  AND2_X1 U40 ( .A1(A[4]), .A2(n31), .ZN(n19) );
  AND2_X1 U41 ( .A1(C[4]), .A2(n32), .ZN(n20) );
  BUF_X2 U42 ( .A(n66), .Z(n36) );
  OR2_X1 U43 ( .A1(SEL[1]), .A2(n38), .ZN(n39) );
  INV_X1 U44 ( .A(n46), .ZN(Y[11]) );
  AND2_X2 U45 ( .A1(n40), .A2(n39), .ZN(n31) );
  INV_X2 U46 ( .A(n49), .ZN(Y[14]) );
  OR3_X2 U47 ( .A1(n26), .A2(n27), .A3(n25), .ZN(Y[0]) );
  AND2_X1 U48 ( .A1(n66), .A2(B[0]), .ZN(n25) );
  AND2_X1 U49 ( .A1(A[0]), .A2(n31), .ZN(n26) );
  AND2_X1 U50 ( .A1(C[0]), .A2(n33), .ZN(n27) );
  AND2_X1 U51 ( .A1(B[2]), .A2(n66), .ZN(n28) );
  AND2_X1 U52 ( .A1(A[2]), .A2(n31), .ZN(n29) );
  AND2_X1 U53 ( .A1(C[2]), .A2(n33), .ZN(n30) );
  INV_X2 U54 ( .A(n61), .ZN(Y[27]) );
  INV_X2 U55 ( .A(n42), .ZN(Y[7]) );
  INV_X2 U56 ( .A(n41), .ZN(Y[6]) );
  INV_X2 U57 ( .A(n57), .ZN(Y[22]) );
  INV_X2 U58 ( .A(n43), .ZN(Y[8]) );
  INV_X1 U59 ( .A(n39), .ZN(n66) );
  INV_X1 U60 ( .A(SEL[0]), .ZN(n38) );
  NAND2_X1 U61 ( .A1(n38), .A2(SEL[1]), .ZN(n40) );
  INV_X1 U62 ( .A(n40), .ZN(n65) );
  AOI222_X1 U63 ( .A1(B[6]), .A2(n36), .B1(A[6]), .B2(n31), .C1(C[6]), .C2(n33), .ZN(n41) );
  AOI222_X1 U64 ( .A1(B[7]), .A2(n37), .B1(A[7]), .B2(n35), .C1(C[7]), .C2(n32), .ZN(n42) );
  AOI222_X1 U65 ( .A1(B[8]), .A2(n36), .B1(A[8]), .B2(n31), .C1(C[8]), .C2(n32), .ZN(n43) );
  AOI222_X1 U66 ( .A1(B[9]), .A2(n36), .B1(A[9]), .B2(n21), .C1(C[9]), .C2(n32), .ZN(n44) );
  AOI222_X1 U67 ( .A1(B[10]), .A2(n36), .B1(A[10]), .B2(n21), .C1(C[10]), .C2(
        n33), .ZN(n45) );
  AOI222_X1 U68 ( .A1(B[11]), .A2(n36), .B1(A[11]), .B2(n35), .C1(C[11]), .C2(
        n22), .ZN(n46) );
  AOI222_X1 U69 ( .A1(B[12]), .A2(n36), .B1(A[12]), .B2(n21), .C1(C[12]), .C2(
        n32), .ZN(n47) );
  AOI222_X1 U70 ( .A1(B[13]), .A2(n37), .B1(A[13]), .B2(n34), .C1(C[13]), .C2(
        n22), .ZN(n48) );
  AOI222_X1 U71 ( .A1(B[14]), .A2(n36), .B1(A[14]), .B2(n21), .C1(C[14]), .C2(
        n33), .ZN(n49) );
  AOI222_X1 U72 ( .A1(B[15]), .A2(n37), .B1(A[15]), .B2(n34), .C1(C[15]), .C2(
        n22), .ZN(n50) );
  AOI222_X1 U73 ( .A1(B[16]), .A2(n37), .B1(A[16]), .B2(n35), .C1(C[16]), .C2(
        n32), .ZN(n51) );
  AOI222_X1 U74 ( .A1(B[17]), .A2(n36), .B1(A[17]), .B2(n21), .C1(C[17]), .C2(
        n22), .ZN(n52) );
  AOI222_X1 U75 ( .A1(B[18]), .A2(n36), .B1(A[18]), .B2(n34), .C1(C[18]), .C2(
        n22), .ZN(n53) );
  AOI222_X1 U76 ( .A1(B[19]), .A2(n36), .B1(A[19]), .B2(n35), .C1(C[19]), .C2(
        n33), .ZN(n54) );
  INV_X1 U77 ( .A(n54), .ZN(Y[19]) );
  AOI222_X1 U78 ( .A1(B[20]), .A2(n37), .B1(A[20]), .B2(n21), .C1(C[20]), .C2(
        n22), .ZN(n55) );
  AOI222_X1 U79 ( .A1(B[21]), .A2(n37), .B1(A[21]), .B2(n21), .C1(C[21]), .C2(
        n22), .ZN(n56) );
  AOI222_X1 U80 ( .A1(B[22]), .A2(n36), .B1(A[22]), .B2(n21), .C1(C[22]), .C2(
        n32), .ZN(n57) );
  AOI222_X1 U81 ( .A1(B[23]), .A2(n36), .B1(A[23]), .B2(n34), .C1(C[23]), .C2(
        n32), .ZN(n58) );
  AOI222_X1 U82 ( .A1(B[24]), .A2(n36), .B1(A[24]), .B2(n31), .C1(C[24]), .C2(
        n22), .ZN(n59) );
  AOI222_X1 U83 ( .A1(B[25]), .A2(n37), .B1(A[25]), .B2(n35), .C1(C[25]), .C2(
        n32), .ZN(n60) );
  AOI222_X1 U84 ( .A1(B[27]), .A2(n37), .B1(A[27]), .B2(n21), .C1(C[27]), .C2(
        n22), .ZN(n61) );
  AOI222_X1 U85 ( .A1(B[28]), .A2(n36), .B1(A[28]), .B2(n21), .C1(C[28]), .C2(
        n32), .ZN(n62) );
  INV_X1 U86 ( .A(n62), .ZN(Y[28]) );
  AOI222_X1 U87 ( .A1(B[29]), .A2(n37), .B1(A[29]), .B2(n21), .C1(C[29]), .C2(
        n33), .ZN(n63) );
  INV_X1 U88 ( .A(n63), .ZN(Y[29]) );
  AOI222_X1 U89 ( .A1(B[30]), .A2(n36), .B1(A[30]), .B2(n34), .C1(C[30]), .C2(
        n32), .ZN(n64) );
  INV_X1 U90 ( .A(n64), .ZN(Y[30]) );
  AOI222_X1 U91 ( .A1(B[31]), .A2(n36), .B1(A[31]), .B2(n34), .C1(C[31]), .C2(
        n22), .ZN(n67) );
  INV_X1 U92 ( .A(n67), .ZN(Y[31]) );
endmodule


module mux_3to1_N32_3 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   net27986, net28019, net29531, net29543, net29814, net37145, net37292,
         net37339, net37338, net37507, net37714, net37886, net37887, net37925,
         net37961, net38041, net38078, net38213, net38721, net38782, net38796,
         net39109, net43925, net28020, net45622, net37351, net37209, net28024,
         n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n28, n29, n30, n31, n32, n33, n35, n36,
         n37, n40, n41, n42, n45, n46, n47, n50, n51, n52, n54, n55, n56, n57,
         n58, n59, n62, n63, n64, n65, n66, n67, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91,
         n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105
;
  assign Y[0] = net37507;
  assign Y[14] = net37886;

  OR3_X2 U1 ( .A1(n35), .A2(n37), .A3(n36), .ZN(Y[18]) );
  NAND3_X2 U2 ( .A1(n14), .A2(n15), .A3(n16), .ZN(Y[23]) );
  CLKBUF_X1 U3 ( .A(net27986), .Z(net29543) );
  CLKBUF_X1 U4 ( .A(net27986), .Z(net37714) );
  NAND3_X1 U5 ( .A1(n54), .A2(n55), .A3(n56), .ZN(Y[22]) );
  OR3_X1 U6 ( .A1(n17), .A2(n18), .A3(n19), .ZN(Y[25]) );
  BUF_X1 U7 ( .A(net27986), .Z(net43925) );
  CLKBUF_X1 U8 ( .A(SEL[0]), .Z(net37351) );
  CLKBUF_X1 U9 ( .A(net28019), .Z(net38721) );
  OR3_X2 U10 ( .A1(n50), .A2(n51), .A3(n52), .ZN(Y[21]) );
  CLKBUF_X1 U11 ( .A(net37145), .Z(n3) );
  CLKBUF_X1 U12 ( .A(net37145), .Z(net37887) );
  NAND3_X1 U13 ( .A1(n74), .A2(n75), .A3(n76), .ZN(Y[17]) );
  NAND2_X1 U14 ( .A1(SEL[1]), .A2(n6), .ZN(net28019) );
  INV_X1 U15 ( .A(SEL[0]), .ZN(n6) );
  INV_X1 U16 ( .A(SEL[1]), .ZN(net28024) );
  NAND3_X1 U17 ( .A1(n8), .A2(n7), .A3(n9), .ZN(net37507) );
  NAND2_X1 U18 ( .A1(net27986), .A2(C[0]), .ZN(n9) );
  INV_X1 U19 ( .A(net28019), .ZN(net27986) );
  NAND2_X1 U20 ( .A1(B[0]), .A2(net29814), .ZN(n7) );
  OR2_X1 U21 ( .A1(n10), .A2(net29814), .ZN(n8) );
  NAND2_X1 U22 ( .A1(net37209), .A2(A[0]), .ZN(n10) );
  BUF_X1 U23 ( .A(net28019), .Z(net37209) );
  INV_X1 U24 ( .A(net37209), .ZN(net37292) );
  AND2_X1 U25 ( .A1(net28024), .A2(net37351), .ZN(net29814) );
  AND2_X2 U26 ( .A1(net28024), .A2(net37351), .ZN(net37925) );
  NAND2_X1 U27 ( .A1(net28024), .A2(net37351), .ZN(net28020) );
  INV_X1 U28 ( .A(net38721), .ZN(net45622) );
  INV_X1 U29 ( .A(net38721), .ZN(net38796) );
  OR3_X1 U30 ( .A1(n45), .A2(n46), .A3(n47), .ZN(Y[19]) );
  AND2_X2 U31 ( .A1(net28020), .A2(net28019), .ZN(net37145) );
  AND2_X2 U32 ( .A1(net28019), .A2(net28020), .ZN(net38041) );
  OR3_X2 U33 ( .A1(n12), .A2(n11), .A3(n13), .ZN(net37886) );
  AND2_X1 U34 ( .A1(net27986), .A2(C[14]), .ZN(n13) );
  AND2_X1 U35 ( .A1(B[14]), .A2(net29814), .ZN(n11) );
  AND2_X1 U36 ( .A1(net37145), .A2(A[14]), .ZN(n12) );
  CLKBUF_X1 U37 ( .A(net37145), .Z(net39109) );
  NAND2_X1 U38 ( .A1(B[23]), .A2(net37961), .ZN(n14) );
  NAND2_X1 U39 ( .A1(A[23]), .A2(net37887), .ZN(n15) );
  NAND2_X1 U40 ( .A1(C[23]), .A2(net37714), .ZN(n16) );
  NAND3_X1 U41 ( .A1(n71), .A2(n72), .A3(n73), .ZN(Y[13]) );
  AND2_X1 U42 ( .A1(B[25]), .A2(net37961), .ZN(n17) );
  AND2_X1 U43 ( .A1(A[25]), .A2(net37887), .ZN(n18) );
  AND2_X1 U44 ( .A1(C[25]), .A2(net29543), .ZN(n19) );
  BUF_X1 U45 ( .A(net29814), .Z(net37961) );
  NAND3_X1 U46 ( .A1(n78), .A2(n77), .A3(n79), .ZN(Y[3]) );
  NAND3_X1 U47 ( .A1(n20), .A2(n21), .A3(n22), .ZN(Y[15]) );
  NAND2_X1 U48 ( .A1(net39109), .A2(A[15]), .ZN(n20) );
  NAND2_X1 U49 ( .A1(net43925), .A2(C[15]), .ZN(n21) );
  NAND2_X1 U50 ( .A1(B[15]), .A2(net29814), .ZN(n22) );
  NAND3_X1 U51 ( .A1(n91), .A2(n90), .A3(n92), .ZN(Y[8]) );
  NAND3_X1 U52 ( .A1(n23), .A2(n24), .A3(n25), .ZN(Y[11]) );
  NAND2_X1 U53 ( .A1(net38041), .A2(A[11]), .ZN(n23) );
  NAND2_X1 U54 ( .A1(net43925), .A2(C[11]), .ZN(n24) );
  NAND2_X1 U55 ( .A1(net29814), .A2(B[11]), .ZN(n25) );
  CLKBUF_X1 U56 ( .A(net37145), .Z(net38782) );
  NAND3_X1 U57 ( .A1(n40), .A2(n41), .A3(n42), .ZN(Y[12]) );
  NAND3_X1 U58 ( .A1(n28), .A2(n29), .A3(n30), .ZN(Y[7]) );
  NAND2_X1 U59 ( .A1(net38041), .A2(A[7]), .ZN(n28) );
  NAND2_X1 U60 ( .A1(net38796), .A2(C[7]), .ZN(n29) );
  NAND2_X1 U61 ( .A1(B[7]), .A2(net37925), .ZN(n30) );
  CLKBUF_X1 U62 ( .A(net29543), .Z(net38213) );
  CLKBUF_X1 U63 ( .A(net37145), .Z(net38078) );
  NAND2_X1 U64 ( .A1(B[20]), .A2(net37961), .ZN(n31) );
  NAND2_X1 U65 ( .A1(A[20]), .A2(net38078), .ZN(n32) );
  NAND2_X1 U66 ( .A1(C[20]), .A2(net37292), .ZN(n33) );
  AND3_X1 U67 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n98) );
  CLKBUF_X1 U68 ( .A(net37925), .Z(net29531) );
  AND2_X1 U69 ( .A1(B[18]), .A2(net37925), .ZN(n35) );
  AND2_X1 U70 ( .A1(net37145), .A2(A[18]), .ZN(n36) );
  AND2_X1 U71 ( .A1(net27986), .A2(C[18]), .ZN(n37) );
  NAND3_X1 U72 ( .A1(n82), .A2(n81), .A3(n80), .ZN(Y[2]) );
  INV_X1 U73 ( .A(net37338), .ZN(net37339) );
  NAND2_X1 U74 ( .A1(B[12]), .A2(net37925), .ZN(n40) );
  NAND2_X1 U75 ( .A1(net38041), .A2(A[12]), .ZN(n41) );
  NAND2_X1 U76 ( .A1(net37292), .A2(C[12]), .ZN(n42) );
  NAND3_X1 U77 ( .A1(n87), .A2(n88), .A3(n89), .ZN(Y[10]) );
  AND2_X1 U78 ( .A1(B[19]), .A2(net37925), .ZN(n45) );
  AND2_X1 U79 ( .A1(net37145), .A2(A[19]), .ZN(n46) );
  AND2_X1 U80 ( .A1(net27986), .A2(C[19]), .ZN(n47) );
  NAND3_X1 U81 ( .A1(n57), .A2(n58), .A3(n59), .ZN(Y[4]) );
  AND2_X1 U82 ( .A1(B[21]), .A2(net37925), .ZN(n50) );
  AND2_X1 U83 ( .A1(n3), .A2(A[21]), .ZN(n51) );
  AND2_X1 U84 ( .A1(C[21]), .A2(net37292), .ZN(n52) );
  NAND3_X1 U85 ( .A1(n62), .A2(n63), .A3(n64), .ZN(Y[5]) );
  NAND2_X1 U86 ( .A1(B[22]), .A2(net37961), .ZN(n54) );
  NAND2_X1 U87 ( .A1(A[22]), .A2(net37887), .ZN(n55) );
  NAND2_X1 U88 ( .A1(C[22]), .A2(net37714), .ZN(n56) );
  NAND3_X1 U89 ( .A1(n94), .A2(n95), .A3(n96), .ZN(Y[1]) );
  NAND2_X1 U90 ( .A1(B[4]), .A2(net37925), .ZN(n57) );
  NAND2_X1 U91 ( .A1(net38041), .A2(A[4]), .ZN(n58) );
  NAND2_X1 U92 ( .A1(C[4]), .A2(net45622), .ZN(n59) );
  NAND3_X1 U93 ( .A1(n83), .A2(n84), .A3(n85), .ZN(Y[9]) );
  NAND3_X1 U94 ( .A1(n65), .A2(n66), .A3(n67), .ZN(Y[6]) );
  NAND2_X1 U95 ( .A1(net37925), .A2(B[5]), .ZN(n62) );
  NAND2_X1 U96 ( .A1(net38041), .A2(A[5]), .ZN(n63) );
  NAND2_X1 U97 ( .A1(net38796), .A2(C[5]), .ZN(n64) );
  NAND2_X1 U98 ( .A1(B[6]), .A2(net37925), .ZN(n65) );
  NAND2_X1 U99 ( .A1(net38041), .A2(A[6]), .ZN(n66) );
  NAND2_X1 U100 ( .A1(net37292), .A2(C[6]), .ZN(n67) );
  NAND2_X1 U101 ( .A1(B[13]), .A2(net37925), .ZN(n71) );
  NAND2_X1 U102 ( .A1(net38041), .A2(A[13]), .ZN(n72) );
  NAND2_X1 U103 ( .A1(C[13]), .A2(net37292), .ZN(n73) );
  NAND2_X1 U104 ( .A1(B[17]), .A2(net37925), .ZN(n74) );
  NAND2_X1 U105 ( .A1(n3), .A2(A[17]), .ZN(n75) );
  NAND2_X1 U106 ( .A1(C[17]), .A2(net38796), .ZN(n76) );
  NAND2_X1 U107 ( .A1(B[3]), .A2(net29814), .ZN(n77) );
  NAND2_X1 U108 ( .A1(net38041), .A2(A[3]), .ZN(n78) );
  NAND2_X1 U109 ( .A1(net38796), .A2(C[3]), .ZN(n79) );
  INV_X1 U110 ( .A(net38041), .ZN(net37338) );
  NAND2_X1 U111 ( .A1(net37925), .A2(B[2]), .ZN(n80) );
  NAND2_X1 U112 ( .A1(net37145), .A2(A[2]), .ZN(n81) );
  NAND2_X1 U113 ( .A1(net45622), .A2(C[2]), .ZN(n82) );
  NAND2_X1 U114 ( .A1(B[9]), .A2(net37925), .ZN(n83) );
  NAND2_X1 U115 ( .A1(net37145), .A2(A[9]), .ZN(n84) );
  NAND2_X1 U116 ( .A1(net27986), .A2(C[9]), .ZN(n85) );
  NAND2_X1 U117 ( .A1(B[10]), .A2(net37925), .ZN(n87) );
  NAND2_X1 U118 ( .A1(net38041), .A2(A[10]), .ZN(n88) );
  NAND2_X1 U119 ( .A1(C[10]), .A2(net45622), .ZN(n89) );
  NAND2_X1 U120 ( .A1(B[8]), .A2(net37925), .ZN(n90) );
  NAND2_X1 U121 ( .A1(net38041), .A2(A[8]), .ZN(n91) );
  NAND2_X1 U122 ( .A1(net37292), .A2(C[8]), .ZN(n92) );
  NAND2_X1 U123 ( .A1(B[1]), .A2(net37925), .ZN(n94) );
  NAND2_X1 U124 ( .A1(net37145), .A2(A[1]), .ZN(n95) );
  NAND2_X1 U125 ( .A1(C[1]), .A2(net27986), .ZN(n96) );
  AOI222_X1 U126 ( .A1(B[16]), .A2(net37925), .B1(net38782), .B2(A[16]), .C1(
        net37714), .C2(C[16]), .ZN(n97) );
  INV_X1 U127 ( .A(n97), .ZN(Y[16]) );
  INV_X1 U128 ( .A(n98), .ZN(Y[20]) );
  AOI222_X1 U129 ( .A1(B[24]), .A2(net29531), .B1(A[24]), .B2(net37339), .C1(
        C[24]), .C2(net29543), .ZN(n99) );
  INV_X1 U130 ( .A(n99), .ZN(Y[24]) );
  AOI222_X1 U131 ( .A1(B[26]), .A2(net37961), .B1(A[26]), .B2(net37339), .C1(
        C[26]), .C2(net29543), .ZN(n100) );
  INV_X1 U132 ( .A(n100), .ZN(Y[26]) );
  AOI222_X1 U133 ( .A1(B[27]), .A2(net29531), .B1(A[27]), .B2(net37339), .C1(
        C[27]), .C2(net29543), .ZN(n101) );
  INV_X1 U134 ( .A(n101), .ZN(Y[27]) );
  AOI222_X1 U135 ( .A1(B[28]), .A2(net29531), .B1(A[28]), .B2(net37339), .C1(
        C[28]), .C2(net29543), .ZN(n102) );
  INV_X1 U136 ( .A(n102), .ZN(Y[28]) );
  AOI222_X1 U137 ( .A1(B[29]), .A2(net29531), .B1(A[29]), .B2(net37339), .C1(
        C[29]), .C2(net38213), .ZN(n103) );
  INV_X1 U138 ( .A(n103), .ZN(Y[29]) );
  AOI222_X1 U139 ( .A1(B[30]), .A2(net29531), .B1(A[30]), .B2(net37339), .C1(
        C[30]), .C2(net29543), .ZN(n104) );
  INV_X1 U140 ( .A(n104), .ZN(Y[30]) );
  AOI222_X1 U141 ( .A1(B[31]), .A2(net29531), .B1(A[31]), .B2(net37339), .C1(
        C[31]), .C2(net38213), .ZN(n105) );
  INV_X1 U142 ( .A(n105), .ZN(Y[31]) );
endmodule


module add_sub_N32_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   net26789, net26755, net26754, net26748, net37260, net37319, net37512,
         net37522, net37543, net37600, net37602, net37633, net37685, net37702,
         net37708, net37710, net37712, net37722, net37727, net37752, net37871,
         net37882, net37954, net37922, net37353, net37243, net36877, net26708,
         net26701, net36876, net26750, net39045, net37930, net37768, net37416,
         net26732, net26707, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92;

  OR2_X1 U3 ( .A1(n10), .A2(n1), .ZN(n89) );
  NAND2_X1 U4 ( .A1(n2), .A2(net37319), .ZN(n1) );
  NOR2_X1 U5 ( .A1(net37602), .A2(net37712), .ZN(n2) );
  INV_X1 U6 ( .A(n28), .ZN(n3) );
  INV_X1 U7 ( .A(n3), .ZN(n4) );
  INV_X1 U8 ( .A(n25), .ZN(n5) );
  CLKBUF_X1 U9 ( .A(net37602), .Z(n6) );
  NOR2_X1 U10 ( .A1(n84), .A2(n85), .ZN(n7) );
  AND2_X1 U11 ( .A1(n37), .A2(n81), .ZN(n8) );
  XNOR2_X1 U12 ( .A(net37543), .B(n9), .ZN(DIFF[6]) );
  NAND2_X1 U13 ( .A1(n64), .A2(net37512), .ZN(n9) );
  OR2_X1 U14 ( .A1(n88), .A2(net26748), .ZN(n10) );
  BUF_X1 U15 ( .A(n33), .Z(net37722) );
  XNOR2_X1 U16 ( .A(n11), .B(net37954), .ZN(DIFF[11]) );
  NOR2_X1 U17 ( .A1(n60), .A2(n43), .ZN(n11) );
  CLKBUF_X1 U18 ( .A(net37243), .Z(net37416) );
  AND4_X2 U19 ( .A1(n71), .A2(n67), .A3(n70), .A4(n50), .ZN(n53) );
  XNOR2_X1 U20 ( .A(n12), .B(n81), .ZN(DIFF[26]) );
  NAND2_X1 U21 ( .A1(n46), .A2(n37), .ZN(n12) );
  AND2_X1 U22 ( .A1(net37243), .A2(n13), .ZN(n17) );
  AND2_X1 U23 ( .A1(net39045), .A2(n18), .ZN(n13) );
  NOR2_X1 U24 ( .A1(net26707), .A2(net26708), .ZN(n14) );
  XNOR2_X1 U25 ( .A(n14), .B(B[20]), .ZN(DIFF[20]) );
  INV_X1 U26 ( .A(net37768), .ZN(net26707) );
  NOR2_X1 U27 ( .A1(net37930), .A2(net26708), .ZN(net37260) );
  INV_X1 U28 ( .A(B[17]), .ZN(n16) );
  AND2_X1 U29 ( .A1(n16), .A2(n19), .ZN(n18) );
  NAND3_X1 U30 ( .A1(n19), .A2(n15), .A3(n16), .ZN(net26708) );
  INV_X1 U31 ( .A(B[19]), .ZN(n15) );
  INV_X1 U32 ( .A(B[18]), .ZN(n19) );
  AND2_X1 U33 ( .A1(net37600), .A2(net39045), .ZN(net37768) );
  CLKBUF_X1 U34 ( .A(net26732), .Z(net39045) );
  XOR2_X1 U35 ( .A(net37416), .B(net39045), .Z(DIFF[16]) );
  AND2_X1 U36 ( .A1(net37600), .A2(net39045), .ZN(net37353) );
  INV_X1 U37 ( .A(B[16]), .ZN(net26732) );
  NAND2_X1 U38 ( .A1(net26732), .A2(net26701), .ZN(net37930) );
  AND2_X1 U39 ( .A1(net26732), .A2(net37882), .ZN(net37752) );
  XNOR2_X1 U40 ( .A(n17), .B(B[19]), .ZN(DIFF[19]) );
  CLKBUF_X1 U41 ( .A(B[18]), .Z(net37922) );
  AND2_X1 U42 ( .A1(net37243), .A2(net37260), .ZN(net37727) );
  NOR2_X1 U43 ( .A1(n21), .A2(net26750), .ZN(net36876) );
  AND2_X1 U44 ( .A1(net36876), .A2(net36877), .ZN(net37600) );
  AND2_X1 U45 ( .A1(net36876), .A2(net36877), .ZN(net37243) );
  NAND4_X1 U46 ( .A1(n24), .A2(n28), .A3(n25), .A4(n20), .ZN(net26750) );
  INV_X1 U47 ( .A(B[8]), .ZN(n20) );
  NAND4_X1 U48 ( .A1(n24), .A2(n28), .A3(n25), .A4(n20), .ZN(net37602) );
  INV_X1 U49 ( .A(B[9]), .ZN(n25) );
  INV_X1 U50 ( .A(B[10]), .ZN(n28) );
  INV_X1 U51 ( .A(B[11]), .ZN(n24) );
  NAND4_X1 U52 ( .A1(n26), .A2(n27), .A3(n22), .A4(n23), .ZN(n21) );
  INV_X1 U53 ( .A(B[13]), .ZN(n23) );
  CLKBUF_X1 U54 ( .A(n23), .Z(net37633) );
  AND2_X1 U55 ( .A1(n23), .A2(net26754), .ZN(net37319) );
  INV_X1 U56 ( .A(B[12]), .ZN(n22) );
  INV_X1 U57 ( .A(B[15]), .ZN(n27) );
  INV_X1 U58 ( .A(B[14]), .ZN(n26) );
  INV_X1 U59 ( .A(B[8]), .ZN(net37702) );
  CLKBUF_X1 U60 ( .A(B[11]), .Z(net37954) );
  CLKBUF_X1 U61 ( .A(B[12]), .Z(net37712) );
  CLKBUF_X1 U62 ( .A(B[15]), .Z(net37710) );
  CLKBUF_X1 U63 ( .A(B[14]), .Z(net37708) );
  INV_X1 U64 ( .A(B[20]), .ZN(net26701) );
  NOR2_X1 U65 ( .A1(net26708), .A2(B[20]), .ZN(net37522) );
  OR2_X2 U66 ( .A1(n30), .A2(n88), .ZN(n60) );
  XNOR2_X1 U67 ( .A(n29), .B(n87), .ZN(DIFF[23]) );
  NAND2_X1 U68 ( .A1(net37243), .A2(n49), .ZN(n29) );
  XOR2_X1 U69 ( .A(n65), .B(n86), .Z(DIFF[22]) );
  NAND4_X1 U70 ( .A1(net37871), .A2(n32), .A3(n33), .A4(n31), .ZN(n30) );
  NOR2_X1 U71 ( .A1(net37685), .A2(n34), .ZN(net36877) );
  NAND4_X1 U72 ( .A1(net37871), .A2(n32), .A3(n33), .A4(n31), .ZN(n34) );
  INV_X1 U73 ( .A(B[6]), .ZN(n31) );
  NAND4_X1 U74 ( .A1(net37871), .A2(n32), .A3(n33), .A4(n31), .ZN(net26748) );
  CLKBUF_X1 U75 ( .A(n31), .Z(net37543) );
  INV_X1 U76 ( .A(B[4]), .ZN(n33) );
  INV_X1 U77 ( .A(B[5]), .ZN(n32) );
  CLKBUF_X1 U78 ( .A(n32), .Z(net37512) );
  XNOR2_X1 U79 ( .A(n35), .B(net37922), .ZN(DIFF[18]) );
  AND2_X1 U80 ( .A1(net37353), .A2(n16), .ZN(n35) );
  INV_X1 U81 ( .A(B[0]), .ZN(n36) );
  INV_X1 U82 ( .A(B[25]), .ZN(n37) );
  INV_X1 U83 ( .A(B[3]), .ZN(n38) );
  XNOR2_X1 U84 ( .A(net37708), .B(n90), .ZN(DIFF[14]) );
  OR2_X1 U85 ( .A1(net37602), .A2(net37712), .ZN(n55) );
  AND2_X2 U86 ( .A1(n53), .A2(net37722), .ZN(n64) );
  OR2_X1 U87 ( .A1(n88), .A2(net26748), .ZN(n59) );
  INV_X1 U88 ( .A(DIFF[0]), .ZN(n39) );
  INV_X1 U89 ( .A(n85), .ZN(n40) );
  NOR2_X1 U90 ( .A1(n41), .A2(n84), .ZN(n46) );
  NAND2_X1 U91 ( .A1(n83), .A2(n40), .ZN(n41) );
  OR2_X1 U92 ( .A1(n79), .A2(n42), .ZN(n76) );
  OR2_X1 U93 ( .A1(n80), .A2(B[28]), .ZN(n42) );
  OR2_X1 U94 ( .A1(n58), .A2(B[10]), .ZN(n43) );
  CLKBUF_X1 U95 ( .A(n70), .Z(n44) );
  NOR2_X1 U96 ( .A1(B[21]), .A2(B[22]), .ZN(net37882) );
  INV_X1 U97 ( .A(B[7]), .ZN(net37871) );
  INV_X1 U98 ( .A(B[21]), .ZN(n45) );
  OR2_X1 U99 ( .A1(n47), .A2(n84), .ZN(n79) );
  OR2_X1 U100 ( .A1(n85), .A2(B[24]), .ZN(n47) );
  NOR2_X1 U101 ( .A1(n60), .A2(n58), .ZN(n92) );
  NOR2_X1 U102 ( .A1(n6), .A2(n60), .ZN(n91) );
  AND2_X1 U103 ( .A1(net37522), .A2(net37752), .ZN(n49) );
  XNOR2_X1 U104 ( .A(n48), .B(n5), .ZN(DIFF[9]) );
  NOR2_X1 U105 ( .A1(n59), .A2(net26789), .ZN(n48) );
  NAND4_X1 U106 ( .A1(n77), .A2(n38), .A3(n36), .A4(n70), .ZN(net37685) );
  INV_X1 U107 ( .A(B[1]), .ZN(n50) );
  NAND2_X1 U108 ( .A1(n64), .A2(n51), .ZN(n68) );
  AND2_X1 U109 ( .A1(net37512), .A2(net37543), .ZN(n51) );
  XNOR2_X1 U110 ( .A(net37727), .B(B[21]), .ZN(DIFF[21]) );
  CLKBUF_X1 U111 ( .A(B[0]), .Z(DIFF[0]) );
  AND2_X1 U112 ( .A1(net37727), .A2(n45), .ZN(n65) );
  NOR2_X1 U113 ( .A1(n60), .A2(n55), .ZN(n54) );
  NOR2_X1 U114 ( .A1(n55), .A2(n10), .ZN(n63) );
  NOR2_X1 U115 ( .A1(n84), .A2(n85), .ZN(n56) );
  AND2_X1 U116 ( .A1(n7), .A2(n57), .ZN(n66) );
  AND2_X1 U117 ( .A1(n8), .A2(n83), .ZN(n57) );
  AND2_X1 U118 ( .A1(n63), .A2(net37633), .ZN(n90) );
  OR2_X1 U119 ( .A1(net26789), .A2(B[9]), .ZN(n58) );
  NAND2_X1 U120 ( .A1(net37600), .A2(net37260), .ZN(n84) );
  XNOR2_X1 U121 ( .A(n89), .B(net26755), .ZN(DIFF[15]) );
  INV_X1 U122 ( .A(n60), .ZN(n61) );
  XOR2_X1 U123 ( .A(n74), .B(n75), .Z(DIFF[30]) );
  NOR2_X1 U124 ( .A1(B[29]), .A2(n76), .ZN(n74) );
  NAND4_X1 U125 ( .A1(n36), .A2(n71), .A3(n50), .A4(n70), .ZN(n88) );
  NOR2_X1 U126 ( .A1(n79), .A2(n80), .ZN(n78) );
  AND2_X1 U127 ( .A1(n77), .A2(n67), .ZN(n62) );
  NAND2_X1 U128 ( .A1(n44), .A2(n62), .ZN(n69) );
  XOR2_X1 U129 ( .A(net37702), .B(n61), .Z(DIFF[8]) );
  XOR2_X1 U130 ( .A(n76), .B(B[29]), .Z(DIFF[29]) );
  XNOR2_X1 U131 ( .A(n72), .B(n73), .ZN(DIFF[31]) );
  INV_X1 U132 ( .A(B[31]), .ZN(n73) );
  NAND2_X1 U133 ( .A1(n74), .A2(n75), .ZN(n72) );
  XNOR2_X1 U134 ( .A(n78), .B(B[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U135 ( .A(n66), .B(B[27]), .ZN(DIFF[27]) );
  XOR2_X1 U136 ( .A(n44), .B(n62), .Z(DIFF[2]) );
  XOR2_X1 U137 ( .A(net37512), .B(n64), .Z(DIFF[5]) );
  XOR2_X1 U138 ( .A(n77), .B(n39), .Z(DIFF[1]) );
  INV_X1 U139 ( .A(B[2]), .ZN(n70) );
  INV_X1 U140 ( .A(net37708), .ZN(net26754) );
  XOR2_X1 U141 ( .A(n4), .B(n92), .Z(DIFF[10]) );
  INV_X1 U142 ( .A(B[26]), .ZN(n81) );
  INV_X1 U143 ( .A(B[22]), .ZN(n86) );
  INV_X1 U144 ( .A(B[3]), .ZN(n71) );
  INV_X1 U145 ( .A(B[1]), .ZN(n77) );
  INV_X1 U146 ( .A(net37710), .ZN(net26755) );
  INV_X1 U147 ( .A(B[24]), .ZN(n83) );
  INV_X1 U148 ( .A(B[30]), .ZN(n75) );
  XNOR2_X1 U149 ( .A(n56), .B(B[24]), .ZN(DIFF[24]) );
  XOR2_X1 U150 ( .A(n22), .B(n91), .Z(DIFF[12]) );
  XOR2_X1 U151 ( .A(n53), .B(net37722), .Z(DIFF[4]) );
  XOR2_X1 U152 ( .A(net37633), .B(n54), .Z(DIFF[13]) );
  XOR2_X1 U153 ( .A(n37), .B(n46), .Z(DIFF[25]) );
  XOR2_X1 U154 ( .A(net37353), .B(n16), .Z(DIFF[17]) );
  INV_X1 U155 ( .A(B[23]), .ZN(n87) );
  INV_X1 U156 ( .A(B[27]), .ZN(n82) );
  XNOR2_X1 U157 ( .A(n38), .B(n69), .ZN(DIFF[3]) );
  XNOR2_X1 U158 ( .A(net37871), .B(n68), .ZN(DIFF[7]) );
  INV_X1 U159 ( .A(B[0]), .ZN(n67) );
  NAND3_X1 U160 ( .A1(n81), .A2(n82), .A3(n37), .ZN(n80) );
  NAND3_X1 U161 ( .A1(n86), .A2(n87), .A3(n45), .ZN(n85) );
  INV_X1 U162 ( .A(net37702), .ZN(net26789) );
endmodule


module add_sub_N32 ( A, .SEL({\SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , \SEL[0] 
        }), O );
  input [31:0] A;
  output [31:0] O;
  input \SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , \SEL[0] ;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, net19775, net29489, net29487, net29485, net37049,
         net37424, net37956, net39102, net37839, net37838, n1, n2, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [4:0] SEL;
  assign O[19] = net19775;

  add_sub_N32_DW01_sub_2 sub_20 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(A), .CI(1'b0), .DIFF({N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2}) );
  NAND2_X1 U4 ( .A1(N17), .A2(n1), .ZN(n2) );
  NAND2_X2 U5 ( .A1(n25), .A2(net37838), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n2), .A2(n5), .ZN(O[15]) );
  INV_X1 U7 ( .A(net37838), .ZN(n1) );
  INV_X2 U8 ( .A(net29487), .ZN(net37838) );
  NOR4_X1 U9 ( .A1(SEL[2]), .A2(n13), .A3(SEL[4]), .A4(SEL[3]), .ZN(n15) );
  NAND2_X1 U10 ( .A1(A[17]), .A2(net37956), .ZN(n21) );
  MUX2_X1 U11 ( .A(A[13]), .B(N15), .S(net29487), .Z(O[13]) );
  MUX2_X1 U12 ( .A(A[24]), .B(N26), .S(net29489), .Z(O[24]) );
  NAND2_X1 U13 ( .A1(A[19]), .A2(net37838), .ZN(net37839) );
  CLKBUF_X1 U14 ( .A(A[5]), .Z(n6) );
  CLKBUF_X1 U15 ( .A(A[10]), .Z(n7) );
  CLKBUF_X1 U16 ( .A(A[14]), .Z(n8) );
  CLKBUF_X1 U17 ( .A(A[0]), .Z(n9) );
  INV_X1 U18 ( .A(net29489), .ZN(net37049) );
  BUF_X1 U19 ( .A(n15), .Z(net29485) );
  BUF_X1 U20 ( .A(n15), .Z(net29487) );
  INV_X1 U21 ( .A(net29489), .ZN(net37424) );
  NAND2_X1 U22 ( .A1(n28), .A2(n10), .ZN(n11) );
  NAND2_X1 U23 ( .A1(N8), .A2(net29485), .ZN(n12) );
  NAND2_X1 U24 ( .A1(n11), .A2(n12), .ZN(O[6]) );
  INV_X1 U25 ( .A(net29485), .ZN(n10) );
  MUX2_X2 U26 ( .A(A[9]), .B(N11), .S(net29485), .Z(O[9]) );
  NAND2_X1 U27 ( .A1(N21), .A2(net29487), .ZN(n16) );
  NAND2_X1 U28 ( .A1(n16), .A2(net37839), .ZN(net19775) );
  CLKBUF_X1 U29 ( .A(n15), .Z(net29489) );
  NAND2_X1 U30 ( .A1(SEL[1]), .A2(n14), .ZN(n13) );
  INV_X1 U31 ( .A(SEL[0]), .ZN(n14) );
  NAND2_X1 U32 ( .A1(N20), .A2(net29489), .ZN(n17) );
  NAND2_X1 U33 ( .A1(A[18]), .A2(net37424), .ZN(n18) );
  NAND2_X1 U34 ( .A1(n17), .A2(n18), .ZN(O[18]) );
  NAND2_X1 U35 ( .A1(A[7]), .A2(net39102), .ZN(n19) );
  NAND2_X1 U36 ( .A1(N9), .A2(net29485), .ZN(n20) );
  NAND2_X1 U37 ( .A1(n20), .A2(n19), .ZN(O[7]) );
  INV_X1 U38 ( .A(net29485), .ZN(net39102) );
  MUX2_X2 U39 ( .A(A[8]), .B(N10), .S(net29485), .Z(O[8]) );
  MUX2_X1 U40 ( .A(A[3]), .B(N5), .S(net29485), .Z(O[3]) );
  MUX2_X1 U41 ( .A(A[25]), .B(N27), .S(net29489), .Z(O[25]) );
  NAND2_X1 U42 ( .A1(N19), .A2(net29487), .ZN(n22) );
  NAND2_X1 U43 ( .A1(n21), .A2(n22), .ZN(O[17]) );
  INV_X1 U44 ( .A(net29487), .ZN(net37956) );
  MUX2_X2 U45 ( .A(A[22]), .B(N24), .S(net29487), .Z(O[22]) );
  NAND2_X1 U46 ( .A1(N29), .A2(net29489), .ZN(n23) );
  NAND2_X1 U47 ( .A1(A[27]), .A2(net37049), .ZN(n24) );
  NAND2_X1 U48 ( .A1(n23), .A2(n24), .ZN(O[27]) );
  MUX2_X2 U49 ( .A(A[23]), .B(N25), .S(net29487), .Z(O[23]) );
  MUX2_X2 U50 ( .A(n6), .B(N7), .S(net29485), .Z(O[5]) );
  CLKBUF_X1 U51 ( .A(A[15]), .Z(n25) );
  MUX2_X2 U52 ( .A(N22), .B(A[20]), .S(net37956), .Z(O[20]) );
  MUX2_X1 U53 ( .A(A[21]), .B(N23), .S(net29487), .Z(O[21]) );
  NAND2_X1 U54 ( .A1(A[11]), .A2(net37838), .ZN(n26) );
  NAND2_X1 U55 ( .A1(N13), .A2(net29485), .ZN(n27) );
  NAND2_X1 U56 ( .A1(n27), .A2(n26), .ZN(O[11]) );
  MUX2_X2 U57 ( .A(A[29]), .B(N31), .S(net29489), .Z(O[29]) );
  CLKBUF_X1 U58 ( .A(A[6]), .Z(n28) );
  NAND2_X1 U59 ( .A1(A[26]), .A2(net37424), .ZN(n29) );
  NAND2_X1 U60 ( .A1(N28), .A2(net29489), .ZN(n30) );
  NAND2_X1 U61 ( .A1(n30), .A2(n29), .ZN(O[26]) );
  MUX2_X2 U62 ( .A(A[28]), .B(N30), .S(net29489), .Z(O[28]) );
  MUX2_X2 U63 ( .A(n8), .B(N16), .S(net29487), .Z(O[14]) );
  MUX2_X1 U64 ( .A(n9), .B(N2), .S(net29485), .Z(O[0]) );
  MUX2_X1 U65 ( .A(A[1]), .B(N3), .S(net29485), .Z(O[1]) );
  MUX2_X1 U66 ( .A(A[2]), .B(N4), .S(net29485), .Z(O[2]) );
  MUX2_X1 U67 ( .A(A[4]), .B(N6), .S(net29485), .Z(O[4]) );
  MUX2_X1 U68 ( .A(n7), .B(N12), .S(net29485), .Z(O[10]) );
  MUX2_X1 U69 ( .A(A[12]), .B(N14), .S(net29487), .Z(O[12]) );
  MUX2_X1 U70 ( .A(A[16]), .B(N18), .S(net29487), .Z(O[16]) );
  MUX2_X1 U71 ( .A(A[30]), .B(N32), .S(net29489), .Z(O[30]) );
  MUX2_X1 U72 ( .A(A[31]), .B(N33), .S(net29489), .Z(O[31]) );
endmodule


module G_0 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(PA), .B2(GB), .A(GA), .ZN(n2) );
endmodule


module xor_gate_0 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_0 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_31 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_31 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_30 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_30 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_29 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_29 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_28 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_28 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_27 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_27 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_26 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_26 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_25 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_25 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_24 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_24 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_23 ( A, B, O );
  input A, B;
  output O;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(n3), .ZN(O) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module and_gate_23 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_22 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_22 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_21 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_21 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_20 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_20 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_19 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_19 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_18 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_18 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_17 ( A, B, O );
  input A, B;
  output O;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(O) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module and_gate_17 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_16 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_16 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_15 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_15 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_14 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(O) );
endmodule


module and_gate_14 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_13 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_13 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_12 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_12 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_11 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_11 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_10 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_10 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_9 ( A, B, O );
  input A, B;
  output O;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(n3), .ZN(O) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module and_gate_9 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_8 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_8 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_7 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_7 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_6 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_6 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_5 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_5 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_4 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_4 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_3 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_3 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_2 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_2 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module xor_gate_1 ( A, B, O );
  input A, B;
  output O;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(O) );
endmodule


module and_gate_1 ( A, B, O );
  input A, B;
  output O;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(O) );
endmodule


module G_9 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(PA), .B2(GB), .A(GA), .ZN(n3) );
endmodule


module PG_0 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n2;

  AND2_X1 U1 ( .A1(PB), .A2(PA), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(GB), .B2(PA), .A(GA), .ZN(n2) );
endmodule


module PG_26 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(PA), .B2(GB), .A(GA), .ZN(n3) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
endmodule


module PG_25 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(PA), .B2(GB), .A(GA), .ZN(n3) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
endmodule


module PG_24 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AND2_X1 U1 ( .A1(PB), .A2(PA), .ZN(P) );
  AOI21_X1 U2 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G) );
endmodule


module PG_23 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(PA), .B2(GB), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_22 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_21 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(PA), .B2(GB), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
endmodule


module PG_20 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_19 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_18 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net20023, net37809, n1, n2;
  assign G = net20023;
  assign net37809 = PA;

  NOR2_X1 U1 ( .A1(net37809), .A2(GA), .ZN(n2) );
  NOR2_X1 U2 ( .A1(GB), .A2(GA), .ZN(n1) );
  NOR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(net20023) );
  AND2_X1 U4 ( .A1(PB), .A2(net37809), .ZN(P) );
endmodule


module PG_17 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_16 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(PA), .B2(GB), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_15 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(PA), .B2(GB), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
endmodule


module PG_14 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  AND2_X1 U1 ( .A1(PB), .A2(PA), .ZN(P) );
  INV_X1 U2 ( .A(n3), .ZN(G) );
  AOI21_X1 U3 ( .B1(GB), .B2(PA), .A(GA), .ZN(n3) );
endmodule


module PG_13 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  AND2_X1 U1 ( .A1(PB), .A2(PA), .ZN(P) );
  INV_X1 U2 ( .A(n3), .ZN(G) );
  AOI21_X1 U3 ( .B1(GB), .B2(PA), .A(GA), .ZN(n3) );
endmodule


module G_8 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(PA), .B2(GB), .A(GA), .ZN(n3) );
endmodule


module PG_12 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n2;

  OR2_X1 U1 ( .A1(n2), .A2(GA), .ZN(G) );
  AND2_X1 U2 ( .A1(PA), .A2(GB), .ZN(n2) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
endmodule


module PG_11 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n2;

  OR2_X1 U1 ( .A1(n2), .A2(GA), .ZN(G) );
  AND2_X1 U2 ( .A1(PA), .A2(GB), .ZN(n2) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_10 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
endmodule


module PG_9 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net37216, n1, n2;
  assign G = net37216;

  NAND2_X1 U1 ( .A1(PA), .A2(GB), .ZN(n2) );
  AND2_X1 U2 ( .A1(PA), .A2(PB), .ZN(P) );
  INV_X1 U3 ( .A(GA), .ZN(n1) );
  NAND2_X1 U4 ( .A1(n2), .A2(n1), .ZN(net37216) );
endmodule


module PG_8 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net20013, n1, n2;
  assign G = net20013;

  INV_X1 U1 ( .A(GA), .ZN(n1) );
  NAND2_X1 U2 ( .A1(PA), .A2(GB), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(net20013) );
  AND2_X1 U4 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module PG_7 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net20012, n1, n2;
  assign G = net20012;

  INV_X1 U1 ( .A(GA), .ZN(n1) );
  NAND2_X1 U2 ( .A1(PA), .A2(GB), .ZN(n2) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
  NAND2_X1 U4 ( .A1(n1), .A2(n2), .ZN(net20012) );
endmodule


module PG_6 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(GB), .B2(PA), .A(GA), .ZN(n3) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module G_7 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n2;

  AND2_X1 U1 ( .A1(PA), .A2(GB), .ZN(n2) );
  OR2_X1 U2 ( .A1(n2), .A2(GA), .ZN(G) );
endmodule


module BUFF_0 ( IG, IP, OG, OP );
  input IG, IP;
  output OG, OP;
  wire   IG, IP;
  assign OG = IG;
  assign OP = IP;

endmodule


module PG_5 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net20010, n1, n2;
  assign G = net20010;

  INV_X1 U1 ( .A(GA), .ZN(n1) );
  NAND2_X1 U2 ( .A1(PA), .A2(GB), .ZN(n2) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
  NAND2_X1 U4 ( .A1(n1), .A2(n2), .ZN(net20010) );
endmodule


module BUFF_4 ( IG, IP, OG, OP );
  input IG, IP;
  output OG, OP;
  wire   IG, IP;
  assign OG = IG;
  assign OP = IP;

endmodule


module PG_4 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net20009, n1;
  assign G = net20009;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net20009) );
  AND2_X1 U3 ( .A1(PB), .A2(PA), .ZN(P) );
endmodule


module BUFF_3 ( IG, IP, OG, OP );
  input IG, IP;
  output OG, OP;
  wire   IG, IP;
  assign OG = IG;
  assign OP = IP;

endmodule


module PG_3 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  AND2_X1 U1 ( .A1(PB), .A2(PA), .ZN(P) );
  INV_X1 U2 ( .A(n3), .ZN(G) );
  AOI21_X1 U3 ( .B1(GB), .B2(PA), .A(GA), .ZN(n3) );
endmodule


module G_6 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
endmodule


module G_5 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n2;

  OR2_X2 U1 ( .A1(GA), .A2(n2), .ZN(G) );
  AND2_X1 U2 ( .A1(GB), .A2(PA), .ZN(n2) );
endmodule


module BUFF_2 ( IG, IP, OG, OP );
  input IG, IP;
  output OG, OP;
  wire   IG, IP;
  assign OG = IG;
  assign OP = IP;

endmodule


module BUFF_1 ( IG, IP, OG, OP );
  input IG, IP;
  output OG, OP;
  wire   IG, IP;
  assign OG = IG;
  assign OP = IP;

endmodule


module PG_2 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   net20007, n1, n2;
  assign G = net20007;

  NAND2_X1 U1 ( .A1(GB), .A2(PA), .ZN(n2) );
  NAND2_X1 U2 ( .A1(n2), .A2(n1), .ZN(net20007) );
  AND2_X1 U3 ( .A1(PA), .A2(PB), .ZN(P) );
  INV_X1 U4 ( .A(GA), .ZN(n1) );
endmodule


module PG_1 ( PA, PB, GA, GB, P, G );
  input PA, PB, GA, GB;
  output P, G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AND2_X1 U2 ( .A1(PB), .A2(PA), .ZN(P) );
  AOI21_X1 U3 ( .B1(GB), .B2(PA), .A(GA), .ZN(n3) );
endmodule


module G_4 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
endmodule


module G_3 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n1;

  AOI21_X1 U1 ( .B1(GB), .B2(PA), .A(GA), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G) );
endmodule


module G_2 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   net19998, n1, n2;
  assign G = net19998;

  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(net19998) );
  NAND2_X1 U2 ( .A1(GB), .A2(PA), .ZN(n2) );
  INV_X1 U3 ( .A(GA), .ZN(n1) );
endmodule


module G_1 ( PA, GA, GB, G );
  input PA, GA, GB;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(PA), .B2(GB), .A(GA), .ZN(n3) );
endmodule


module CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   n8, n9, n10, Psubtractor, Gsubtractor, \matrixG[4][31] ,
         \matrixG[4][27] , \matrixG[4][23] , \matrixG[4][19] ,
         \matrixG[3][31] , \matrixG[3][27] , \matrixG[3][23] ,
         \matrixG[3][19] , \matrixG[3][15] , \matrixG[3][11] ,
         \matrixG[2][31] , \matrixG[2][27] , \matrixG[2][23] ,
         \matrixG[2][19] , \matrixG[2][15] , \matrixG[2][11] , \matrixG[2][7] ,
         \matrixG[1][31] , \matrixG[1][29] , \matrixG[1][27] ,
         \matrixG[1][25] , \matrixG[1][23] , \matrixG[1][21] ,
         \matrixG[1][19] , \matrixG[1][17] , \matrixG[1][15] ,
         \matrixG[1][13] , \matrixG[1][11] , \matrixG[1][9] , \matrixG[1][7] ,
         \matrixG[1][5] , \matrixG[1][3] , \matrixG[1][1] , \matrixG[0][31] ,
         \matrixG[0][30] , \matrixG[0][29] , \matrixG[0][28] ,
         \matrixG[0][27] , \matrixG[0][26] , \matrixG[0][25] ,
         \matrixG[0][24] , \matrixG[0][23] , \matrixG[0][22] ,
         \matrixG[0][21] , \matrixG[0][20] , \matrixG[0][19] ,
         \matrixG[0][18] , \matrixG[0][17] , \matrixG[0][16] ,
         \matrixG[0][15] , \matrixG[0][14] , \matrixG[0][13] ,
         \matrixG[0][12] , \matrixG[0][11] , \matrixG[0][10] , \matrixG[0][9] ,
         \matrixG[0][8] , \matrixG[0][7] , \matrixG[0][6] , \matrixG[0][5] ,
         \matrixG[0][4] , \matrixG[0][3] , \matrixG[0][2] , \matrixG[0][1] ,
         \matrixG[0][0] , \matrixP[4][31] , \matrixP[4][27] , \matrixP[4][23] ,
         \matrixP[4][19] , \matrixP[3][31] , \matrixP[3][27] ,
         \matrixP[3][23] , \matrixP[3][19] , \matrixP[3][15] ,
         \matrixP[3][11] , \matrixP[2][31] , \matrixP[2][27] ,
         \matrixP[2][23] , \matrixP[2][19] , \matrixP[2][15] ,
         \matrixP[2][11] , \matrixP[2][7] , \matrixP[1][31] , \matrixP[1][29] ,
         \matrixP[1][27] , \matrixP[1][25] , \matrixP[1][23] ,
         \matrixP[1][21] , \matrixP[1][19] , \matrixP[1][17] ,
         \matrixP[1][15] , \matrixP[1][13] , \matrixP[1][11] , \matrixP[1][9] ,
         \matrixP[1][7] , \matrixP[1][5] , \matrixP[1][3] , \matrixP[0][31] ,
         \matrixP[0][30] , \matrixP[0][29] , \matrixP[0][28] ,
         \matrixP[0][27] , \matrixP[0][26] , \matrixP[0][25] ,
         \matrixP[0][24] , \matrixP[0][23] , \matrixP[0][22] ,
         \matrixP[0][21] , \matrixP[0][20] , \matrixP[0][19] ,
         \matrixP[0][18] , \matrixP[0][17] , \matrixP[0][16] ,
         \matrixP[0][15] , \matrixP[0][14] , \matrixP[0][13] ,
         \matrixP[0][12] , \matrixP[0][11] , \matrixP[0][10] , \matrixP[0][9] ,
         \matrixP[0][8] , \matrixP[0][7] , \matrixP[0][6] , \matrixP[0][5] ,
         \matrixP[0][4] , \matrixP[0][3] , \matrixP[0][2] , \matrixP[0][1] ,
         n1, n2, n5, n7;

  G_0 Gsub ( .PA(Psubtractor), .GA(Gsubtractor), .GB(Cin), .G(\matrixG[0][0] )
         );
  xor_gate_0 Xor_gsi_0_0 ( .A(A[0]), .B(B[0]), .O(Psubtractor) );
  and_gate_0 and_gsi_0_0 ( .A(A[0]), .B(B[0]), .O(Gsubtractor) );
  xor_gate_31 Xor_gsi_0_1 ( .A(A[1]), .B(B[1]), .O(\matrixP[0][1] ) );
  and_gate_31 and_gsi_0_1 ( .A(A[1]), .B(B[1]), .O(\matrixG[0][1] ) );
  xor_gate_30 Xor_gsi_0_2 ( .A(A[2]), .B(B[2]), .O(\matrixP[0][2] ) );
  and_gate_30 and_gsi_0_2 ( .A(A[2]), .B(B[2]), .O(\matrixG[0][2] ) );
  xor_gate_29 Xor_gsi_0_3 ( .A(A[3]), .B(B[3]), .O(\matrixP[0][3] ) );
  and_gate_29 and_gsi_0_3 ( .A(A[3]), .B(B[3]), .O(\matrixG[0][3] ) );
  xor_gate_28 Xor_gsi_0_4 ( .A(A[4]), .B(B[4]), .O(\matrixP[0][4] ) );
  and_gate_28 and_gsi_0_4 ( .A(A[4]), .B(B[4]), .O(\matrixG[0][4] ) );
  xor_gate_27 Xor_gsi_0_5 ( .A(A[5]), .B(B[5]), .O(\matrixP[0][5] ) );
  and_gate_27 and_gsi_0_5 ( .A(A[5]), .B(B[5]), .O(\matrixG[0][5] ) );
  xor_gate_26 Xor_gsi_0_6 ( .A(A[6]), .B(B[6]), .O(\matrixP[0][6] ) );
  and_gate_26 and_gsi_0_6 ( .A(A[6]), .B(B[6]), .O(\matrixG[0][6] ) );
  xor_gate_25 Xor_gsi_0_7 ( .A(A[7]), .B(B[7]), .O(\matrixP[0][7] ) );
  and_gate_25 and_gsi_0_7 ( .A(A[7]), .B(n1), .O(\matrixG[0][7] ) );
  xor_gate_24 Xor_gsi_0_8 ( .A(A[8]), .B(B[8]), .O(\matrixP[0][8] ) );
  and_gate_24 and_gsi_0_8 ( .A(A[8]), .B(B[8]), .O(\matrixG[0][8] ) );
  xor_gate_23 Xor_gsi_0_9 ( .A(A[9]), .B(B[9]), .O(\matrixP[0][9] ) );
  and_gate_23 and_gsi_0_9 ( .A(A[9]), .B(B[9]), .O(\matrixG[0][9] ) );
  xor_gate_22 Xor_gsi_0_10 ( .A(A[10]), .B(B[10]), .O(\matrixP[0][10] ) );
  and_gate_22 and_gsi_0_10 ( .A(A[10]), .B(B[10]), .O(\matrixG[0][10] ) );
  xor_gate_21 Xor_gsi_0_11 ( .A(A[11]), .B(B[11]), .O(\matrixP[0][11] ) );
  and_gate_21 and_gsi_0_11 ( .A(A[11]), .B(B[11]), .O(\matrixG[0][11] ) );
  xor_gate_20 Xor_gsi_0_12 ( .A(A[12]), .B(B[12]), .O(\matrixP[0][12] ) );
  and_gate_20 and_gsi_0_12 ( .A(A[12]), .B(B[12]), .O(\matrixG[0][12] ) );
  xor_gate_19 Xor_gsi_0_13 ( .A(A[13]), .B(B[13]), .O(\matrixP[0][13] ) );
  and_gate_19 and_gsi_0_13 ( .A(A[13]), .B(B[13]), .O(\matrixG[0][13] ) );
  xor_gate_18 Xor_gsi_0_14 ( .A(A[14]), .B(B[14]), .O(\matrixP[0][14] ) );
  and_gate_18 and_gsi_0_14 ( .A(A[14]), .B(B[14]), .O(\matrixG[0][14] ) );
  xor_gate_17 Xor_gsi_0_15 ( .A(A[15]), .B(B[15]), .O(\matrixP[0][15] ) );
  and_gate_17 and_gsi_0_15 ( .A(A[15]), .B(B[15]), .O(\matrixG[0][15] ) );
  xor_gate_16 Xor_gsi_0_16 ( .A(A[16]), .B(B[16]), .O(\matrixP[0][16] ) );
  and_gate_16 and_gsi_0_16 ( .A(A[16]), .B(B[16]), .O(\matrixG[0][16] ) );
  xor_gate_15 Xor_gsi_0_17 ( .A(A[17]), .B(B[17]), .O(\matrixP[0][17] ) );
  and_gate_15 and_gsi_0_17 ( .A(A[17]), .B(B[17]), .O(\matrixG[0][17] ) );
  xor_gate_14 Xor_gsi_0_18 ( .A(A[18]), .B(B[18]), .O(\matrixP[0][18] ) );
  and_gate_14 and_gsi_0_18 ( .A(A[18]), .B(B[18]), .O(\matrixG[0][18] ) );
  xor_gate_13 Xor_gsi_0_19 ( .A(A[19]), .B(B[19]), .O(\matrixP[0][19] ) );
  and_gate_13 and_gsi_0_19 ( .A(A[19]), .B(B[19]), .O(\matrixG[0][19] ) );
  xor_gate_12 Xor_gsi_0_20 ( .A(A[20]), .B(B[20]), .O(\matrixP[0][20] ) );
  and_gate_12 and_gsi_0_20 ( .A(A[20]), .B(B[20]), .O(\matrixG[0][20] ) );
  xor_gate_11 Xor_gsi_0_21 ( .A(A[21]), .B(B[21]), .O(\matrixP[0][21] ) );
  and_gate_11 and_gsi_0_21 ( .A(A[21]), .B(B[21]), .O(\matrixG[0][21] ) );
  xor_gate_10 Xor_gsi_0_22 ( .A(A[22]), .B(B[22]), .O(\matrixP[0][22] ) );
  and_gate_10 and_gsi_0_22 ( .A(A[22]), .B(B[22]), .O(\matrixG[0][22] ) );
  xor_gate_9 Xor_gsi_0_23 ( .A(A[23]), .B(B[23]), .O(\matrixP[0][23] ) );
  and_gate_9 and_gsi_0_23 ( .A(A[23]), .B(B[23]), .O(\matrixG[0][23] ) );
  xor_gate_8 Xor_gsi_0_24 ( .A(A[24]), .B(B[24]), .O(\matrixP[0][24] ) );
  and_gate_8 and_gsi_0_24 ( .A(A[24]), .B(B[24]), .O(\matrixG[0][24] ) );
  xor_gate_7 Xor_gsi_0_25 ( .A(A[25]), .B(B[25]), .O(\matrixP[0][25] ) );
  and_gate_7 and_gsi_0_25 ( .A(A[25]), .B(B[25]), .O(\matrixG[0][25] ) );
  xor_gate_6 Xor_gsi_0_26 ( .A(A[26]), .B(B[26]), .O(\matrixP[0][26] ) );
  and_gate_6 and_gsi_0_26 ( .A(A[26]), .B(B[26]), .O(\matrixG[0][26] ) );
  xor_gate_5 Xor_gsi_0_27 ( .A(A[27]), .B(B[27]), .O(\matrixP[0][27] ) );
  and_gate_5 and_gsi_0_27 ( .A(A[27]), .B(B[27]), .O(\matrixG[0][27] ) );
  xor_gate_4 Xor_gsi_0_28 ( .A(A[28]), .B(B[28]), .O(\matrixP[0][28] ) );
  and_gate_4 and_gsi_0_28 ( .A(A[28]), .B(B[28]), .O(\matrixG[0][28] ) );
  xor_gate_3 Xor_gsi_0_29 ( .A(A[29]), .B(B[29]), .O(\matrixP[0][29] ) );
  and_gate_3 and_gsi_0_29 ( .A(A[29]), .B(B[29]), .O(\matrixG[0][29] ) );
  xor_gate_2 Xor_gsi_0_30 ( .A(A[30]), .B(B[30]), .O(\matrixP[0][30] ) );
  and_gate_2 and_gsi_0_30 ( .A(A[30]), .B(B[30]), .O(\matrixG[0][30] ) );
  xor_gate_1 Xor_gsi_0_31 ( .A(A[31]), .B(B[31]), .O(\matrixP[0][31] ) );
  and_gate_1 and_gsi_0_31 ( .A(A[31]), .B(B[31]), .O(\matrixG[0][31] ) );
  G_9 Gs_d_1_1 ( .PA(\matrixP[0][1] ), .GA(\matrixG[0][1] ), .GB(
        \matrixG[0][0] ), .G(\matrixG[1][1] ) );
  PG_0 PGsi_1_3 ( .PA(\matrixP[0][3] ), .PB(\matrixP[0][2] ), .GA(
        \matrixG[0][3] ), .GB(\matrixG[0][2] ), .P(\matrixP[1][3] ), .G(
        \matrixG[1][3] ) );
  PG_26 PGsi_1_5 ( .PA(\matrixP[0][5] ), .PB(\matrixP[0][4] ), .GA(
        \matrixG[0][5] ), .GB(\matrixG[0][4] ), .P(\matrixP[1][5] ), .G(
        \matrixG[1][5] ) );
  PG_25 PGsi_1_7 ( .PA(\matrixP[0][7] ), .PB(\matrixP[0][6] ), .GA(
        \matrixG[0][7] ), .GB(\matrixG[0][6] ), .P(\matrixP[1][7] ), .G(
        \matrixG[1][7] ) );
  PG_24 PGsi_1_9 ( .PA(\matrixP[0][9] ), .PB(\matrixP[0][8] ), .GA(
        \matrixG[0][9] ), .GB(\matrixG[0][8] ), .P(\matrixP[1][9] ), .G(
        \matrixG[1][9] ) );
  PG_23 PGsi_1_11 ( .PA(\matrixP[0][11] ), .PB(\matrixP[0][10] ), .GA(
        \matrixG[0][11] ), .GB(\matrixG[0][10] ), .P(\matrixP[1][11] ), .G(
        \matrixG[1][11] ) );
  PG_22 PGsi_1_13 ( .PA(\matrixP[0][13] ), .PB(\matrixP[0][12] ), .GA(
        \matrixG[0][13] ), .GB(\matrixG[0][12] ), .P(\matrixP[1][13] ), .G(
        \matrixG[1][13] ) );
  PG_21 PGsi_1_15 ( .PA(\matrixP[0][15] ), .PB(\matrixP[0][14] ), .GA(
        \matrixG[0][15] ), .GB(\matrixG[0][14] ), .P(\matrixP[1][15] ), .G(
        \matrixG[1][15] ) );
  PG_20 PGsi_1_17 ( .PA(\matrixP[0][17] ), .PB(\matrixP[0][16] ), .GA(
        \matrixG[0][17] ), .GB(\matrixG[0][16] ), .P(\matrixP[1][17] ), .G(
        \matrixG[1][17] ) );
  PG_19 PGsi_1_19 ( .PA(\matrixP[0][19] ), .PB(\matrixP[0][18] ), .GA(
        \matrixG[0][19] ), .GB(\matrixG[0][18] ), .P(\matrixP[1][19] ), .G(
        \matrixG[1][19] ) );
  PG_18 PGsi_1_21 ( .PA(\matrixP[0][21] ), .PB(\matrixP[0][20] ), .GA(
        \matrixG[0][21] ), .GB(\matrixG[0][20] ), .P(\matrixP[1][21] ), .G(
        \matrixG[1][21] ) );
  PG_17 PGsi_1_23 ( .PA(\matrixP[0][23] ), .PB(\matrixP[0][22] ), .GA(
        \matrixG[0][23] ), .GB(\matrixG[0][22] ), .P(\matrixP[1][23] ), .G(
        \matrixG[1][23] ) );
  PG_16 PGsi_1_25 ( .PA(\matrixP[0][25] ), .PB(\matrixP[0][24] ), .GA(
        \matrixG[0][25] ), .GB(\matrixG[0][24] ), .P(\matrixP[1][25] ), .G(
        \matrixG[1][25] ) );
  PG_15 PGsi_1_27 ( .PA(\matrixP[0][27] ), .PB(\matrixP[0][26] ), .GA(
        \matrixG[0][27] ), .GB(\matrixG[0][26] ), .P(\matrixP[1][27] ), .G(
        \matrixG[1][27] ) );
  PG_14 PGsi_1_29 ( .PA(\matrixP[0][29] ), .PB(\matrixP[0][28] ), .GA(
        \matrixG[0][29] ), .GB(\matrixG[0][28] ), .P(\matrixP[1][29] ), .G(
        \matrixG[1][29] ) );
  PG_13 PGsi_1_31 ( .PA(\matrixP[0][31] ), .PB(\matrixP[0][30] ), .GA(
        \matrixG[0][31] ), .GB(\matrixG[0][30] ), .P(\matrixP[1][31] ), .G(
        \matrixG[1][31] ) );
  G_8 Gs_d_2_3 ( .PA(\matrixP[1][3] ), .GA(\matrixG[1][3] ), .GB(
        \matrixG[1][1] ), .G(n10) );
  PG_12 PGsi_2_7 ( .PA(\matrixP[1][7] ), .PB(\matrixP[1][5] ), .GA(
        \matrixG[1][7] ), .GB(\matrixG[1][5] ), .P(\matrixP[2][7] ), .G(
        \matrixG[2][7] ) );
  PG_11 PGsi_2_11 ( .PA(\matrixP[1][11] ), .PB(\matrixP[1][9] ), .GA(
        \matrixG[1][11] ), .GB(\matrixG[1][9] ), .P(\matrixP[2][11] ), .G(
        \matrixG[2][11] ) );
  PG_10 PGsi_2_15 ( .PA(\matrixP[1][15] ), .PB(\matrixP[1][13] ), .GA(
        \matrixG[1][15] ), .GB(\matrixG[1][13] ), .P(\matrixP[2][15] ), .G(
        \matrixG[2][15] ) );
  PG_9 PGsi_2_19 ( .PA(\matrixP[1][19] ), .PB(\matrixP[1][17] ), .GA(
        \matrixG[1][19] ), .GB(\matrixG[1][17] ), .P(\matrixP[2][19] ), .G(
        \matrixG[2][19] ) );
  PG_8 PGsi_2_23 ( .PA(\matrixP[1][23] ), .PB(\matrixP[1][21] ), .GA(
        \matrixG[1][23] ), .GB(\matrixG[1][21] ), .P(\matrixP[2][23] ), .G(
        \matrixG[2][23] ) );
  PG_7 PGsi_2_27 ( .PA(\matrixP[1][27] ), .PB(\matrixP[1][25] ), .GA(
        \matrixG[1][27] ), .GB(\matrixG[1][25] ), .P(\matrixP[2][27] ), .G(
        \matrixG[2][27] ) );
  PG_6 PGsi_2_31 ( .PA(\matrixP[1][31] ), .PB(\matrixP[1][29] ), .GA(
        \matrixG[1][31] ), .GB(\matrixG[1][29] ), .P(\matrixP[2][31] ), .G(
        \matrixG[2][31] ) );
  G_7 Gs_h_3_7 ( .PA(\matrixP[2][7] ), .GA(\matrixG[2][7] ), .GB(n10), .G(n9)
         );
  BUFF_0 Buf_h_3_11 ( .IG(\matrixG[2][11] ), .IP(\matrixP[2][11] ), .OG(
        \matrixG[3][11] ), .OP(\matrixP[3][11] ) );
  PG_5 PGsi_3_15 ( .PA(\matrixP[2][15] ), .PB(\matrixP[3][11] ), .GA(
        \matrixG[2][15] ), .GB(\matrixG[2][11] ), .P(\matrixP[3][15] ), .G(
        \matrixG[3][15] ) );
  BUFF_4 Buf_h_3_19 ( .IG(n2), .IP(\matrixP[2][19] ), .OG(\matrixG[3][19] ), 
        .OP(\matrixP[3][19] ) );
  PG_4 PGsi_3_23 ( .PA(\matrixP[2][23] ), .PB(\matrixP[3][19] ), .GA(
        \matrixG[2][23] ), .GB(\matrixG[2][19] ), .P(\matrixP[3][23] ), .G(
        \matrixG[3][23] ) );
  BUFF_3 Buf_h_3_27 ( .IG(\matrixG[2][27] ), .IP(\matrixP[2][27] ), .OG(
        \matrixG[3][27] ), .OP(\matrixP[3][27] ) );
  PG_3 PGsi_3_31 ( .PA(\matrixP[2][31] ), .PB(\matrixP[3][27] ), .GA(
        \matrixG[2][31] ), .GB(\matrixG[2][27] ), .P(\matrixP[3][31] ), .G(
        \matrixG[3][31] ) );
  G_6 Gs_h_4_11 ( .PA(\matrixP[3][11] ), .GA(\matrixG[3][11] ), .GB(Co[1]), 
        .G(Co[2]) );
  G_5 Gs_h_4_15 ( .PA(\matrixP[3][15] ), .GA(\matrixG[3][15] ), .GB(n9), .G(n8) );
  BUFF_2 Buf_h_4_19_0 ( .IG(\matrixG[3][19] ), .IP(\matrixP[3][19] ), .OG(
        \matrixG[4][19] ), .OP(\matrixP[4][19] ) );
  BUFF_1 Buf_h_4_23_0 ( .IG(n7), .IP(\matrixP[3][23] ), .OG(\matrixG[4][23] ), 
        .OP(\matrixP[4][23] ) );
  PG_2 PGsi_4_27_0 ( .PA(\matrixP[3][27] ), .PB(\matrixP[3][23] ), .GA(
        \matrixG[3][27] ), .GB(\matrixG[3][23] ), .P(\matrixP[4][27] ), .G(
        \matrixG[4][27] ) );
  PG_1 PGsi_4_31_0 ( .PA(\matrixP[3][31] ), .PB(\matrixP[3][23] ), .GA(
        \matrixG[3][31] ), .GB(n7), .P(\matrixP[4][31] ), .G(\matrixG[4][31] )
         );
  G_4 Gs_h_5_19 ( .PA(\matrixP[4][19] ), .GA(\matrixG[4][19] ), .GB(n8), .G(
        Co[4]) );
  G_3 Gs_h_5_23 ( .PA(\matrixP[4][23] ), .GA(\matrixG[4][23] ), .GB(n8), .G(
        Co[5]) );
  G_2 Gs_h_5_27 ( .PA(\matrixP[4][27] ), .GA(\matrixG[4][27] ), .GB(n8), .G(
        Co[6]) );
  G_1 Gs_h_5_31 ( .PA(\matrixP[4][31] ), .GA(\matrixG[4][31] ), .GB(Co[3]), 
        .G(Co[7]) );
  INV_X2 U1 ( .A(n5), .ZN(Co[3]) );
  CLKBUF_X1 U2 ( .A(B[7]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(\matrixG[2][19] ), .Z(n2) );
  BUF_X1 U4 ( .A(\matrixG[3][23] ), .Z(n7) );
  CLKBUF_X1 U5 ( .A(n9), .Z(Co[1]) );
  CLKBUF_X1 U6 ( .A(n10), .Z(Co[0]) );
  INV_X1 U7 ( .A(n8), .ZN(n5) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n5;

  INV_X1 U1 ( .A(n8), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n5), .ZN(n8) );
  INV_X1 U3 ( .A(n7), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n5), .ZN(n7) );
  INV_X1 U5 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U6 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n6) );
  INV_X1 U7 ( .A(n9), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n5), .ZN(n9) );
  INV_X1 U9 ( .A(SEL), .ZN(n5) );
endmodule


module carry_select_block_N4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_0 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_15 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_0 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n5, n10, n11, n12, n13;

  INV_X1 U1 ( .A(SEL), .ZN(n5) );
  INV_X1 U2 ( .A(n13), .ZN(Y[3]) );
  AOI22_X1 U3 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n13) );
  INV_X1 U4 ( .A(n12), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n5), .ZN(n12) );
  INV_X1 U6 ( .A(n11), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n5), .ZN(n11) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n5), .ZN(n10) );
endmodule


module carry_select_block_N4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_14 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_13 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_7 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n1) );
  INV_X1 U2 ( .A(n5), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n1), .A2(n9), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n1) );
  INV_X1 U6 ( .A(n9), .ZN(n4) );
  INV_X1 U7 ( .A(n8), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(Ci), .ZN(n8) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n5, n10, n11, n12, n13;

  INV_X1 U1 ( .A(SEL), .ZN(n5) );
  INV_X1 U2 ( .A(n12), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n5), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n5), .ZN(n13) );
  INV_X1 U6 ( .A(n11), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n5), .ZN(n11) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n5), .ZN(n10) );
endmodule


module carry_select_block_N4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_12 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_11 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_6 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(B[0]), .B(A[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(B[1]), .B(A[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(B[3]), .B(A[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_10 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_9 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_5 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(B[0]), .B(A[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(B[1]), .B(A[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(B[3]), .B(A[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_8 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_7 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_4 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5, n6;

  INV_X1 U1 ( .A(n3), .ZN(n1) );
  XNOR2_X1 U2 ( .A(A), .B(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n2), .ZN(S) );
  INV_X1 U5 ( .A(A), .ZN(n4) );
  INV_X1 U6 ( .A(Ci), .ZN(n5) );
  INV_X1 U7 ( .A(B), .ZN(n3) );
  OAI22_X1 U8 ( .A1(n6), .A2(n5), .B1(n4), .B2(n3), .ZN(Co) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n3), .A2(n4), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5, n6;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n1) );
  INV_X1 U2 ( .A(A), .ZN(n3) );
  XOR2_X1 U3 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U4 ( .A(Ci), .ZN(n4) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n5), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
  INV_X1 U7 ( .A(n5), .ZN(n6) );
  XOR2_X1 U8 ( .A(n1), .B(n6), .Z(S) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n5), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n1) );
  INV_X1 U3 ( .A(A), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U5 ( .A(n1), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n2) );
  OAI22_X1 U7 ( .A1(n5), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(n4), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(S) );
  INV_X1 U3 ( .A(A), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n2) );
  OAI22_X1 U7 ( .A1(n5), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U2 ( .A(B[3]), .B(A[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U3 ( .A(B[0]), .B(A[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(B[1]), .B(A[1]), .S(SEL), .Z(Y[1]) );
endmodule


module carry_select_block_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_6 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_5 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_3 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n4) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U3 ( .A(A), .ZN(n2) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(B[3]), .B(A[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U3 ( .A(B[0]), .B(A[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(B[1]), .B(A[1]), .S(SEL), .Z(Y[1]) );
endmodule


module carry_select_block_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_4 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_3 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_2 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n5) );
  XNOR2_X1 U3 ( .A(Ci), .B(n5), .ZN(S) );
  INV_X1 U4 ( .A(A), .ZN(n3) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n2) );
  OAI22_X1 U7 ( .A1(n1), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(n4), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(S) );
  INV_X1 U3 ( .A(A), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n2) );
  OAI22_X1 U7 ( .A1(n5), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5, n6;

  INV_X1 U1 ( .A(n4), .ZN(n1) );
  INV_X1 U2 ( .A(A), .ZN(n3) );
  XOR2_X1 U3 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U4 ( .A(Ci), .ZN(n4) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n4), .A2(n5), .B1(n3), .B2(n2), .ZN(Co) );
  INV_X1 U7 ( .A(n5), .ZN(n6) );
  XOR2_X1 U8 ( .A(n6), .B(n1), .Z(S) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n5), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n1) );
  INV_X1 U3 ( .A(A), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U5 ( .A(n1), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n2) );
  OAI22_X1 U7 ( .A1(n5), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  XOR2_X1 U2 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U3 ( .A(Ci), .ZN(n3) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  OAI22_X1 U5 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
  XOR2_X1 U7 ( .A(Ci), .B(n5), .Z(S) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(n4), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(S) );
  INV_X1 U3 ( .A(A), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(B), .Z(n5) );
  INV_X1 U5 ( .A(Ci), .ZN(n4) );
  INV_X1 U6 ( .A(B), .ZN(n2) );
  OAI22_X1 U7 ( .A1(n5), .A2(n4), .B1(n3), .B2(n2), .ZN(Co) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  XOR2_X1 U3 ( .A(n2), .B(B), .Z(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3;

  NAND2_X1 U1 ( .A1(n1), .A2(B[3]), .ZN(n2) );
  NAND2_X1 U2 ( .A1(SEL), .A2(A[3]), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(Y[3]) );
  INV_X1 U4 ( .A(SEL), .ZN(n1) );
  MUX2_X1 U5 ( .A(B[0]), .B(A[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(B[1]), .B(A[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(B[2]), .B(A[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_N4_2 RCA0 ( .A(A), .B(B), .Ci(1'b1), .S(S0) );
  RCA_N4_1 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  MUX21_GENERIC_N4_1 MUXSUM ( .A(S0), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Cin, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Cin;
  output [31:0] S;


  carry_select_block_N4_0 BLI_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Cin[0]), .S(
        S[3:0]) );
  carry_select_block_N4_7 BLI_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Cin[1]), .S(
        S[7:4]) );
  carry_select_block_N4_6 BLI_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Cin[2]), .S(
        S[11:8]) );
  carry_select_block_N4_5 BLI_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Cin[3]), .S(
        S[15:12]) );
  carry_select_block_N4_4 BLI_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Cin[4]), .S(
        S[19:16]) );
  carry_select_block_N4_3 BLI_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Cin[5]), .S(
        S[23:20]) );
  carry_select_block_N4_2 BLI_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Cin[6]), .S(
        S[27:24]) );
  carry_select_block_N4_1 BLI_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Cin[7]), .S(
        S[31:28]) );
endmodule


module P4_ADDER_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;
  wire   [6:0] carryv;

  CARRY_GENERATOR_PARAMETRIC_NBIT32_NBIT_PER_BLOCK4 C_GEN ( .A(A), .B({
        B[31:30], n1, n5, B[27:0]}), .Cin(Cin), .Co({Cout, carryv}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 S_GEN ( .A(A), .B({B[31:28], n12, n21, 
        n18, B[24], n19, n17, n11, n14, n20, n9, n13, B[16], n16, B[14:12], n6, 
        B[10], n8, B[8], n15, n4, n2, B[4], n3, B[2:0]}), .Cin({carryv, Cin}), 
        .S(S) );
  BUF_X1 U1 ( .A(B[20]), .Z(n14) );
  CLKBUF_X1 U2 ( .A(B[29]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(B[5]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(B[3]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[6]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(B[28]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[25]), .Z(n18) );
  CLKBUF_X1 U8 ( .A(B[11]), .Z(n6) );
  INV_X1 U9 ( .A(B[9]), .ZN(n7) );
  INV_X1 U10 ( .A(n7), .ZN(n8) );
  CLKBUF_X1 U11 ( .A(B[18]), .Z(n9) );
  INV_X1 U12 ( .A(B[21]), .ZN(n10) );
  INV_X1 U13 ( .A(n10), .ZN(n11) );
  CLKBUF_X1 U14 ( .A(B[27]), .Z(n12) );
  CLKBUF_X1 U15 ( .A(B[17]), .Z(n13) );
  CLKBUF_X1 U16 ( .A(B[7]), .Z(n15) );
  CLKBUF_X1 U17 ( .A(B[15]), .Z(n16) );
  CLKBUF_X1 U18 ( .A(B[22]), .Z(n17) );
  CLKBUF_X1 U19 ( .A(B[23]), .Z(n19) );
  CLKBUF_X1 U20 ( .A(B[19]), .Z(n20) );
  CLKBUF_X1 U21 ( .A(B[26]), .Z(n21) );
endmodule


module add_wrapper_N32 ( A, B, .SEL({\SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , 
        \SEL[0] }), O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  input \SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , \SEL[0] ;

  wire   [4:0] SEL;
  wire   [31:0] outp;

  add_sub_N32 sign ( .A(B), .SEL({\SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , 
        \SEL[0] }), .O(outp) );
  P4_ADDER_NBIT32 adder ( .A(A), .B(outp), .Cin(1'b0), .S(O) );
endmodule


module logic_N32 ( A, B, .SEL({\SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , 
        \SEL[0] }), O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  input \SEL[4] , \SEL[3] , \SEL[2] , \SEL[1] , \SEL[0] ;
  wire   n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n69, n135, n136, n137, n138, n139, n140, n141, n142;
  wire   [4:0] SEL;

  INV_X1 U2 ( .A(SEL[2]), .ZN(n142) );
  AOI22_X1 U3 ( .A1(n8), .A2(n16), .B1(A[0]), .B2(n2), .ZN(n132) );
  AOI22_X1 U4 ( .A1(n9), .A2(n41), .B1(A[3]), .B2(n4), .ZN(n82) );
  AOI21_X1 U5 ( .B1(n10), .B2(n11), .A(n5), .ZN(n133) );
  AOI21_X1 U6 ( .B1(n10), .B2(n12), .A(n5), .ZN(n111) );
  AOI21_X1 U7 ( .B1(n9), .B2(n13), .A(n6), .ZN(n89) );
  AOI21_X1 U8 ( .B1(n8), .B2(n14), .A(n7), .ZN(n83) );
  INV_X1 U9 ( .A(A[3]), .ZN(n41) );
  INV_X1 U10 ( .A(A[0]), .ZN(n16) );
  INV_X1 U11 ( .A(n1), .ZN(n10) );
  BUF_X1 U12 ( .A(n70), .Z(n5) );
  BUF_X1 U13 ( .A(n70), .Z(n6) );
  OAI22_X1 U14 ( .A1(n116), .A2(n55), .B1(n117), .B2(n24), .ZN(O[17]) );
  AOI21_X1 U15 ( .B1(n10), .B2(n55), .A(n5), .ZN(n117) );
  AOI22_X1 U16 ( .A1(n9), .A2(n24), .B1(A[17]), .B2(n2), .ZN(n116) );
  INV_X1 U17 ( .A(B[17]), .ZN(n55) );
  OAI22_X1 U18 ( .A1(n106), .A2(n59), .B1(n107), .B2(n29), .ZN(O[21]) );
  AOI21_X1 U19 ( .B1(n10), .B2(n59), .A(n6), .ZN(n107) );
  AOI22_X1 U20 ( .A1(n9), .A2(n29), .B1(A[21]), .B2(n3), .ZN(n106) );
  INV_X1 U21 ( .A(B[21]), .ZN(n59) );
  OAI22_X1 U22 ( .A1(n80), .A2(n15), .B1(n81), .B2(n42), .ZN(O[4]) );
  AOI21_X1 U23 ( .B1(n9), .B2(n15), .A(n7), .ZN(n81) );
  OAI22_X1 U24 ( .A1(n78), .A2(n137), .B1(n79), .B2(n43), .ZN(O[5]) );
  AOI21_X1 U25 ( .B1(n8), .B2(n137), .A(n7), .ZN(n79) );
  INV_X1 U26 ( .A(B[5]), .ZN(n137) );
  OAI22_X1 U27 ( .A1(n74), .A2(n139), .B1(n75), .B2(n45), .ZN(O[7]) );
  AOI21_X1 U28 ( .B1(n8), .B2(n139), .A(n7), .ZN(n75) );
  AOI22_X1 U29 ( .A1(n8), .A2(n45), .B1(A[7]), .B2(n4), .ZN(n74) );
  INV_X1 U30 ( .A(B[7]), .ZN(n139) );
  OAI22_X1 U31 ( .A1(n76), .A2(n138), .B1(n77), .B2(n44), .ZN(O[6]) );
  AOI21_X1 U32 ( .B1(n8), .B2(n138), .A(n7), .ZN(n77) );
  AOI22_X1 U33 ( .A1(n8), .A2(n44), .B1(A[6]), .B2(n4), .ZN(n76) );
  INV_X1 U34 ( .A(B[6]), .ZN(n138) );
  OAI22_X1 U35 ( .A1(n67), .A2(n141), .B1(n68), .B2(n47), .ZN(O[9]) );
  AOI21_X1 U36 ( .B1(n9), .B2(n141), .A(n7), .ZN(n68) );
  AOI22_X1 U37 ( .A1(n8), .A2(n47), .B1(n4), .B2(A[9]), .ZN(n67) );
  INV_X1 U38 ( .A(B[9]), .ZN(n141) );
  OAI22_X1 U39 ( .A1(n72), .A2(n140), .B1(n73), .B2(n46), .ZN(O[8]) );
  AOI21_X1 U40 ( .B1(n8), .B2(n140), .A(n7), .ZN(n73) );
  AOI22_X1 U41 ( .A1(n8), .A2(n46), .B1(A[8]), .B2(n4), .ZN(n72) );
  INV_X1 U42 ( .A(B[8]), .ZN(n140) );
  OAI22_X1 U43 ( .A1(n130), .A2(n48), .B1(n131), .B2(n17), .ZN(O[10]) );
  AOI21_X1 U44 ( .B1(n8), .B2(n48), .A(n5), .ZN(n131) );
  AOI22_X1 U45 ( .A1(n8), .A2(n17), .B1(A[10]), .B2(n2), .ZN(n130) );
  INV_X1 U46 ( .A(B[10]), .ZN(n48) );
  OAI22_X1 U47 ( .A1(n128), .A2(n49), .B1(n129), .B2(n18), .ZN(O[11]) );
  AOI21_X1 U48 ( .B1(n9), .B2(n49), .A(n5), .ZN(n129) );
  AOI22_X1 U49 ( .A1(n8), .A2(n18), .B1(A[11]), .B2(n2), .ZN(n128) );
  INV_X1 U50 ( .A(B[11]), .ZN(n49) );
  OAI22_X1 U51 ( .A1(n112), .A2(n57), .B1(n113), .B2(n26), .ZN(O[19]) );
  AOI21_X1 U52 ( .B1(n10), .B2(n57), .A(n5), .ZN(n113) );
  AOI22_X1 U53 ( .A1(n9), .A2(n26), .B1(A[19]), .B2(n2), .ZN(n112) );
  INV_X1 U54 ( .A(B[19]), .ZN(n57) );
  OAI22_X1 U55 ( .A1(n108), .A2(n58), .B1(n109), .B2(n28), .ZN(O[20]) );
  AOI21_X1 U56 ( .B1(n10), .B2(n58), .A(n6), .ZN(n109) );
  AOI22_X1 U57 ( .A1(n9), .A2(n28), .B1(A[20]), .B2(n3), .ZN(n108) );
  INV_X1 U58 ( .A(B[20]), .ZN(n58) );
  BUF_X1 U59 ( .A(n71), .Z(n2) );
  BUF_X1 U60 ( .A(n71), .Z(n3) );
  OAI22_X1 U61 ( .A1(n86), .A2(n135), .B1(n87), .B2(n39), .ZN(O[30]) );
  AOI21_X1 U62 ( .B1(n8), .B2(n135), .A(n6), .ZN(n87) );
  AOI22_X1 U63 ( .A1(n9), .A2(n39), .B1(A[30]), .B2(n3), .ZN(n86) );
  INV_X1 U64 ( .A(B[30]), .ZN(n135) );
  INV_X1 U65 ( .A(A[7]), .ZN(n45) );
  OAI22_X1 U66 ( .A1(n102), .A2(n61), .B1(n103), .B2(n31), .ZN(O[23]) );
  AOI21_X1 U67 ( .B1(n10), .B2(n61), .A(n6), .ZN(n103) );
  AOI22_X1 U68 ( .A1(n9), .A2(n31), .B1(A[23]), .B2(n3), .ZN(n102) );
  INV_X1 U69 ( .A(B[23]), .ZN(n61) );
  OAI22_X1 U70 ( .A1(n126), .A2(n50), .B1(n127), .B2(n19), .ZN(O[12]) );
  AOI21_X1 U71 ( .B1(n10), .B2(n50), .A(n5), .ZN(n127) );
  AOI22_X1 U72 ( .A1(n8), .A2(n19), .B1(A[12]), .B2(n2), .ZN(n126) );
  INV_X1 U73 ( .A(B[12]), .ZN(n50) );
  OAI22_X1 U74 ( .A1(n122), .A2(n52), .B1(n123), .B2(n21), .ZN(O[14]) );
  AOI21_X1 U75 ( .B1(n10), .B2(n52), .A(n5), .ZN(n123) );
  AOI22_X1 U76 ( .A1(n8), .A2(n21), .B1(A[14]), .B2(n2), .ZN(n122) );
  INV_X1 U77 ( .A(B[14]), .ZN(n52) );
  OAI22_X1 U78 ( .A1(n124), .A2(n51), .B1(n125), .B2(n20), .ZN(O[13]) );
  AOI21_X1 U79 ( .B1(n8), .B2(n51), .A(n5), .ZN(n125) );
  AOI22_X1 U80 ( .A1(n8), .A2(n20), .B1(A[13]), .B2(n2), .ZN(n124) );
  INV_X1 U81 ( .A(B[13]), .ZN(n51) );
  OAI22_X1 U82 ( .A1(n120), .A2(n53), .B1(n121), .B2(n22), .ZN(O[15]) );
  AOI21_X1 U83 ( .B1(n10), .B2(n53), .A(n5), .ZN(n121) );
  AOI22_X1 U84 ( .A1(n8), .A2(n22), .B1(A[15]), .B2(n2), .ZN(n120) );
  INV_X1 U85 ( .A(B[15]), .ZN(n53) );
  OAI22_X1 U86 ( .A1(n118), .A2(n54), .B1(n119), .B2(n23), .ZN(O[16]) );
  AOI21_X1 U87 ( .B1(n10), .B2(n54), .A(n5), .ZN(n119) );
  AOI22_X1 U88 ( .A1(n8), .A2(n23), .B1(A[16]), .B2(n2), .ZN(n118) );
  INV_X1 U89 ( .A(B[16]), .ZN(n54) );
  OAI22_X1 U90 ( .A1(n94), .A2(n65), .B1(n95), .B2(n35), .ZN(O[27]) );
  AOI21_X1 U91 ( .B1(n10), .B2(n65), .A(n6), .ZN(n95) );
  AOI22_X1 U92 ( .A1(n10), .A2(n35), .B1(A[27]), .B2(n3), .ZN(n94) );
  INV_X1 U93 ( .A(B[27]), .ZN(n65) );
  OAI22_X1 U94 ( .A1(n96), .A2(n64), .B1(n97), .B2(n34), .ZN(O[26]) );
  AOI21_X1 U95 ( .B1(n8), .B2(n64), .A(n6), .ZN(n97) );
  AOI22_X1 U96 ( .A1(n9), .A2(n34), .B1(A[26]), .B2(n3), .ZN(n96) );
  INV_X1 U97 ( .A(B[26]), .ZN(n64) );
  OAI22_X1 U98 ( .A1(n84), .A2(n136), .B1(n85), .B2(n40), .ZN(O[31]) );
  AOI21_X1 U99 ( .B1(n9), .B2(n136), .A(n7), .ZN(n85) );
  AOI22_X1 U100 ( .A1(n8), .A2(n40), .B1(A[31]), .B2(n4), .ZN(n84) );
  INV_X1 U101 ( .A(B[31]), .ZN(n136) );
  OAI22_X1 U102 ( .A1(n92), .A2(n66), .B1(n93), .B2(n36), .ZN(O[28]) );
  AOI21_X1 U103 ( .B1(n10), .B2(n66), .A(n6), .ZN(n93) );
  AOI22_X1 U104 ( .A1(n9), .A2(n36), .B1(A[28]), .B2(n3), .ZN(n92) );
  INV_X1 U105 ( .A(B[28]), .ZN(n66) );
  OAI22_X1 U106 ( .A1(n114), .A2(n56), .B1(n115), .B2(n25), .ZN(O[18]) );
  AOI21_X1 U107 ( .B1(n10), .B2(n56), .A(n5), .ZN(n115) );
  AOI22_X1 U108 ( .A1(n9), .A2(n25), .B1(A[18]), .B2(n2), .ZN(n114) );
  INV_X1 U109 ( .A(B[18]), .ZN(n56) );
  OAI22_X1 U110 ( .A1(n90), .A2(n69), .B1(n91), .B2(n37), .ZN(O[29]) );
  AOI21_X1 U111 ( .B1(n8), .B2(n69), .A(n6), .ZN(n91) );
  AOI22_X1 U112 ( .A1(n8), .A2(n37), .B1(A[29]), .B2(n3), .ZN(n90) );
  INV_X1 U113 ( .A(B[29]), .ZN(n69) );
  INV_X1 U114 ( .A(A[6]), .ZN(n44) );
  OAI22_X1 U115 ( .A1(n104), .A2(n60), .B1(n105), .B2(n30), .ZN(O[22]) );
  AOI21_X1 U116 ( .B1(n10), .B2(n60), .A(n6), .ZN(n105) );
  AOI22_X1 U117 ( .A1(n9), .A2(n30), .B1(A[22]), .B2(n3), .ZN(n104) );
  INV_X1 U118 ( .A(B[22]), .ZN(n60) );
  OAI22_X1 U119 ( .A1(n100), .A2(n62), .B1(n101), .B2(n32), .ZN(O[24]) );
  AOI21_X1 U120 ( .B1(n10), .B2(n62), .A(n6), .ZN(n101) );
  AOI22_X1 U121 ( .A1(n9), .A2(n32), .B1(A[24]), .B2(n3), .ZN(n100) );
  INV_X1 U122 ( .A(B[24]), .ZN(n62) );
  OAI22_X1 U123 ( .A1(n98), .A2(n63), .B1(n99), .B2(n33), .ZN(O[25]) );
  AOI21_X1 U124 ( .B1(n9), .B2(n63), .A(n6), .ZN(n99) );
  AOI22_X1 U125 ( .A1(n9), .A2(n33), .B1(A[25]), .B2(n3), .ZN(n98) );
  INV_X1 U126 ( .A(B[25]), .ZN(n63) );
  INV_X1 U127 ( .A(A[12]), .ZN(n19) );
  INV_X1 U128 ( .A(A[14]), .ZN(n21) );
  BUF_X1 U129 ( .A(n70), .Z(n7) );
  INV_X1 U130 ( .A(A[17]), .ZN(n24) );
  INV_X1 U131 ( .A(A[21]), .ZN(n29) );
  INV_X1 U132 ( .A(A[13]), .ZN(n20) );
  INV_X1 U133 ( .A(A[15]), .ZN(n22) );
  INV_X1 U134 ( .A(A[16]), .ZN(n23) );
  INV_X1 U135 ( .A(A[27]), .ZN(n35) );
  INV_X1 U136 ( .A(A[26]), .ZN(n34) );
  INV_X1 U137 ( .A(A[31]), .ZN(n40) );
  BUF_X1 U138 ( .A(n71), .Z(n4) );
  INV_X1 U139 ( .A(A[28]), .ZN(n36) );
  INV_X1 U140 ( .A(A[18]), .ZN(n25) );
  INV_X1 U141 ( .A(A[29]), .ZN(n37) );
  INV_X1 U142 ( .A(A[19]), .ZN(n26) );
  INV_X1 U143 ( .A(A[20]), .ZN(n28) );
  INV_X1 U144 ( .A(A[30]), .ZN(n39) );
  INV_X1 U145 ( .A(A[9]), .ZN(n47) );
  INV_X1 U146 ( .A(A[8]), .ZN(n46) );
  INV_X1 U147 ( .A(A[10]), .ZN(n17) );
  INV_X1 U148 ( .A(A[11]), .ZN(n18) );
  INV_X1 U149 ( .A(A[23]), .ZN(n31) );
  INV_X1 U150 ( .A(A[22]), .ZN(n30) );
  INV_X1 U151 ( .A(A[24]), .ZN(n32) );
  INV_X1 U152 ( .A(A[25]), .ZN(n33) );
  OAI22_X1 U153 ( .A1(n132), .A2(n11), .B1(n133), .B2(n16), .ZN(O[0]) );
  NOR2_X1 U154 ( .A1(n1), .A2(SEL[0]), .ZN(n70) );
  AND3_X1 U155 ( .A1(SEL[1]), .A2(SEL[0]), .A3(n134), .ZN(n71) );
  NOR3_X1 U156 ( .A1(SEL[2]), .A2(SEL[4]), .A3(SEL[3]), .ZN(n134) );
  OR4_X1 U157 ( .A1(n142), .A2(SEL[1]), .A3(SEL[3]), .A4(SEL[4]), .ZN(n1) );
  OAI22_X1 U158 ( .A1(n110), .A2(n12), .B1(n111), .B2(n27), .ZN(O[1]) );
  OAI22_X1 U159 ( .A1(n88), .A2(n13), .B1(n89), .B2(n38), .ZN(O[2]) );
  OAI22_X1 U160 ( .A1(n82), .A2(n14), .B1(n83), .B2(n41), .ZN(O[3]) );
  AOI22_X1 U161 ( .A1(n8), .A2(n38), .B1(A[2]), .B2(n3), .ZN(n88) );
  INV_X1 U162 ( .A(A[2]), .ZN(n38) );
  AOI22_X1 U163 ( .A1(n9), .A2(n43), .B1(A[5]), .B2(n4), .ZN(n78) );
  INV_X1 U164 ( .A(A[5]), .ZN(n43) );
  AOI22_X1 U165 ( .A1(n9), .A2(n42), .B1(A[4]), .B2(n4), .ZN(n80) );
  INV_X1 U166 ( .A(A[4]), .ZN(n42) );
  AOI22_X1 U167 ( .A1(n9), .A2(n27), .B1(A[1]), .B2(n2), .ZN(n110) );
  INV_X1 U168 ( .A(A[1]), .ZN(n27) );
  INV_X1 U169 ( .A(n1), .ZN(n8) );
  INV_X1 U170 ( .A(n1), .ZN(n9) );
  INV_X1 U171 ( .A(B[0]), .ZN(n11) );
  INV_X1 U172 ( .A(B[1]), .ZN(n12) );
  INV_X1 U173 ( .A(B[2]), .ZN(n13) );
  INV_X1 U174 ( .A(B[3]), .ZN(n14) );
  INV_X1 U175 ( .A(B[4]), .ZN(n15) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  INV_X1 U2 ( .A(SH[1]), .ZN(n6) );
  AOI221_X1 U3 ( .B1(n95), .B2(A[14]), .C1(n96), .C2(A[15]), .A(n17), .ZN(n150) );
  AOI221_X1 U4 ( .B1(n95), .B2(A[8]), .C1(n96), .C2(A[9]), .A(n107), .ZN(n79)
         );
  AOI221_X1 U5 ( .B1(n95), .B2(A[9]), .C1(n96), .C2(A[10]), .A(n97), .ZN(n74)
         );
  AOI221_X1 U6 ( .B1(n95), .B2(A[11]), .C1(n96), .C2(A[12]), .A(n131), .ZN(n61) );
  AOI221_X1 U7 ( .B1(n112), .B2(n113), .C1(n114), .C2(n115), .A(n46), .ZN(n63)
         );
  NOR2_X2 U8 ( .A1(n6), .A2(SH[0]), .ZN(n95) );
  AOI221_X1 U9 ( .B1(n118), .B2(n113), .C1(n119), .C2(n115), .A(n46), .ZN(n75)
         );
  NOR2_X2 U10 ( .A1(SH[2]), .A2(SH[3]), .ZN(n115) );
  INV_X1 U11 ( .A(n99), .ZN(n1) );
  NAND2_X1 U12 ( .A1(n60), .A2(n12), .ZN(n2) );
  NAND2_X1 U13 ( .A1(n65), .A2(n16), .ZN(n3) );
  NAND2_X1 U14 ( .A1(n67), .A2(n72), .ZN(n4) );
  AND3_X1 U15 ( .A1(n2), .A2(n3), .A3(n4), .ZN(n88) );
  INV_X1 U16 ( .A(n99), .ZN(n57) );
  INV_X2 U17 ( .A(n89), .ZN(n60) );
  AND2_X2 U18 ( .A1(SH[2]), .A2(n167), .ZN(n67) );
  AOI221_X1 U19 ( .B1(n95), .B2(A[10]), .C1(n96), .C2(A[11]), .A(n166), .ZN(
        n69) );
  INV_X2 U20 ( .A(n98), .ZN(n55) );
  NAND2_X2 U21 ( .A1(n5), .A2(n6), .ZN(n99) );
  INV_X2 U22 ( .A(n95), .ZN(n58) );
  NAND2_X2 U23 ( .A1(n115), .A2(n8), .ZN(n62) );
  INV_X1 U24 ( .A(n96), .ZN(n56) );
  INV_X1 U25 ( .A(SH[4]), .ZN(n8) );
  INV_X1 U26 ( .A(n62), .ZN(n59) );
  INV_X1 U27 ( .A(n138), .ZN(n24) );
  INV_X1 U28 ( .A(n139), .ZN(n33) );
  INV_X1 U29 ( .A(n127), .ZN(n39) );
  INV_X1 U30 ( .A(n135), .ZN(n36) );
  INV_X1 U31 ( .A(n170), .ZN(n32) );
  INV_X1 U32 ( .A(n126), .ZN(n40) );
  INV_X1 U33 ( .A(n122), .ZN(n43) );
  NOR2_X2 U34 ( .A1(n5), .A2(n6), .ZN(n96) );
  INV_X1 U35 ( .A(n101), .ZN(n47) );
  INV_X1 U36 ( .A(n78), .ZN(n26) );
  AND2_X2 U37 ( .A1(n167), .A2(n7), .ZN(n65) );
  INV_X1 U38 ( .A(n133), .ZN(n18) );
  INV_X1 U39 ( .A(n150), .ZN(n16) );
  INV_X1 U40 ( .A(n142), .ZN(n20) );
  INV_X1 U41 ( .A(n136), .ZN(n46) );
  INV_X1 U42 ( .A(n69), .ZN(n12) );
  INV_X1 U43 ( .A(n61), .ZN(n10) );
  INV_X1 U44 ( .A(n105), .ZN(n9) );
  INV_X1 U45 ( .A(n93), .ZN(n13) );
  INV_X1 U46 ( .A(n77), .ZN(n22) );
  INV_X1 U47 ( .A(A[3]), .ZN(n48) );
  INV_X1 U48 ( .A(A[17]), .ZN(n23) );
  INV_X1 U49 ( .A(A[12]), .ZN(n15) );
  INV_X1 U50 ( .A(n149), .ZN(n19) );
  INV_X1 U51 ( .A(n161), .ZN(n21) );
  INV_X1 U52 ( .A(A[23]), .ZN(n30) );
  INV_X1 U53 ( .A(A[21]), .ZN(n29) );
  INV_X1 U54 ( .A(A[6]), .ZN(n51) );
  INV_X1 U55 ( .A(A[7]), .ZN(n52) );
  INV_X1 U56 ( .A(\A[31] ), .ZN(n45) );
  INV_X1 U57 ( .A(A[18]), .ZN(n25) );
  INV_X1 U58 ( .A(A[19]), .ZN(n27) );
  INV_X1 U59 ( .A(A[29]), .ZN(n41) );
  INV_X1 U60 ( .A(A[27]), .ZN(n37) );
  INV_X1 U61 ( .A(A[26]), .ZN(n35) );
  INV_X1 U62 ( .A(A[28]), .ZN(n38) );
  INV_X1 U63 ( .A(A[20]), .ZN(n28) );
  INV_X1 U64 ( .A(A[30]), .ZN(n44) );
  INV_X1 U65 ( .A(A[9]), .ZN(n54) );
  INV_X1 U66 ( .A(A[8]), .ZN(n53) );
  INV_X1 U67 ( .A(A[10]), .ZN(n11) );
  INV_X1 U68 ( .A(A[11]), .ZN(n14) );
  INV_X1 U69 ( .A(A[24]), .ZN(n31) );
  INV_X1 U70 ( .A(A[25]), .ZN(n34) );
  INV_X1 U71 ( .A(n169), .ZN(n17) );
  INV_X1 U72 ( .A(A[2]), .ZN(n42) );
  NAND2_X1 U73 ( .A1(SH[0]), .A2(n6), .ZN(n98) );
  INV_X1 U74 ( .A(A[5]), .ZN(n50) );
  INV_X1 U75 ( .A(A[4]), .ZN(n49) );
  INV_X1 U76 ( .A(SH[0]), .ZN(n5) );
  INV_X1 U77 ( .A(SH[2]), .ZN(n7) );
  OAI221_X1 U78 ( .B1(n61), .B2(n62), .C1(n63), .C2(n8), .A(n64), .ZN(B[9]) );
  AOI222_X1 U79 ( .A1(n60), .A2(n18), .B1(n65), .B2(n66), .C1(n67), .C2(n68), 
        .ZN(n64) );
  OAI221_X1 U80 ( .B1(n69), .B2(n62), .C1(n70), .C2(n8), .A(n71), .ZN(B[8]) );
  AOI222_X1 U81 ( .A1(n60), .A2(n16), .B1(n65), .B2(n72), .C1(n67), .C2(n73), 
        .ZN(n71) );
  OAI221_X1 U82 ( .B1(n74), .B2(n62), .C1(n75), .C2(n8), .A(n76), .ZN(B[7]) );
  AOI222_X1 U83 ( .A1(n60), .A2(n13), .B1(n65), .B2(n77), .C1(n67), .C2(n78), 
        .ZN(n76) );
  OAI221_X1 U84 ( .B1(n79), .B2(n62), .C1(n80), .C2(n8), .A(n81), .ZN(B[6]) );
  AOI222_X1 U85 ( .A1(n60), .A2(n9), .B1(n65), .B2(n20), .C1(n67), .C2(n82), 
        .ZN(n81) );
  OAI221_X1 U86 ( .B1(n83), .B2(n62), .C1(n84), .C2(n8), .A(n85), .ZN(B[5]) );
  AOI222_X1 U87 ( .A1(n60), .A2(n10), .B1(n65), .B2(n18), .C1(n67), .C2(n66), 
        .ZN(n85) );
  OAI221_X1 U88 ( .B1(n86), .B2(n62), .C1(n87), .C2(n8), .A(n88), .ZN(B[4]) );
  OAI221_X1 U89 ( .B1(n74), .B2(n89), .C1(n90), .C2(n8), .A(n91), .ZN(B[3]) );
  AOI222_X1 U90 ( .A1(n67), .A2(n77), .B1(n59), .B2(n92), .C1(n65), .C2(n13), 
        .ZN(n91) );
  OAI221_X1 U91 ( .B1(n58), .B2(n50), .C1(n56), .C2(n51), .A(n94), .ZN(n92) );
  AOI22_X1 U92 ( .A1(A[4]), .A2(n55), .B1(A[3]), .B2(n1), .ZN(n94) );
  OAI22_X1 U93 ( .A1(n53), .A2(n98), .B1(n52), .B2(n99), .ZN(n97) );
  OAI21_X1 U94 ( .B1(SH[4]), .B2(n100), .A(n101), .ZN(B[30]) );
  OAI221_X1 U95 ( .B1(n79), .B2(n89), .C1(n102), .C2(n8), .A(n103), .ZN(B[2])
         );
  AOI222_X1 U96 ( .A1(n67), .A2(n20), .B1(n59), .B2(n104), .C1(n65), .C2(n9), 
        .ZN(n103) );
  OAI221_X1 U97 ( .B1(n58), .B2(n49), .C1(n56), .C2(n50), .A(n106), .ZN(n104)
         );
  AOI22_X1 U98 ( .A1(A[3]), .A2(n55), .B1(A[2]), .B2(n1), .ZN(n106) );
  OAI22_X1 U99 ( .A1(n52), .A2(n98), .B1(n51), .B2(n99), .ZN(n107) );
  OAI21_X1 U100 ( .B1(SH[4]), .B2(n108), .A(n101), .ZN(B[29]) );
  OAI21_X1 U101 ( .B1(SH[4]), .B2(n109), .A(n101), .ZN(B[28]) );
  OAI21_X1 U102 ( .B1(SH[4]), .B2(n110), .A(n101), .ZN(B[27]) );
  OAI21_X1 U103 ( .B1(SH[4]), .B2(n111), .A(n101), .ZN(B[26]) );
  OAI21_X1 U104 ( .B1(SH[4]), .B2(n63), .A(n101), .ZN(B[25]) );
  OAI21_X1 U105 ( .B1(SH[4]), .B2(n70), .A(n101), .ZN(B[24]) );
  AOI221_X1 U106 ( .B1(n116), .B2(n113), .C1(n117), .C2(n115), .A(n46), .ZN(
        n70) );
  OAI21_X1 U107 ( .B1(SH[4]), .B2(n75), .A(n101), .ZN(B[23]) );
  OAI21_X1 U108 ( .B1(SH[4]), .B2(n80), .A(n101), .ZN(B[22]) );
  AOI221_X1 U109 ( .B1(n120), .B2(n113), .C1(n121), .C2(n115), .A(n43), .ZN(
        n80) );
  AOI21_X1 U110 ( .B1(n123), .B2(n124), .A(n125), .ZN(n122) );
  OAI21_X1 U111 ( .B1(SH[4]), .B2(n84), .A(n101), .ZN(B[21]) );
  AOI221_X1 U112 ( .B1(n114), .B2(n113), .C1(n68), .C2(n115), .A(n40), .ZN(n84) );
  AOI21_X1 U113 ( .B1(n123), .B2(n112), .A(n125), .ZN(n126) );
  OAI21_X1 U114 ( .B1(SH[4]), .B2(n87), .A(n101), .ZN(B[20]) );
  AOI221_X1 U115 ( .B1(n117), .B2(n113), .C1(n73), .C2(n115), .A(n39), .ZN(n87) );
  AOI21_X1 U116 ( .B1(n123), .B2(n116), .A(n125), .ZN(n127) );
  OAI221_X1 U117 ( .B1(n83), .B2(n89), .C1(n128), .C2(n8), .A(n129), .ZN(B[1])
         );
  AOI222_X1 U118 ( .A1(n67), .A2(n18), .B1(n59), .B2(n130), .C1(n65), .C2(n10), 
        .ZN(n129) );
  OAI22_X1 U119 ( .A1(n11), .A2(n98), .B1(n54), .B2(n99), .ZN(n131) );
  OAI221_X1 U120 ( .B1(n58), .B2(n48), .C1(n56), .C2(n49), .A(n132), .ZN(n130)
         );
  AOI22_X1 U121 ( .A1(A[2]), .A2(n55), .B1(A[1]), .B2(n1), .ZN(n132) );
  AOI221_X1 U122 ( .B1(n95), .B2(A[7]), .C1(n96), .C2(A[8]), .A(n134), .ZN(n83) );
  OAI22_X1 U123 ( .A1(n51), .A2(n98), .B1(n50), .B2(n99), .ZN(n134) );
  OAI21_X1 U124 ( .B1(SH[4]), .B2(n90), .A(n101), .ZN(B[19]) );
  AOI221_X1 U125 ( .B1(n119), .B2(n113), .C1(n78), .C2(n115), .A(n36), .ZN(n90) );
  AOI21_X1 U126 ( .B1(n123), .B2(n118), .A(n125), .ZN(n135) );
  NOR2_X1 U127 ( .A1(n136), .A2(n7), .ZN(n125) );
  OAI21_X1 U128 ( .B1(SH[4]), .B2(n102), .A(n101), .ZN(B[18]) );
  AOI221_X1 U129 ( .B1(n124), .B2(n137), .C1(n120), .C2(n123), .A(n24), .ZN(
        n102) );
  AOI22_X1 U130 ( .A1(n113), .A2(n121), .B1(n115), .B2(n82), .ZN(n138) );
  OAI21_X1 U131 ( .B1(SH[4]), .B2(n128), .A(n101), .ZN(B[17]) );
  AOI221_X1 U132 ( .B1(n68), .B2(n113), .C1(n66), .C2(n115), .A(n33), .ZN(n128) );
  AOI22_X1 U133 ( .A1(n137), .A2(n112), .B1(n123), .B2(n114), .ZN(n139) );
  OAI21_X1 U134 ( .B1(SH[4]), .B2(n140), .A(n101), .ZN(B[16]) );
  OAI221_X1 U135 ( .B1(n26), .B2(n89), .C1(n22), .C2(n62), .A(n141), .ZN(B[15]) );
  AOI221_X1 U136 ( .B1(n67), .B2(n118), .C1(n65), .C2(n119), .A(n47), .ZN(n141) );
  NAND2_X1 U137 ( .A1(SH[4]), .A2(\A[31] ), .ZN(n101) );
  OAI221_X1 U138 ( .B1(n142), .B2(n62), .C1(n100), .C2(n8), .A(n143), .ZN(
        B[14]) );
  AOI222_X1 U139 ( .A1(n60), .A2(n82), .B1(n65), .B2(n121), .C1(n67), .C2(n120), .ZN(n143) );
  AOI21_X1 U140 ( .B1(n124), .B2(n115), .A(n144), .ZN(n100) );
  OAI221_X1 U141 ( .B1(n133), .B2(n62), .C1(n108), .C2(n8), .A(n145), .ZN(
        B[13]) );
  AOI222_X1 U142 ( .A1(n60), .A2(n66), .B1(n65), .B2(n68), .C1(n67), .C2(n114), 
        .ZN(n145) );
  OAI221_X1 U143 ( .B1(n58), .B2(n37), .C1(n56), .C2(n38), .A(n146), .ZN(n114)
         );
  AOI22_X1 U144 ( .A1(A[26]), .A2(n55), .B1(A[25]), .B2(n57), .ZN(n146) );
  OAI221_X1 U145 ( .B1(n58), .B2(n30), .C1(n56), .C2(n31), .A(n147), .ZN(n68)
         );
  AOI22_X1 U146 ( .A1(A[22]), .A2(n55), .B1(A[21]), .B2(n57), .ZN(n147) );
  OAI221_X1 U147 ( .B1(n58), .B2(n27), .C1(n56), .C2(n28), .A(n148), .ZN(n66)
         );
  AOI22_X1 U148 ( .A1(A[18]), .A2(n55), .B1(A[17]), .B2(n57), .ZN(n148) );
  AOI21_X1 U149 ( .B1(n112), .B2(n115), .A(n144), .ZN(n108) );
  OAI222_X1 U150 ( .A1(n99), .A2(n41), .B1(n98), .B2(n44), .C1(n6), .C2(n45), 
        .ZN(n112) );
  AOI221_X1 U151 ( .B1(n95), .B2(A[15]), .C1(n96), .C2(A[16]), .A(n19), .ZN(
        n133) );
  AOI22_X1 U152 ( .A1(A[14]), .A2(n55), .B1(A[13]), .B2(n57), .ZN(n149) );
  OAI221_X1 U153 ( .B1(n150), .B2(n62), .C1(n109), .C2(n8), .A(n151), .ZN(
        B[12]) );
  AOI222_X1 U154 ( .A1(n60), .A2(n72), .B1(n65), .B2(n73), .C1(n67), .C2(n117), 
        .ZN(n151) );
  AOI21_X1 U155 ( .B1(n116), .B2(n115), .A(n144), .ZN(n109) );
  OAI221_X1 U156 ( .B1(n93), .B2(n62), .C1(n110), .C2(n8), .A(n152), .ZN(B[11]) );
  AOI222_X1 U157 ( .A1(n60), .A2(n77), .B1(n65), .B2(n78), .C1(n67), .C2(n119), 
        .ZN(n152) );
  OAI221_X1 U158 ( .B1(n58), .B2(n34), .C1(n56), .C2(n35), .A(n153), .ZN(n119)
         );
  AOI22_X1 U159 ( .A1(A[24]), .A2(n55), .B1(A[23]), .B2(n57), .ZN(n153) );
  OAI221_X1 U160 ( .B1(n28), .B2(n98), .C1(n27), .C2(n99), .A(n154), .ZN(n78)
         );
  AOI22_X1 U161 ( .A1(A[21]), .A2(n95), .B1(A[22]), .B2(n96), .ZN(n154) );
  OAI221_X1 U162 ( .B1(n58), .B2(n23), .C1(n56), .C2(n25), .A(n155), .ZN(n77)
         );
  AOI22_X1 U163 ( .A1(A[16]), .A2(n55), .B1(A[15]), .B2(n1), .ZN(n155) );
  AOI21_X1 U164 ( .B1(n118), .B2(n115), .A(n144), .ZN(n110) );
  OAI21_X1 U165 ( .B1(n7), .B2(n45), .A(n136), .ZN(n144) );
  OAI221_X1 U166 ( .B1(n58), .B2(n41), .C1(n56), .C2(n44), .A(n156), .ZN(n118)
         );
  AOI22_X1 U167 ( .A1(A[28]), .A2(n55), .B1(A[27]), .B2(n57), .ZN(n156) );
  AOI221_X1 U168 ( .B1(n95), .B2(A[13]), .C1(n96), .C2(A[14]), .A(n157), .ZN(
        n93) );
  OAI22_X1 U169 ( .A1(n15), .A2(n98), .B1(n14), .B2(n99), .ZN(n157) );
  OAI221_X1 U170 ( .B1(n105), .B2(n62), .C1(n111), .C2(n8), .A(n158), .ZN(
        B[10]) );
  AOI222_X1 U171 ( .A1(n60), .A2(n20), .B1(n65), .B2(n82), .C1(n67), .C2(n121), 
        .ZN(n158) );
  OAI221_X1 U172 ( .B1(n58), .B2(n31), .C1(n56), .C2(n34), .A(n159), .ZN(n121)
         );
  AOI22_X1 U173 ( .A1(A[23]), .A2(n55), .B1(A[22]), .B2(n57), .ZN(n159) );
  OAI221_X1 U174 ( .B1(n27), .B2(n98), .C1(n25), .C2(n99), .A(n160), .ZN(n82)
         );
  AOI22_X1 U175 ( .A1(A[20]), .A2(n95), .B1(A[21]), .B2(n96), .ZN(n160) );
  AOI221_X1 U176 ( .B1(n95), .B2(A[16]), .C1(n96), .C2(A[17]), .A(n21), .ZN(
        n142) );
  AOI22_X1 U177 ( .A1(A[15]), .A2(n55), .B1(A[14]), .B2(n57), .ZN(n161) );
  AOI221_X1 U178 ( .B1(n124), .B2(n113), .C1(n120), .C2(n115), .A(n46), .ZN(
        n111) );
  NAND2_X1 U179 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n136) );
  OAI221_X1 U180 ( .B1(n58), .B2(n38), .C1(n56), .C2(n41), .A(n162), .ZN(n120)
         );
  AOI22_X1 U181 ( .A1(A[27]), .A2(n55), .B1(A[26]), .B2(n57), .ZN(n162) );
  MUX2_X1 U182 ( .A(A[30]), .B(\A[31] ), .S(n99), .Z(n124) );
  AOI221_X1 U183 ( .B1(n95), .B2(A[12]), .C1(n96), .C2(A[13]), .A(n163), .ZN(
        n105) );
  OAI22_X1 U184 ( .A1(n14), .A2(n98), .B1(n11), .B2(n99), .ZN(n163) );
  OAI221_X1 U185 ( .B1(n86), .B2(n89), .C1(n140), .C2(n8), .A(n164), .ZN(B[0])
         );
  AOI222_X1 U186 ( .A1(n67), .A2(n16), .B1(n59), .B2(n165), .C1(n65), .C2(n12), 
        .ZN(n164) );
  OAI22_X1 U187 ( .A1(n54), .A2(n98), .B1(n53), .B2(n99), .ZN(n166) );
  OAI221_X1 U188 ( .B1(n58), .B2(n42), .C1(n56), .C2(n48), .A(n168), .ZN(n165)
         );
  AOI22_X1 U189 ( .A1(A[1]), .A2(n55), .B1(A[0]), .B2(n1), .ZN(n168) );
  AOI22_X1 U190 ( .A1(A[13]), .A2(n55), .B1(A[12]), .B2(n57), .ZN(n169) );
  AND2_X1 U191 ( .A1(SH[3]), .A2(n8), .ZN(n167) );
  AOI221_X1 U192 ( .B1(n73), .B2(n113), .C1(n72), .C2(n115), .A(n32), .ZN(n140) );
  AOI22_X1 U193 ( .A1(n137), .A2(n116), .B1(n123), .B2(n117), .ZN(n170) );
  OAI221_X1 U194 ( .B1(n58), .B2(n35), .C1(n56), .C2(n37), .A(n171), .ZN(n117)
         );
  AOI22_X1 U195 ( .A1(A[25]), .A2(n55), .B1(A[24]), .B2(n57), .ZN(n171) );
  AND2_X1 U196 ( .A1(SH[3]), .A2(n7), .ZN(n123) );
  OAI221_X1 U197 ( .B1(n58), .B2(n44), .C1(n56), .C2(n45), .A(n172), .ZN(n116)
         );
  AOI22_X1 U198 ( .A1(A[29]), .A2(n55), .B1(A[28]), .B2(n57), .ZN(n172) );
  AND2_X1 U199 ( .A1(SH[2]), .A2(SH[3]), .ZN(n137) );
  OAI221_X1 U200 ( .B1(n58), .B2(n25), .C1(n27), .C2(n56), .A(n173), .ZN(n72)
         );
  AOI22_X1 U201 ( .A1(A[17]), .A2(n55), .B1(A[16]), .B2(n57), .ZN(n173) );
  OAI221_X1 U202 ( .B1(n98), .B2(n29), .C1(n28), .C2(n99), .A(n174), .ZN(n73)
         );
  AOI22_X1 U203 ( .A1(A[22]), .A2(n95), .B1(A[23]), .B2(n96), .ZN(n174) );
  NAND2_X1 U204 ( .A1(n113), .A2(n8), .ZN(n89) );
  NOR2_X1 U205 ( .A1(n7), .A2(SH[3]), .ZN(n113) );
  AOI221_X1 U206 ( .B1(n95), .B2(A[6]), .C1(n96), .C2(A[7]), .A(n175), .ZN(n86) );
  OAI22_X1 U207 ( .A1(n50), .A2(n98), .B1(n49), .B2(n99), .ZN(n175) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;

  CLKBUF_X1 U3 ( .A(SH[4]), .Z(n5) );
  AOI221_X1 U4 ( .B1(n54), .B2(A[7]), .C1(n52), .C2(A[6]), .A(n165), .ZN(n86)
         );
  AOI221_X1 U5 ( .B1(n54), .B2(A[11]), .C1(n52), .C2(A[10]), .A(n156), .ZN(n67) );
  AOI221_X1 U6 ( .B1(n54), .B2(A[13]), .C1(n52), .C2(A[12]), .A(n153), .ZN(
        n105) );
  INV_X1 U7 ( .A(n140), .ZN(n57) );
  AOI221_X1 U8 ( .B1(n54), .B2(A[10]), .C1(n52), .C2(A[9]), .A(n99), .ZN(n73)
         );
  NAND2_X2 U9 ( .A1(SH[1]), .A2(SH[0]), .ZN(n94) );
  INV_X1 U10 ( .A(n97), .ZN(n53) );
  NOR2_X2 U11 ( .A1(SH[0]), .A2(SH[1]), .ZN(n98) );
  AOI221_X1 U12 ( .B1(n54), .B2(A[12]), .C1(n52), .C2(A[11]), .A(n122), .ZN(
        n58) );
  NOR2_X2 U13 ( .A1(n2), .A2(SH[1]), .ZN(n97) );
  INV_X1 U14 ( .A(n59), .ZN(n56) );
  INV_X1 U15 ( .A(SH[4]), .ZN(n6) );
  INV_X1 U16 ( .A(n89), .ZN(n55) );
  INV_X1 U17 ( .A(n160), .ZN(n32) );
  INV_X1 U18 ( .A(n126), .ZN(n35) );
  INV_X1 U19 ( .A(n139), .ZN(n27) );
  INV_X1 U20 ( .A(n94), .ZN(n54) );
  INV_X1 U21 ( .A(n128), .ZN(n33) );
  INV_X1 U22 ( .A(n95), .ZN(n52) );
  INV_X1 U23 ( .A(n81), .ZN(n16) );
  INV_X1 U24 ( .A(n138), .ZN(B[12]) );
  AND2_X2 U25 ( .A1(n157), .A2(n3), .ZN(n63) );
  INV_X1 U26 ( .A(n58), .ZN(n8) );
  INV_X1 U27 ( .A(n105), .ZN(n7) );
  INV_X1 U28 ( .A(n67), .ZN(n10) );
  INV_X1 U29 ( .A(n93), .ZN(n11) );
  INV_X1 U30 ( .A(n76), .ZN(n18) );
  INV_X1 U31 ( .A(n62), .ZN(n15) );
  INV_X1 U32 ( .A(n64), .ZN(n21) );
  INV_X1 U33 ( .A(n82), .ZN(n23) );
  INV_X1 U34 ( .A(n77), .ZN(n25) );
  INV_X1 U35 ( .A(A[3]), .ZN(n44) );
  INV_X1 U36 ( .A(n125), .ZN(n37) );
  INV_X1 U37 ( .A(A[14]), .ZN(n17) );
  INV_X1 U38 ( .A(A[23]), .ZN(n30) );
  INV_X1 U39 ( .A(A[12]), .ZN(n13) );
  INV_X1 U40 ( .A(A[6]), .ZN(n47) );
  INV_X1 U41 ( .A(A[7]), .ZN(n48) );
  INV_X1 U42 ( .A(A[31]), .ZN(n43) );
  INV_X1 U43 ( .A(A[17]), .ZN(n22) );
  INV_X1 U44 ( .A(A[21]), .ZN(n29) );
  INV_X1 U45 ( .A(A[20]), .ZN(n28) );
  INV_X1 U46 ( .A(A[15]), .ZN(n19) );
  INV_X1 U47 ( .A(A[16]), .ZN(n20) );
  INV_X1 U48 ( .A(A[29]), .ZN(n40) );
  INV_X1 U49 ( .A(A[27]), .ZN(n38) );
  INV_X1 U50 ( .A(A[26]), .ZN(n36) );
  INV_X1 U51 ( .A(A[30]), .ZN(n42) );
  INV_X1 U52 ( .A(A[28]), .ZN(n39) );
  INV_X1 U53 ( .A(A[18]), .ZN(n24) );
  INV_X1 U54 ( .A(A[19]), .ZN(n26) );
  INV_X1 U55 ( .A(A[9]), .ZN(n50) );
  INV_X1 U56 ( .A(A[8]), .ZN(n49) );
  INV_X1 U57 ( .A(A[10]), .ZN(n9) );
  INV_X1 U58 ( .A(A[11]), .ZN(n12) );
  INV_X1 U59 ( .A(A[24]), .ZN(n31) );
  INV_X1 U60 ( .A(A[25]), .ZN(n34) );
  AND2_X1 U61 ( .A1(SH[2]), .A2(n157), .ZN(n65) );
  INV_X1 U62 ( .A(A[2]), .ZN(n41) );
  NAND2_X1 U63 ( .A1(SH[1]), .A2(n2), .ZN(n95) );
  INV_X1 U64 ( .A(A[5]), .ZN(n46) );
  INV_X1 U65 ( .A(A[4]), .ZN(n45) );
  NAND2_X1 U66 ( .A1(SH[1]), .A2(n2), .ZN(n1) );
  INV_X1 U67 ( .A(SH[0]), .ZN(n2) );
  INV_X1 U68 ( .A(SH[2]), .ZN(n3) );
  INV_X1 U69 ( .A(SH[3]), .ZN(n4) );
  INV_X2 U70 ( .A(n98), .ZN(n51) );
  OAI221_X1 U71 ( .B1(n58), .B2(n59), .C1(n60), .C2(n6), .A(n61), .ZN(B[9]) );
  AOI222_X1 U72 ( .A1(n55), .A2(n62), .B1(n63), .B2(n64), .C1(n65), .C2(n66), 
        .ZN(n61) );
  OAI221_X1 U73 ( .B1(n67), .B2(n59), .C1(n68), .C2(n6), .A(n69), .ZN(B[8]) );
  AOI222_X1 U74 ( .A1(n55), .A2(n70), .B1(n63), .B2(n71), .C1(n65), .C2(n72), 
        .ZN(n69) );
  OAI221_X1 U75 ( .B1(n73), .B2(n59), .C1(n74), .C2(n6), .A(n75), .ZN(B[7]) );
  AOI222_X1 U76 ( .A1(n55), .A2(n11), .B1(n63), .B2(n76), .C1(n65), .C2(n77), 
        .ZN(n75) );
  OAI221_X1 U77 ( .B1(n78), .B2(n59), .C1(n79), .C2(n6), .A(n80), .ZN(B[6]) );
  AOI222_X1 U78 ( .A1(n55), .A2(n7), .B1(n63), .B2(n81), .C1(n65), .C2(n82), 
        .ZN(n80) );
  OAI221_X1 U79 ( .B1(n83), .B2(n59), .C1(n84), .C2(n6), .A(n85), .ZN(B[5]) );
  AOI222_X1 U80 ( .A1(n55), .A2(n8), .B1(n63), .B2(n62), .C1(n65), .C2(n64), 
        .ZN(n85) );
  OAI221_X1 U81 ( .B1(n86), .B2(n59), .C1(n87), .C2(n6), .A(n88), .ZN(B[4]) );
  AOI222_X1 U82 ( .A1(n55), .A2(n10), .B1(n63), .B2(n70), .C1(n65), .C2(n71), 
        .ZN(n88) );
  OAI221_X1 U83 ( .B1(n73), .B2(n89), .C1(n90), .C2(n6), .A(n91), .ZN(B[3]) );
  AOI222_X1 U84 ( .A1(n65), .A2(n76), .B1(n56), .B2(n92), .C1(n63), .C2(n11), 
        .ZN(n91) );
  OAI221_X1 U85 ( .B1(n94), .B2(n47), .C1(n95), .C2(n46), .A(n96), .ZN(n92) );
  AOI22_X1 U86 ( .A1(A[4]), .A2(n97), .B1(A[3]), .B2(n98), .ZN(n96) );
  OAI22_X1 U87 ( .A1(n49), .A2(n53), .B1(n48), .B2(n51), .ZN(n99) );
  AND2_X1 U88 ( .A1(n56), .A2(n100), .ZN(B[31]) );
  AND2_X1 U89 ( .A1(n101), .A2(n56), .ZN(B[30]) );
  OAI221_X1 U90 ( .B1(n78), .B2(n89), .C1(n102), .C2(n6), .A(n103), .ZN(B[2])
         );
  AOI222_X1 U91 ( .A1(n65), .A2(n81), .B1(n56), .B2(n104), .C1(n63), .C2(n7), 
        .ZN(n103) );
  OAI221_X1 U92 ( .B1(n94), .B2(n46), .C1(n1), .C2(n45), .A(n106), .ZN(n104)
         );
  AOI22_X1 U93 ( .A1(A[3]), .A2(n97), .B1(A[2]), .B2(n98), .ZN(n106) );
  AOI221_X1 U94 ( .B1(n54), .B2(A[9]), .C1(n52), .C2(A[8]), .A(n107), .ZN(n78)
         );
  OAI22_X1 U95 ( .A1(n48), .A2(n53), .B1(n47), .B2(n51), .ZN(n107) );
  AND2_X1 U96 ( .A1(n108), .A2(n56), .ZN(B[29]) );
  AND2_X1 U97 ( .A1(n109), .A2(n56), .ZN(B[28]) );
  NOR3_X1 U98 ( .A1(n37), .A2(n5), .A3(SH[3]), .ZN(B[27]) );
  NOR2_X1 U99 ( .A1(n5), .A2(n110), .ZN(B[26]) );
  NOR2_X1 U100 ( .A1(n5), .A2(n60), .ZN(B[25]) );
  AOI22_X1 U101 ( .A1(n111), .A2(n57), .B1(n108), .B2(n112), .ZN(n60) );
  NOR2_X1 U102 ( .A1(n5), .A2(n68), .ZN(B[24]) );
  AOI22_X1 U103 ( .A1(n113), .A2(n57), .B1(n109), .B2(n112), .ZN(n68) );
  NOR2_X1 U104 ( .A1(n5), .A2(n74), .ZN(B[23]) );
  AOI222_X1 U105 ( .A1(n114), .A2(n112), .B1(n100), .B2(n115), .C1(n116), .C2(
        n57), .ZN(n74) );
  NOR2_X1 U106 ( .A1(n5), .A2(n79), .ZN(B[22]) );
  AOI222_X1 U107 ( .A1(n117), .A2(n112), .B1(n101), .B2(n115), .C1(n118), .C2(
        n57), .ZN(n79) );
  NOR2_X1 U108 ( .A1(n5), .A2(n84), .ZN(B[21]) );
  AOI222_X1 U109 ( .A1(n111), .A2(n112), .B1(n108), .B2(n115), .C1(n66), .C2(
        n57), .ZN(n84) );
  NOR2_X1 U110 ( .A1(n5), .A2(n87), .ZN(B[20]) );
  AOI222_X1 U111 ( .A1(n113), .A2(n112), .B1(n109), .B2(n115), .C1(n72), .C2(
        n57), .ZN(n87) );
  OAI221_X1 U112 ( .B1(n83), .B2(n89), .C1(n119), .C2(n6), .A(n120), .ZN(B[1])
         );
  AOI222_X1 U113 ( .A1(n65), .A2(n62), .B1(n56), .B2(n121), .C1(n63), .C2(n8), 
        .ZN(n120) );
  OAI22_X1 U114 ( .A1(n9), .A2(n53), .B1(n50), .B2(n51), .ZN(n122) );
  OAI221_X1 U115 ( .B1(n94), .B2(n45), .C1(n1), .C2(n44), .A(n123), .ZN(n121)
         );
  AOI22_X1 U116 ( .A1(A[2]), .A2(n97), .B1(A[1]), .B2(n98), .ZN(n123) );
  AOI221_X1 U117 ( .B1(n54), .B2(A[8]), .C1(n52), .C2(A[7]), .A(n124), .ZN(n83) );
  OAI22_X1 U118 ( .A1(n47), .A2(n53), .B1(n46), .B2(n51), .ZN(n124) );
  NOR2_X1 U119 ( .A1(n5), .A2(n90), .ZN(B[19]) );
  AOI222_X1 U120 ( .A1(n77), .A2(n57), .B1(n116), .B2(n112), .C1(n125), .C2(
        SH[3]), .ZN(n90) );
  NOR2_X1 U121 ( .A1(n5), .A2(n102), .ZN(B[18]) );
  AOI221_X1 U122 ( .B1(n118), .B2(n112), .C1(n82), .C2(n57), .A(n35), .ZN(n102) );
  AOI22_X1 U123 ( .A1(n127), .A2(n101), .B1(n115), .B2(n117), .ZN(n126) );
  NOR2_X1 U124 ( .A1(n5), .A2(n119), .ZN(B[17]) );
  AOI221_X1 U125 ( .B1(n66), .B2(n112), .C1(n64), .C2(n57), .A(n33), .ZN(n119)
         );
  AOI22_X1 U126 ( .A1(n127), .A2(n108), .B1(n115), .B2(n111), .ZN(n128) );
  NOR2_X1 U127 ( .A1(n5), .A2(n129), .ZN(B[16]) );
  OAI221_X1 U128 ( .B1(n25), .B2(n89), .C1(n18), .C2(n59), .A(n130), .ZN(B[15]) );
  AOI222_X1 U129 ( .A1(n65), .A2(n114), .B1(n131), .B2(n100), .C1(n63), .C2(
        n116), .ZN(n130) );
  OAI221_X1 U130 ( .B1(n23), .B2(n89), .C1(n16), .C2(n59), .A(n132), .ZN(B[14]) );
  AOI222_X1 U131 ( .A1(n65), .A2(n117), .B1(n131), .B2(n101), .C1(n63), .C2(
        n118), .ZN(n132) );
  OAI221_X1 U132 ( .B1(n21), .B2(n89), .C1(n15), .C2(n59), .A(n133), .ZN(B[13]) );
  AOI222_X1 U133 ( .A1(n65), .A2(n111), .B1(n131), .B2(n108), .C1(n63), .C2(
        n66), .ZN(n133) );
  OAI221_X1 U134 ( .B1(n94), .B2(n31), .C1(n95), .C2(n30), .A(n134), .ZN(n66)
         );
  AOI22_X1 U135 ( .A1(A[22]), .A2(n97), .B1(A[21]), .B2(n98), .ZN(n134) );
  OAI222_X1 U136 ( .A1(n53), .A2(n42), .B1(n95), .B2(n43), .C1(n51), .C2(n40), 
        .ZN(n108) );
  OAI221_X1 U137 ( .B1(n94), .B2(n39), .C1(n1), .C2(n38), .A(n135), .ZN(n111)
         );
  AOI22_X1 U138 ( .A1(A[26]), .A2(n97), .B1(A[25]), .B2(n98), .ZN(n135) );
  OAI221_X1 U139 ( .B1(n94), .B2(n20), .C1(n95), .C2(n19), .A(n136), .ZN(n62)
         );
  AOI22_X1 U140 ( .A1(A[14]), .A2(n97), .B1(A[13]), .B2(n98), .ZN(n136) );
  OAI221_X1 U141 ( .B1(n94), .B2(n28), .C1(n1), .C2(n26), .A(n137), .ZN(n64)
         );
  AOI22_X1 U142 ( .A1(A[18]), .A2(n97), .B1(A[17]), .B2(n98), .ZN(n137) );
  AOI221_X1 U143 ( .B1(n71), .B2(n55), .C1(n70), .C2(n56), .A(n27), .ZN(n138)
         );
  AOI222_X1 U144 ( .A1(n65), .A2(n113), .B1(n131), .B2(n109), .C1(n63), .C2(
        n72), .ZN(n139) );
  NOR2_X1 U145 ( .A1(n6), .A2(n140), .ZN(n131) );
  OAI221_X1 U146 ( .B1(n18), .B2(n89), .C1(n93), .C2(n59), .A(n141), .ZN(B[11]) );
  AOI221_X1 U147 ( .B1(n65), .B2(n116), .C1(n63), .C2(n77), .A(n142), .ZN(n141) );
  NOR3_X1 U148 ( .A1(n6), .A2(SH[3]), .A3(n37), .ZN(n142) );
  MUX2_X1 U149 ( .A(n114), .B(n100), .S(SH[2]), .Z(n125) );
  NOR2_X1 U150 ( .A1(n43), .A2(n51), .ZN(n100) );
  OAI221_X1 U151 ( .B1(n94), .B2(n42), .C1(n95), .C2(n40), .A(n143), .ZN(n114)
         );
  AOI22_X1 U152 ( .A1(A[28]), .A2(n97), .B1(A[27]), .B2(n98), .ZN(n143) );
  OAI221_X1 U153 ( .B1(n28), .B2(n53), .C1(n26), .C2(n51), .A(n144), .ZN(n77)
         );
  AOI22_X1 U154 ( .A1(A[22]), .A2(n54), .B1(A[21]), .B2(n52), .ZN(n144) );
  OAI221_X1 U155 ( .B1(n94), .B2(n36), .C1(n1), .C2(n34), .A(n145), .ZN(n116)
         );
  AOI22_X1 U156 ( .A1(A[24]), .A2(n97), .B1(A[23]), .B2(n98), .ZN(n145) );
  AOI221_X1 U157 ( .B1(n54), .B2(A[14]), .C1(n52), .C2(A[13]), .A(n146), .ZN(
        n93) );
  OAI22_X1 U158 ( .A1(n13), .A2(n53), .B1(n12), .B2(n51), .ZN(n146) );
  OAI221_X1 U159 ( .B1(n94), .B2(n24), .C1(n95), .C2(n22), .A(n147), .ZN(n76)
         );
  AOI22_X1 U160 ( .A1(A[16]), .A2(n97), .B1(A[15]), .B2(n98), .ZN(n147) );
  OAI221_X1 U161 ( .B1(n105), .B2(n59), .C1(n110), .C2(n6), .A(n148), .ZN(
        B[10]) );
  AOI222_X1 U162 ( .A1(n55), .A2(n81), .B1(n63), .B2(n82), .C1(n65), .C2(n118), 
        .ZN(n148) );
  OAI221_X1 U163 ( .B1(n94), .B2(n34), .C1(n1), .C2(n31), .A(n149), .ZN(n118)
         );
  AOI22_X1 U164 ( .A1(A[23]), .A2(n97), .B1(A[22]), .B2(n98), .ZN(n149) );
  OAI221_X1 U165 ( .B1(n94), .B2(n29), .C1(n28), .C2(n1), .A(n150), .ZN(n82)
         );
  AOI22_X1 U166 ( .A1(n97), .A2(A[19]), .B1(n98), .B2(A[18]), .ZN(n150) );
  OAI221_X1 U167 ( .B1(n94), .B2(n22), .C1(n95), .C2(n20), .A(n151), .ZN(n81)
         );
  AOI22_X1 U168 ( .A1(A[15]), .A2(n97), .B1(A[14]), .B2(n98), .ZN(n151) );
  AOI22_X1 U169 ( .A1(n117), .A2(n57), .B1(n101), .B2(n112), .ZN(n110) );
  OAI22_X1 U170 ( .A1(n51), .A2(n42), .B1(n53), .B2(n43), .ZN(n101) );
  OAI221_X1 U171 ( .B1(n94), .B2(n40), .C1(n1), .C2(n39), .A(n152), .ZN(n117)
         );
  AOI22_X1 U172 ( .A1(A[27]), .A2(n97), .B1(A[26]), .B2(n98), .ZN(n152) );
  OAI22_X1 U173 ( .A1(n12), .A2(n53), .B1(n9), .B2(n51), .ZN(n153) );
  OAI221_X1 U174 ( .B1(n86), .B2(n89), .C1(n129), .C2(n6), .A(n154), .ZN(B[0])
         );
  AOI222_X1 U175 ( .A1(n65), .A2(n70), .B1(n56), .B2(n155), .C1(n63), .C2(n10), 
        .ZN(n154) );
  OAI22_X1 U176 ( .A1(n50), .A2(n53), .B1(n49), .B2(n51), .ZN(n156) );
  OAI221_X1 U177 ( .B1(n94), .B2(n44), .C1(n95), .C2(n41), .A(n158), .ZN(n155)
         );
  AOI22_X1 U178 ( .A1(A[1]), .A2(n97), .B1(A[0]), .B2(n98), .ZN(n158) );
  NAND2_X1 U179 ( .A1(n57), .A2(n6), .ZN(n59) );
  OAI221_X1 U180 ( .B1(n94), .B2(n19), .C1(n1), .C2(n17), .A(n159), .ZN(n70)
         );
  AOI22_X1 U181 ( .A1(A[13]), .A2(n97), .B1(A[12]), .B2(n98), .ZN(n159) );
  NOR2_X1 U182 ( .A1(n4), .A2(SH[4]), .ZN(n157) );
  AOI221_X1 U183 ( .B1(n72), .B2(n112), .C1(n71), .C2(n57), .A(n32), .ZN(n129)
         );
  AOI22_X1 U184 ( .A1(n127), .A2(n109), .B1(n115), .B2(n113), .ZN(n160) );
  OAI221_X1 U185 ( .B1(n94), .B2(n38), .C1(n95), .C2(n36), .A(n161), .ZN(n113)
         );
  AOI22_X1 U186 ( .A1(A[25]), .A2(n97), .B1(A[24]), .B2(n98), .ZN(n161) );
  NOR2_X1 U187 ( .A1(n4), .A2(SH[2]), .ZN(n115) );
  OAI221_X1 U188 ( .B1(n94), .B2(n43), .C1(n1), .C2(n42), .A(n162), .ZN(n109)
         );
  AOI22_X1 U189 ( .A1(A[29]), .A2(n97), .B1(A[28]), .B2(n98), .ZN(n162) );
  NOR2_X1 U190 ( .A1(n3), .A2(n4), .ZN(n127) );
  NAND2_X1 U191 ( .A1(n3), .A2(n4), .ZN(n140) );
  OAI221_X1 U192 ( .B1(n94), .B2(n26), .C1(n1), .C2(n24), .A(n163), .ZN(n71)
         );
  AOI22_X1 U193 ( .A1(A[17]), .A2(n97), .B1(A[16]), .B2(n98), .ZN(n163) );
  OAI221_X1 U194 ( .B1(n53), .B2(n29), .C1(n28), .C2(n51), .A(n164), .ZN(n72)
         );
  AOI22_X1 U195 ( .A1(A[23]), .A2(n54), .B1(A[22]), .B2(n52), .ZN(n164) );
  NAND2_X1 U196 ( .A1(n112), .A2(n6), .ZN(n89) );
  NOR2_X1 U197 ( .A1(n3), .A2(SH[3]), .ZN(n112) );
  OAI22_X1 U198 ( .A1(n46), .A2(n53), .B1(n45), .B2(n51), .ZN(n165) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][15] , \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] ,
         \ML_int[5][11] , \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] ,
         \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] ,
         \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(SH[4]), .Z(
        \ML_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(SH[4]), .Z(
        \ML_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(SH[4]), .Z(
        \ML_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(SH[4]), .Z(
        \ML_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(SH[4]), .Z(
        \ML_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(SH[4]), .Z(
        \ML_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(SH[4]), .Z(
        \ML_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(SH[4]), .Z(
        \ML_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(n23), .S(SH[4]), .Z(
        \ML_int[5][23] ) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(n19), .S(SH[4]), .Z(
        \ML_int[5][22] ) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(n21), .S(SH[4]), .Z(
        \ML_int[5][21] ) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(n17), .S(SH[4]), .Z(
        \ML_int[5][20] ) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(n22), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(n18), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(n20), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(n16), .S(SH[4]), .Z(
        \ML_int[5][16] ) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n13), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n13), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n13), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n13), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n13), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n13), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n13), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n13), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n13), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n13), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n13), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n13), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n12), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n12), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n12), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n12), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n12), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n12), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n12), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n12), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n12), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n12), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n12), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n12), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n10), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n10), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n10), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n10), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n10), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n10), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n10), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n10), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n10), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n10), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n10), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n10), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n10), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n10), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n10), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n9), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n9), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n9), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n9), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n9), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n9), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n9), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n9), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n9), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n9), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n9), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n9), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n7), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n7), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n7), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n7), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n7), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n7), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n6), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n6), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n6), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n6), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n6), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n6), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n6), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n6), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n6), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n6), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n6), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n6), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n5), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n5), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n5), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n5), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n5), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n5), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n5), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n5), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n5), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n5), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n5), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n5), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n3), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n3), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n2), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n2), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n2), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n3), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n1), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n2), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n3), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n3), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n1), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n2), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n1), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n2), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n1), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n3), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n1), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n2), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n1), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n3), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n1), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n2), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n1), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n2), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n1), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n3), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n1), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n2), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n2), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n2), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n2), .Z(\ML_int[1][1] ) );
  MUX2_X1 U3 ( .A(\ML_int[2][15] ), .B(\ML_int[2][19] ), .S(n11), .Z(
        \ML_int[3][19] ) );
  INV_X2 U4 ( .A(n11), .ZN(n10) );
  INV_X1 U5 ( .A(n11), .ZN(n9) );
  INV_X1 U6 ( .A(n30), .ZN(n20) );
  INV_X1 U7 ( .A(n31), .ZN(n16) );
  INV_X1 U8 ( .A(n29), .ZN(n18) );
  INV_X1 U9 ( .A(n28), .ZN(n22) );
  INV_X1 U10 ( .A(n26), .ZN(n21) );
  INV_X1 U11 ( .A(n27), .ZN(n17) );
  INV_X1 U12 ( .A(n25), .ZN(n19) );
  INV_X1 U13 ( .A(n24), .ZN(n23) );
  INV_X1 U14 ( .A(SH[3]), .ZN(n14) );
  INV_X1 U15 ( .A(SH[1]), .ZN(n8) );
  INV_X1 U16 ( .A(SH[0]), .ZN(n4) );
  INV_X2 U17 ( .A(n4), .ZN(n1) );
  INV_X2 U18 ( .A(n4), .ZN(n2) );
  INV_X2 U19 ( .A(n8), .ZN(n5) );
  INV_X2 U20 ( .A(n8), .ZN(n6) );
  INV_X1 U21 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(n8), .ZN(n7) );
  INV_X1 U23 ( .A(SH[2]), .ZN(n11) );
  INV_X1 U24 ( .A(n14), .ZN(n12) );
  INV_X1 U25 ( .A(n14), .ZN(n13) );
  INV_X1 U26 ( .A(SH[4]), .ZN(n15) );
  AND2_X1 U27 ( .A1(\ML_int[4][9] ), .A2(n15), .ZN(\ML_int[5][9] ) );
  AND2_X1 U28 ( .A1(\ML_int[4][8] ), .A2(n15), .ZN(\ML_int[5][8] ) );
  NOR2_X1 U29 ( .A1(SH[4]), .A2(n24), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U30 ( .A1(SH[4]), .A2(n25), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U31 ( .A1(SH[4]), .A2(n26), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U32 ( .A1(SH[4]), .A2(n27), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U33 ( .A1(SH[4]), .A2(n28), .ZN(\ML_int[5][3] ) );
  NOR2_X1 U34 ( .A1(SH[4]), .A2(n29), .ZN(\ML_int[5][2] ) );
  NOR2_X1 U35 ( .A1(SH[4]), .A2(n30), .ZN(\ML_int[5][1] ) );
  AND2_X1 U36 ( .A1(\ML_int[4][15] ), .A2(n15), .ZN(\ML_int[5][15] ) );
  AND2_X1 U37 ( .A1(\ML_int[4][14] ), .A2(n15), .ZN(\ML_int[5][14] ) );
  AND2_X1 U38 ( .A1(\ML_int[4][13] ), .A2(n15), .ZN(\ML_int[5][13] ) );
  AND2_X1 U39 ( .A1(\ML_int[4][12] ), .A2(n15), .ZN(\ML_int[5][12] ) );
  AND2_X1 U40 ( .A1(\ML_int[4][11] ), .A2(n15), .ZN(\ML_int[5][11] ) );
  AND2_X1 U41 ( .A1(\ML_int[4][10] ), .A2(n15), .ZN(\ML_int[5][10] ) );
  NOR2_X1 U42 ( .A1(SH[4]), .A2(n31), .ZN(\ML_int[5][0] ) );
  NAND2_X1 U43 ( .A1(\ML_int[3][7] ), .A2(n14), .ZN(n24) );
  NAND2_X1 U44 ( .A1(\ML_int[3][6] ), .A2(n14), .ZN(n25) );
  NAND2_X1 U45 ( .A1(\ML_int[3][5] ), .A2(n14), .ZN(n26) );
  NAND2_X1 U46 ( .A1(\ML_int[3][4] ), .A2(n14), .ZN(n27) );
  NAND2_X1 U47 ( .A1(\ML_int[3][3] ), .A2(n14), .ZN(n28) );
  NAND2_X1 U48 ( .A1(\ML_int[3][2] ), .A2(n14), .ZN(n29) );
  NAND2_X1 U49 ( .A1(\ML_int[3][1] ), .A2(n14), .ZN(n30) );
  NAND2_X1 U50 ( .A1(\ML_int[3][0] ), .A2(n14), .ZN(n31) );
  AND2_X1 U51 ( .A1(\ML_int[2][3] ), .A2(n11), .ZN(\ML_int[3][3] ) );
  AND2_X1 U52 ( .A1(\ML_int[2][2] ), .A2(n11), .ZN(\ML_int[3][2] ) );
  AND2_X1 U53 ( .A1(\ML_int[2][1] ), .A2(n11), .ZN(\ML_int[3][1] ) );
  AND2_X1 U54 ( .A1(\ML_int[2][0] ), .A2(n11), .ZN(\ML_int[3][0] ) );
  AND2_X1 U55 ( .A1(\ML_int[1][1] ), .A2(n8), .ZN(\ML_int[2][1] ) );
  AND2_X1 U56 ( .A1(\ML_int[1][0] ), .A2(n8), .ZN(\ML_int[2][0] ) );
  AND2_X1 U57 ( .A1(A[0]), .A2(n4), .ZN(\ML_int[1][0] ) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, .sel({\sel[4] , \sel[3] , \sel[2] , 
        \sel[1] , \sel[0] }), OUTPUT );
  input [31:0] A;
  input [31:0] B;
  output [31:0] OUTPUT;
  input \sel[4] , \sel[3] , \sel[2] , \sel[1] , \sel[0] ;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n1, n2, n3, n4, n5, n6, n10, n11, n12, n82, n83, n84, n85,
         n86, n87, n88;
  wire   [4:0] sel;

  NAND3_X1 U110 ( .A1(sel[1]), .A2(n87), .A3(sel[2]), .ZN(n81) );
  SHIFTER_GENERIC_N32_DW_sra_0 sra_28 ( .A(A), .SH({n85, B[3:0]}), .SH_TC(1'b0), .B({N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82}) );
  SHIFTER_GENERIC_N32_DW_rash_0 srl_26 ( .A(A), .DATA_TC(1'b0), .SH({n85, 
        B[3:0]}), .SH_TC(1'b0), .B({N81, N80, N79, N78, N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50}) );
  SHIFTER_GENERIC_N32_DW01_ash_0 sll_27 ( .A(A), .DATA_TC(1'b0), .SH({n85, 
        B[3:0]}), .SH_TC(1'b0), .B({N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18}) );
  BUF_X4 U3 ( .A(B[4]), .Z(n85) );
  AOI22_X1 U4 ( .A1(N87), .A2(n84), .B1(N55), .B2(n12), .ZN(n26) );
  AOI22_X1 U5 ( .A1(N86), .A2(n84), .B1(N54), .B2(n12), .ZN(n28) );
  AOI22_X1 U7 ( .A1(N88), .A2(n84), .B1(N56), .B2(n12), .ZN(n24) );
  AOI22_X1 U8 ( .A1(N91), .A2(n84), .B1(N59), .B2(n12), .ZN(n14) );
  AOI22_X1 U9 ( .A1(N90), .A2(n84), .B1(N58), .B2(n12), .ZN(n20) );
  AOI22_X1 U10 ( .A1(N89), .A2(n84), .B1(N57), .B2(n12), .ZN(n22) );
  AOI22_X1 U11 ( .A1(N110), .A2(n83), .B1(N78), .B2(n11), .ZN(n40) );
  AOI22_X1 U12 ( .A1(N111), .A2(n83), .B1(N79), .B2(n11), .ZN(n38) );
  AOI22_X1 U13 ( .A1(N112), .A2(n83), .B1(N80), .B2(n11), .ZN(n34) );
  AOI22_X1 U14 ( .A1(N104), .A2(n83), .B1(N72), .B2(n11), .ZN(n52) );
  AOI22_X1 U15 ( .A1(N105), .A2(n83), .B1(N73), .B2(n11), .ZN(n50) );
  AOI22_X1 U16 ( .A1(N106), .A2(n83), .B1(N74), .B2(n11), .ZN(n48) );
  AOI22_X1 U17 ( .A1(N107), .A2(n83), .B1(N75), .B2(n11), .ZN(n46) );
  AOI22_X1 U18 ( .A1(N108), .A2(n83), .B1(N76), .B2(n11), .ZN(n44) );
  AOI22_X1 U19 ( .A1(N95), .A2(n82), .B1(N63), .B2(n10), .ZN(n72) );
  AOI22_X1 U20 ( .A1(N96), .A2(n82), .B1(N64), .B2(n10), .ZN(n70) );
  AOI22_X1 U21 ( .A1(N97), .A2(n82), .B1(N65), .B2(n10), .ZN(n68) );
  AOI22_X1 U22 ( .A1(N93), .A2(n82), .B1(N61), .B2(n10), .ZN(n76) );
  AOI22_X1 U23 ( .A1(N92), .A2(n82), .B1(N60), .B2(n10), .ZN(n78) );
  AOI22_X1 U24 ( .A1(N94), .A2(n82), .B1(N62), .B2(n10), .ZN(n74) );
  AOI22_X1 U25 ( .A1(N99), .A2(n82), .B1(N67), .B2(n10), .ZN(n64) );
  AOI22_X1 U26 ( .A1(N98), .A2(n82), .B1(N66), .B2(n10), .ZN(n66) );
  AOI22_X1 U27 ( .A1(N100), .A2(n82), .B1(N68), .B2(n10), .ZN(n62) );
  AOI22_X1 U28 ( .A1(N102), .A2(n83), .B1(N70), .B2(n11), .ZN(n56) );
  AOI22_X1 U29 ( .A1(N101), .A2(n82), .B1(N69), .B2(n10), .ZN(n60) );
  AOI22_X1 U30 ( .A1(N103), .A2(n83), .B1(N71), .B2(n11), .ZN(n54) );
  NAND2_X1 U31 ( .A1(n57), .A2(n58), .ZN(OUTPUT[1]) );
  AOI22_X1 U32 ( .A1(N83), .A2(n82), .B1(N51), .B2(n10), .ZN(n58) );
  NAND2_X1 U33 ( .A1(n29), .A2(n30), .ZN(OUTPUT[3]) );
  AOI22_X1 U34 ( .A1(N21), .A2(n6), .B1(A[3]), .B2(n3), .ZN(n29) );
  AOI22_X1 U35 ( .A1(N85), .A2(n84), .B1(N53), .B2(n12), .ZN(n30) );
  NAND2_X1 U36 ( .A1(n79), .A2(n80), .ZN(OUTPUT[0]) );
  AOI22_X1 U37 ( .A1(N18), .A2(n4), .B1(A[0]), .B2(n1), .ZN(n79) );
  AOI22_X1 U38 ( .A1(N82), .A2(n82), .B1(N50), .B2(n10), .ZN(n80) );
  AOI22_X1 U39 ( .A1(N25), .A2(n6), .B1(A[7]), .B2(n3), .ZN(n21) );
  AOI22_X1 U40 ( .A1(N24), .A2(n6), .B1(A[6]), .B2(n3), .ZN(n23) );
  AOI22_X1 U41 ( .A1(N30), .A2(n4), .B1(A[12]), .B2(n1), .ZN(n73) );
  AOI22_X1 U42 ( .A1(N32), .A2(n4), .B1(A[14]), .B2(n1), .ZN(n69) );
  AOI22_X1 U43 ( .A1(N35), .A2(n4), .B1(A[17]), .B2(n1), .ZN(n63) );
  AOI22_X1 U44 ( .A1(N31), .A2(n4), .B1(A[13]), .B2(n1), .ZN(n71) );
  AOI22_X1 U45 ( .A1(N33), .A2(n4), .B1(A[15]), .B2(n1), .ZN(n67) );
  AOI22_X1 U46 ( .A1(N34), .A2(n4), .B1(A[16]), .B2(n1), .ZN(n65) );
  AOI22_X1 U47 ( .A1(N45), .A2(n5), .B1(A[27]), .B2(n2), .ZN(n41) );
  AOI22_X1 U48 ( .A1(N44), .A2(n5), .B1(A[26]), .B2(n2), .ZN(n43) );
  AOI22_X1 U49 ( .A1(N49), .A2(n6), .B1(A[31]), .B2(n3), .ZN(n31) );
  AOI22_X1 U50 ( .A1(N46), .A2(n5), .B1(A[28]), .B2(n2), .ZN(n39) );
  AOI22_X1 U51 ( .A1(N36), .A2(n4), .B1(A[18]), .B2(n1), .ZN(n61) );
  AOI22_X1 U52 ( .A1(N113), .A2(n84), .B1(N81), .B2(n12), .ZN(n32) );
  AOI22_X1 U53 ( .A1(N47), .A2(n5), .B1(A[29]), .B2(n2), .ZN(n37) );
  BUF_X1 U54 ( .A(n15), .Z(n82) );
  BUF_X1 U55 ( .A(n15), .Z(n83) );
  BUF_X1 U56 ( .A(n16), .Z(n10) );
  BUF_X1 U57 ( .A(n16), .Z(n11) );
  AOI22_X1 U58 ( .A1(N37), .A2(n4), .B1(A[19]), .B2(n1), .ZN(n59) );
  BUF_X1 U59 ( .A(n17), .Z(n4) );
  BUF_X1 U60 ( .A(n17), .Z(n5) );
  BUF_X1 U61 ( .A(n18), .Z(n1) );
  BUF_X1 U62 ( .A(n18), .Z(n2) );
  AOI22_X1 U63 ( .A1(N48), .A2(n5), .B1(A[30]), .B2(n2), .ZN(n33) );
  BUF_X1 U64 ( .A(n15), .Z(n84) );
  BUF_X1 U65 ( .A(n16), .Z(n12) );
  AOI22_X1 U66 ( .A1(N109), .A2(n83), .B1(N77), .B2(n11), .ZN(n42) );
  BUF_X1 U67 ( .A(n17), .Z(n6) );
  AOI22_X1 U68 ( .A1(N26), .A2(n6), .B1(A[8]), .B2(n3), .ZN(n19) );
  AOI22_X1 U69 ( .A1(N27), .A2(n6), .B1(A[9]), .B2(n3), .ZN(n13) );
  BUF_X1 U70 ( .A(n18), .Z(n3) );
  AOI22_X1 U71 ( .A1(N28), .A2(n4), .B1(A[10]), .B2(n1), .ZN(n77) );
  AOI22_X1 U72 ( .A1(N42), .A2(n5), .B1(A[24]), .B2(n2), .ZN(n47) );
  AOI22_X1 U73 ( .A1(N43), .A2(n5), .B1(A[25]), .B2(n2), .ZN(n45) );
  AOI22_X1 U74 ( .A1(N29), .A2(n4), .B1(A[11]), .B2(n1), .ZN(n75) );
  INV_X1 U75 ( .A(n81), .ZN(n86) );
  NAND2_X1 U76 ( .A1(n35), .A2(n36), .ZN(OUTPUT[2]) );
  AOI22_X1 U77 ( .A1(N84), .A2(n83), .B1(N52), .B2(n11), .ZN(n36) );
  AOI22_X1 U78 ( .A1(N39), .A2(n5), .B1(A[21]), .B2(n2), .ZN(n53) );
  AOI22_X1 U79 ( .A1(N38), .A2(n5), .B1(A[20]), .B2(n2), .ZN(n55) );
  AOI22_X1 U80 ( .A1(N40), .A2(n5), .B1(A[22]), .B2(n2), .ZN(n51) );
  AOI22_X1 U81 ( .A1(N41), .A2(n5), .B1(A[23]), .B2(n2), .ZN(n49) );
  NOR3_X1 U82 ( .A1(sel[0]), .A2(sel[3]), .A3(n81), .ZN(n17) );
  INV_X1 U83 ( .A(sel[4]), .ZN(n87) );
  OAI21_X1 U84 ( .B1(sel[0]), .B2(n88), .A(n86), .ZN(n18) );
  INV_X1 U85 ( .A(sel[3]), .ZN(n88) );
  AND3_X1 U86 ( .A1(sel[0]), .A2(n86), .A3(sel[3]), .ZN(n15) );
  AND3_X1 U87 ( .A1(n86), .A2(n88), .A3(sel[0]), .ZN(n16) );
  NAND2_X1 U88 ( .A1(n39), .A2(n40), .ZN(OUTPUT[28]) );
  NAND2_X1 U89 ( .A1(n37), .A2(n38), .ZN(OUTPUT[29]) );
  NAND2_X1 U90 ( .A1(n33), .A2(n34), .ZN(OUTPUT[30]) );
  NAND2_X1 U91 ( .A1(n55), .A2(n56), .ZN(OUTPUT[20]) );
  NAND2_X1 U92 ( .A1(n53), .A2(n54), .ZN(OUTPUT[21]) );
  NAND2_X1 U93 ( .A1(n51), .A2(n52), .ZN(OUTPUT[22]) );
  NAND2_X1 U94 ( .A1(n49), .A2(n50), .ZN(OUTPUT[23]) );
  NAND2_X1 U95 ( .A1(n47), .A2(n48), .ZN(OUTPUT[24]) );
  NAND2_X1 U96 ( .A1(n45), .A2(n46), .ZN(OUTPUT[25]) );
  NAND2_X1 U97 ( .A1(n43), .A2(n44), .ZN(OUTPUT[26]) );
  NAND2_X1 U98 ( .A1(n41), .A2(n42), .ZN(OUTPUT[27]) );
  NAND2_X1 U99 ( .A1(n63), .A2(n64), .ZN(OUTPUT[17]) );
  NAND2_X1 U100 ( .A1(n61), .A2(n62), .ZN(OUTPUT[18]) );
  NAND2_X1 U101 ( .A1(n59), .A2(n60), .ZN(OUTPUT[19]) );
  NAND2_X1 U102 ( .A1(n65), .A2(n66), .ZN(OUTPUT[16]) );
  NAND2_X1 U103 ( .A1(n73), .A2(n74), .ZN(OUTPUT[12]) );
  NAND2_X1 U104 ( .A1(n71), .A2(n72), .ZN(OUTPUT[13]) );
  NAND2_X1 U105 ( .A1(n69), .A2(n70), .ZN(OUTPUT[14]) );
  NAND2_X1 U106 ( .A1(n67), .A2(n68), .ZN(OUTPUT[15]) );
  NAND2_X1 U107 ( .A1(n31), .A2(n32), .ZN(OUTPUT[31]) );
  NAND2_X1 U108 ( .A1(n13), .A2(n14), .ZN(OUTPUT[9]) );
  NAND2_X1 U109 ( .A1(n19), .A2(n20), .ZN(OUTPUT[8]) );
  NAND2_X1 U111 ( .A1(n77), .A2(n78), .ZN(OUTPUT[10]) );
  NAND2_X1 U112 ( .A1(n75), .A2(n76), .ZN(OUTPUT[11]) );
  NAND2_X1 U113 ( .A1(n21), .A2(n22), .ZN(OUTPUT[7]) );
  NAND2_X1 U114 ( .A1(n23), .A2(n24), .ZN(OUTPUT[6]) );
  NAND2_X1 U115 ( .A1(n27), .A2(n28), .ZN(OUTPUT[4]) );
  NAND2_X1 U116 ( .A1(n25), .A2(n26), .ZN(OUTPUT[5]) );
  AOI22_X1 U117 ( .A1(N20), .A2(n5), .B1(A[2]), .B2(n2), .ZN(n35) );
  AOI22_X1 U118 ( .A1(N23), .A2(n6), .B1(A[5]), .B2(n3), .ZN(n25) );
  AOI22_X1 U119 ( .A1(N22), .A2(n6), .B1(A[4]), .B2(n3), .ZN(n27) );
  AOI22_X1 U120 ( .A1(N19), .A2(n4), .B1(A[1]), .B2(n1), .ZN(n57) );
endmodule


module comparator_N32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[0]), .ZN(n2) );
  INV_X1 U2 ( .A(A[1]), .ZN(n3) );
  INV_X1 U3 ( .A(B[1]), .ZN(n1) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n3), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n2), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n1), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n2), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module comparator_N32 ( inA, inB, .op({\op[4] , \op[3] , \op[2] , \op[1] , 
        \op[0] }), res );
  input [31:0] inA;
  input [31:0] inB;
  output [31:0] res;
  input \op[4] , \op[3] , \op[2] , \op[1] , \op[0] ;
  wire   N8, net27627, net27642, net27652, net27653, net27661, net27665,
         net27668, net27736, net27753, net28489, net36280, net36538, net36884,
         net36937, net36956, net36967, net36976, net36998, net37153, net37179,
         net37276, net37323, net37334, net37410, net37531, net37588, net37593,
         net37592, net37658, net37657, net37746, net37745, net38175, net38169,
         net38153, net27641, net27636, net27650, net27647, net27646, net27644,
         net37765, net37406, net36906, net27658, net27657, net27655, net35853,
         net35852, net29761, net27659, net27651, net27649, net27648, net27645,
         net27643, net27640, net27639, net27637, net27635, net27632, net27631,
         net27630, net27629, net27628, net38080, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178;
  wire   [4:0] op;
  assign res[1] = 1'b0;
  assign res[2] = 1'b0;
  assign res[3] = 1'b0;
  assign res[4] = 1'b0;
  assign res[5] = 1'b0;
  assign res[6] = 1'b0;
  assign res[7] = 1'b0;
  assign res[8] = 1'b0;
  assign res[9] = 1'b0;
  assign res[10] = 1'b0;
  assign res[11] = 1'b0;
  assign res[12] = 1'b0;
  assign res[13] = 1'b0;
  assign res[14] = 1'b0;
  assign res[15] = 1'b0;
  assign res[16] = 1'b0;
  assign res[17] = 1'b0;
  assign res[18] = 1'b0;
  assign res[19] = 1'b0;
  assign res[20] = 1'b0;
  assign res[21] = 1'b0;
  assign res[22] = 1'b0;
  assign res[23] = 1'b0;
  assign res[24] = 1'b0;
  assign res[25] = 1'b0;
  assign res[26] = 1'b0;
  assign res[27] = 1'b0;
  assign res[28] = 1'b0;
  assign res[29] = 1'b0;
  assign res[30] = 1'b0;
  assign res[31] = 1'b0;
  assign net28489 = inB[4];
  assign net36998 = inB[3];
  assign net37276 = inA[0];

  comparator_N32_DW01_cmp6_0 r57 ( .A({inA[31:1], net37276}), .B({inB[31:5], 
        net28489, net36998, inB[2:1], net36956}), .TC(1'b0), .EQ(N8) );
  OR2_X2 U2 ( .A1(net37593), .A2(net37334), .ZN(net37592) );
  INV_X1 U3 ( .A(inB[5]), .ZN(n41) );
  OR2_X1 U4 ( .A1(n23), .A2(n108), .ZN(net36976) );
  NAND2_X1 U5 ( .A1(net37153), .A2(net36976), .ZN(n22) );
  INV_X1 U6 ( .A(net36976), .ZN(net37593) );
  NAND2_X1 U7 ( .A1(n16), .A2(n27), .ZN(net37746) );
  INV_X1 U8 ( .A(net37153), .ZN(n16) );
  INV_X1 U10 ( .A(inB[30]), .ZN(n25) );
  INV_X1 U11 ( .A(inB[2]), .ZN(net38175) );
  INV_X1 U12 ( .A(net28489), .ZN(n42) );
  NAND2_X1 U13 ( .A1(n41), .A2(inA[5]), .ZN(net36937) );
  NAND2_X1 U14 ( .A1(inB[28]), .A2(net27668), .ZN(n24) );
  INV_X1 U15 ( .A(inB[29]), .ZN(n21) );
  INV_X1 U16 ( .A(n22), .ZN(net37531) );
  NAND2_X1 U17 ( .A1(n17), .A2(n18), .ZN(net37765) );
  NAND2_X1 U18 ( .A1(net37588), .A2(n4), .ZN(net37406) );
  OAI21_X1 U19 ( .B1(net37765), .B2(net27659), .A(net27658), .ZN(net27639) );
  NAND2_X1 U20 ( .A1(net37323), .A2(n4), .ZN(net36906) );
  AND2_X1 U21 ( .A1(n127), .A2(n128), .ZN(n1) );
  AND2_X1 U22 ( .A1(n125), .A2(n126), .ZN(n2) );
  AND2_X1 U23 ( .A1(n89), .A2(n90), .ZN(n3) );
  AND2_X1 U24 ( .A1(n19), .A2(n20), .ZN(n4) );
  AND2_X1 U25 ( .A1(n102), .A2(n103), .ZN(n5) );
  AND2_X1 U26 ( .A1(net27643), .A2(op[1]), .ZN(n6) );
  AND2_X1 U27 ( .A1(net27643), .A2(op[0]), .ZN(n7) );
  INV_X1 U28 ( .A(n23), .ZN(net36280) );
  OAI211_X1 U29 ( .C1(inA[29]), .C2(n21), .A(n24), .B(net27665), .ZN(n23) );
  AND2_X1 U30 ( .A1(n129), .A2(n130), .ZN(n8) );
  AND2_X1 U31 ( .A1(n69), .A2(n68), .ZN(n9) );
  AND2_X1 U32 ( .A1(n105), .A2(n104), .ZN(n10) );
  AND2_X1 U33 ( .A1(n78), .A2(n79), .ZN(n11) );
  AND2_X1 U34 ( .A1(n100), .A2(n101), .ZN(n12) );
  AND2_X1 U35 ( .A1(n120), .A2(n119), .ZN(n14) );
  AND2_X1 U36 ( .A1(n99), .A2(n98), .ZN(n15) );
  NAND3_X1 U37 ( .A1(net37410), .A2(n27), .A3(net37179), .ZN(net37745) );
  NAND3_X1 U38 ( .A1(inA[29]), .A2(n21), .A3(net27665), .ZN(n20) );
  NAND3_X1 U39 ( .A1(net37410), .A2(net37592), .A3(net37179), .ZN(n18) );
  NAND2_X1 U40 ( .A1(inA[30]), .A2(n25), .ZN(n19) );
  INV_X1 U41 ( .A(inA[30]), .ZN(net27661) );
  BUF_X1 U42 ( .A(net37334), .Z(n27) );
  AND2_X1 U43 ( .A1(net37592), .A2(net37410), .ZN(net37658) );
  NAND2_X1 U44 ( .A1(net37592), .A2(n22), .ZN(n26) );
  AND2_X1 U45 ( .A1(n4), .A2(n26), .ZN(n17) );
  AOI21_X1 U46 ( .B1(n31), .B2(net38080), .A(inB[1]), .ZN(n28) );
  NOR2_X1 U47 ( .A1(n29), .A2(n28), .ZN(net38153) );
  INV_X1 U48 ( .A(inA[1]), .ZN(net38080) );
  OAI22_X1 U49 ( .A1(n32), .A2(net38080), .B1(inB[2]), .B2(net38169), .ZN(n29)
         );
  NOR2_X1 U50 ( .A1(net37276), .A2(n30), .ZN(n31) );
  INV_X1 U51 ( .A(inB[0]), .ZN(n30) );
  NOR2_X1 U52 ( .A1(net37276), .A2(n30), .ZN(n32) );
  OAI211_X1 U53 ( .C1(net27627), .C2(net27628), .A(net27630), .B(net27629), 
        .ZN(res[0]) );
  OAI211_X1 U54 ( .C1(op[0]), .C2(net27643), .A(net27648), .B(net27649), .ZN(
        net27629) );
  NAND2_X1 U55 ( .A1(net36967), .A2(n7), .ZN(net27649) );
  INV_X1 U56 ( .A(N8), .ZN(net27643) );
  NAND2_X1 U57 ( .A1(net36884), .A2(net27643), .ZN(net27632) );
  NOR4_X1 U58 ( .A1(op[1]), .A2(op[2]), .A3(op[4]), .A4(net27651), .ZN(
        net27648) );
  INV_X1 U59 ( .A(op[3]), .ZN(net27651) );
  NAND2_X1 U60 ( .A1(op[4]), .A2(net27651), .ZN(net27627) );
  NOR3_X1 U61 ( .A1(n34), .A2(net27635), .A3(net29761), .ZN(net27630) );
  NOR2_X1 U62 ( .A1(net35852), .A2(net35853), .ZN(net29761) );
  OR3_X1 U63 ( .A1(net27644), .A2(op[4]), .A3(net27640), .ZN(net35853) );
  INV_X1 U64 ( .A(op[1]), .ZN(net27640) );
  NAND2_X1 U65 ( .A1(op[0]), .A2(net27640), .ZN(net27637) );
  NOR2_X1 U66 ( .A1(net27650), .A2(N8), .ZN(net35852) );
  OAI33_X1 U67 ( .A1(net27636), .A2(net27637), .A3(net27632), .B1(n33), .B2(
        op[0]), .B3(net27636), .ZN(net27635) );
  AOI21_X1 U68 ( .B1(net27639), .B2(op[1]), .A(N8), .ZN(n33) );
  INV_X1 U69 ( .A(net27657), .ZN(net27659) );
  OAI21_X1 U70 ( .B1(net36906), .B2(net27659), .A(net27658), .ZN(net36884) );
  AND2_X1 U71 ( .A1(net27632), .A2(net27631), .ZN(n34) );
  NOR3_X1 U72 ( .A1(net27644), .A2(op[1]), .A3(net27645), .ZN(net27631) );
  INV_X1 U73 ( .A(op[4]), .ZN(net27645) );
  NAND3_X1 U74 ( .A1(net27652), .A2(net27653), .A3(n6), .ZN(net27628) );
  NAND2_X1 U75 ( .A1(inB[31]), .A2(n35), .ZN(net27658) );
  INV_X1 U76 ( .A(net27658), .ZN(net27655) );
  INV_X1 U77 ( .A(inA[31]), .ZN(n35) );
  NAND2_X1 U78 ( .A1(inA[31]), .A2(n36), .ZN(net27657) );
  OAI21_X1 U79 ( .B1(net37406), .B2(net27655), .A(net27657), .ZN(net27650) );
  OAI21_X1 U80 ( .B1(net27655), .B2(net37765), .A(net27657), .ZN(net36967) );
  INV_X1 U81 ( .A(inB[31]), .ZN(n36) );
  NAND3_X1 U82 ( .A1(op[3]), .A2(net27646), .A3(net27647), .ZN(net27644) );
  INV_X1 U83 ( .A(op[2]), .ZN(net27647) );
  INV_X1 U84 ( .A(op[0]), .ZN(net27646) );
  NOR2_X1 U85 ( .A1(op[2]), .A2(net27646), .ZN(n37) );
  OAI21_X1 U86 ( .B1(op[2]), .B2(net27642), .A(net27646), .ZN(net27653) );
  AOI22_X1 U87 ( .A1(op[2]), .A2(net36884), .B1(net27650), .B2(n37), .ZN(
        net27652) );
  NAND2_X1 U88 ( .A1(op[2]), .A2(net27641), .ZN(net27636) );
  INV_X1 U89 ( .A(net27627), .ZN(net27641) );
  NOR2_X1 U90 ( .A1(n38), .A2(net37593), .ZN(net37588) );
  NAND2_X1 U91 ( .A1(net37745), .A2(net37746), .ZN(n38) );
  NAND2_X1 U92 ( .A1(n57), .A2(n55), .ZN(n39) );
  NAND2_X1 U93 ( .A1(n1), .A2(n40), .ZN(n84) );
  NAND2_X1 U94 ( .A1(n124), .A2(n123), .ZN(n40) );
  NAND2_X1 U95 ( .A1(inA[3]), .A2(n48), .ZN(n50) );
  INV_X1 U96 ( .A(net36998), .ZN(n48) );
  NAND2_X1 U97 ( .A1(inB[5]), .A2(n47), .ZN(n43) );
  OAI21_X1 U98 ( .B1(inA[4]), .B2(n42), .A(n43), .ZN(n51) );
  OAI22_X1 U99 ( .A1(inA[2]), .A2(net38175), .B1(inA[3]), .B2(n48), .ZN(n49)
         );
  OAI21_X1 U100 ( .B1(net38153), .B2(n49), .A(n50), .ZN(n44) );
  NOR2_X1 U101 ( .A1(n51), .A2(net36538), .ZN(n46) );
  AOI21_X1 U102 ( .B1(n44), .B2(n45), .A(n46), .ZN(net27736) );
  INV_X1 U103 ( .A(n51), .ZN(n45) );
  INV_X1 U104 ( .A(inA[5]), .ZN(n47) );
  INV_X1 U105 ( .A(inA[4]), .ZN(net27753) );
  INV_X1 U106 ( .A(inA[2]), .ZN(net38169) );
  INV_X1 U107 ( .A(n30), .ZN(net36956) );
  NAND2_X1 U108 ( .A1(n39), .A2(n5), .ZN(n52) );
  AND2_X1 U109 ( .A1(n83), .A2(n75), .ZN(n53) );
  NOR2_X1 U110 ( .A1(n53), .A2(n54), .ZN(net37410) );
  NOR2_X1 U111 ( .A1(n82), .A2(n85), .ZN(n54) );
  AND2_X1 U112 ( .A1(n58), .A2(n9), .ZN(n55) );
  NAND2_X1 U113 ( .A1(n52), .A2(n70), .ZN(n56) );
  AND2_X1 U114 ( .A1(n109), .A2(n84), .ZN(n83) );
  NAND2_X1 U115 ( .A1(n72), .A2(n59), .ZN(n57) );
  OR2_X1 U116 ( .A1(n62), .A2(n3), .ZN(n58) );
  AND2_X1 U117 ( .A1(n64), .A2(n63), .ZN(n59) );
  NAND2_X1 U118 ( .A1(n56), .A2(net37658), .ZN(n60) );
  AND2_X1 U119 ( .A1(n60), .A2(n61), .ZN(net37323) );
  OR2_X1 U120 ( .A1(net37657), .A2(net37531), .ZN(n61) );
  INV_X1 U121 ( .A(net37592), .ZN(net37657) );
  NAND2_X1 U122 ( .A1(n81), .A2(n80), .ZN(n62) );
  INV_X1 U123 ( .A(n62), .ZN(n63) );
  AND2_X1 U124 ( .A1(n71), .A2(n86), .ZN(net37334) );
  AND2_X1 U125 ( .A1(n73), .A2(n10), .ZN(n64) );
  NOR2_X1 U126 ( .A1(n66), .A2(n67), .ZN(n65) );
  NOR2_X1 U127 ( .A1(inA[6]), .A2(n133), .ZN(n66) );
  NOR2_X1 U128 ( .A1(inA[7]), .A2(n134), .ZN(n67) );
  OR2_X1 U129 ( .A1(inB[16]), .A2(n155), .ZN(n68) );
  OR2_X1 U130 ( .A1(inB[15]), .A2(n154), .ZN(n69) );
  NAND2_X1 U131 ( .A1(n52), .A2(n70), .ZN(net37179) );
  AND2_X1 U132 ( .A1(n106), .A2(n83), .ZN(n70) );
  OR2_X1 U133 ( .A1(n76), .A2(n2), .ZN(n71) );
  AND2_X1 U134 ( .A1(n11), .A2(n77), .ZN(net37153) );
  NAND2_X1 U135 ( .A1(n141), .A2(n74), .ZN(n72) );
  OR2_X1 U136 ( .A1(n110), .A2(n87), .ZN(n73) );
  AND2_X1 U137 ( .A1(n14), .A2(n88), .ZN(n74) );
  NAND2_X1 U138 ( .A1(n97), .A2(n96), .ZN(n75) );
  NAND2_X1 U139 ( .A1(n138), .A2(n8), .ZN(n141) );
  NAND2_X1 U140 ( .A1(n92), .A2(n91), .ZN(n76) );
  INV_X1 U141 ( .A(n76), .ZN(n77) );
  OR2_X1 U142 ( .A1(inB[26]), .A2(n175), .ZN(n91) );
  OR2_X1 U143 ( .A1(inB[14]), .A2(n151), .ZN(n89) );
  OR2_X1 U144 ( .A1(inB[24]), .A2(n171), .ZN(n78) );
  OR2_X1 U145 ( .A1(inB[23]), .A2(n170), .ZN(n79) );
  OR2_X1 U146 ( .A1(inA[15]), .A2(n153), .ZN(n80) );
  OR2_X1 U147 ( .A1(inA[14]), .A2(n152), .ZN(n81) );
  INV_X1 U148 ( .A(n84), .ZN(n82) );
  NAND2_X1 U149 ( .A1(n132), .A2(n65), .ZN(n135) );
  AND2_X1 U150 ( .A1(n12), .A2(n1), .ZN(n85) );
  AND2_X1 U151 ( .A1(n15), .A2(net36280), .ZN(n86) );
  NAND2_X1 U152 ( .A1(n95), .A2(n94), .ZN(n87) );
  INV_X1 U153 ( .A(n87), .ZN(n88) );
  OR2_X1 U154 ( .A1(inB[12]), .A2(n147), .ZN(n94) );
  OR2_X1 U155 ( .A1(inB[13]), .A2(n150), .ZN(n90) );
  OR2_X1 U156 ( .A1(inB[25]), .A2(n174), .ZN(n92) );
  OR2_X1 U157 ( .A1(inB[6]), .A2(n131), .ZN(n93) );
  NAND3_X1 U158 ( .A1(net27736), .A2(net36937), .A3(n93), .ZN(n132) );
  OR2_X1 U159 ( .A1(inB[11]), .A2(n146), .ZN(n95) );
  OR2_X1 U160 ( .A1(inA[19]), .A2(n161), .ZN(n96) );
  OR2_X1 U161 ( .A1(inA[18]), .A2(n160), .ZN(n97) );
  OR2_X1 U162 ( .A1(inA[27]), .A2(n177), .ZN(n98) );
  OR2_X1 U163 ( .A1(inA[26]), .A2(n176), .ZN(n99) );
  OR2_X1 U164 ( .A1(inA[21]), .A2(n165), .ZN(n100) );
  OR2_X1 U165 ( .A1(inA[20]), .A2(n164), .ZN(n101) );
  OR2_X1 U166 ( .A1(inA[17]), .A2(n157), .ZN(n102) );
  OR2_X1 U167 ( .A1(inA[16]), .A2(n156), .ZN(n103) );
  OR2_X1 U168 ( .A1(inA[13]), .A2(n149), .ZN(n104) );
  OR2_X1 U169 ( .A1(inA[12]), .A2(n148), .ZN(n105) );
  OR2_X1 U170 ( .A1(net28489), .A2(net27753), .ZN(net36538) );
  AND2_X1 U171 ( .A1(n114), .A2(n113), .ZN(n106) );
  AND2_X1 U172 ( .A1(n116), .A2(n115), .ZN(n107) );
  AND2_X1 U173 ( .A1(n121), .A2(n122), .ZN(n108) );
  AND2_X1 U174 ( .A1(n118), .A2(n117), .ZN(n109) );
  NOR2_X1 U175 ( .A1(n111), .A2(n112), .ZN(n110) );
  NOR2_X1 U176 ( .A1(n144), .A2(inA[10]), .ZN(n111) );
  NOR2_X1 U177 ( .A1(inA[11]), .A2(n145), .ZN(n112) );
  NAND2_X1 U178 ( .A1(n135), .A2(n107), .ZN(n138) );
  OR2_X1 U179 ( .A1(inB[18]), .A2(n159), .ZN(n113) );
  OR2_X1 U180 ( .A1(inB[17]), .A2(n158), .ZN(n114) );
  OR2_X1 U181 ( .A1(inB[8]), .A2(n137), .ZN(n115) );
  OR2_X1 U182 ( .A1(inB[7]), .A2(n136), .ZN(n116) );
  OR2_X1 U183 ( .A1(inB[20]), .A2(n163), .ZN(n117) );
  OR2_X1 U184 ( .A1(inB[19]), .A2(n162), .ZN(n118) );
  OR2_X1 U185 ( .A1(inB[10]), .A2(n143), .ZN(n119) );
  OR2_X1 U186 ( .A1(inB[9]), .A2(n142), .ZN(n120) );
  OR2_X1 U187 ( .A1(inB[28]), .A2(net27668), .ZN(n121) );
  OR2_X1 U188 ( .A1(inB[27]), .A2(n178), .ZN(n122) );
  OR2_X1 U189 ( .A1(inB[22]), .A2(n167), .ZN(n123) );
  OR2_X1 U190 ( .A1(inB[21]), .A2(n166), .ZN(n124) );
  OR2_X1 U191 ( .A1(inA[25]), .A2(n173), .ZN(n125) );
  OR2_X1 U192 ( .A1(inA[24]), .A2(n172), .ZN(n126) );
  OR2_X1 U193 ( .A1(inA[23]), .A2(n169), .ZN(n127) );
  OR2_X1 U194 ( .A1(inA[22]), .A2(n168), .ZN(n128) );
  OR2_X1 U195 ( .A1(inA[9]), .A2(n140), .ZN(n129) );
  OR2_X1 U196 ( .A1(inA[8]), .A2(n139), .ZN(n130) );
  NAND2_X1 U197 ( .A1(inB[30]), .A2(net27661), .ZN(net27665) );
  INV_X1 U198 ( .A(inA[28]), .ZN(net27668) );
  INV_X1 U199 ( .A(inA[27]), .ZN(n178) );
  INV_X1 U200 ( .A(inB[27]), .ZN(n177) );
  INV_X1 U201 ( .A(inB[26]), .ZN(n176) );
  INV_X1 U202 ( .A(inA[26]), .ZN(n175) );
  INV_X1 U203 ( .A(inA[25]), .ZN(n174) );
  INV_X1 U204 ( .A(inB[25]), .ZN(n173) );
  INV_X1 U205 ( .A(inB[24]), .ZN(n172) );
  INV_X1 U206 ( .A(inA[24]), .ZN(n171) );
  INV_X1 U207 ( .A(inA[23]), .ZN(n170) );
  INV_X1 U208 ( .A(inB[23]), .ZN(n169) );
  INV_X1 U209 ( .A(inB[22]), .ZN(n168) );
  INV_X1 U210 ( .A(inA[22]), .ZN(n167) );
  INV_X1 U211 ( .A(inA[21]), .ZN(n166) );
  INV_X1 U212 ( .A(inB[21]), .ZN(n165) );
  INV_X1 U213 ( .A(inB[20]), .ZN(n164) );
  INV_X1 U214 ( .A(inA[20]), .ZN(n163) );
  INV_X1 U215 ( .A(inA[19]), .ZN(n162) );
  INV_X1 U216 ( .A(inB[19]), .ZN(n161) );
  INV_X1 U217 ( .A(inB[18]), .ZN(n160) );
  INV_X1 U218 ( .A(inA[18]), .ZN(n159) );
  INV_X1 U219 ( .A(inA[17]), .ZN(n158) );
  INV_X1 U220 ( .A(inB[17]), .ZN(n157) );
  INV_X1 U221 ( .A(inB[16]), .ZN(n156) );
  INV_X1 U222 ( .A(inA[16]), .ZN(n155) );
  INV_X1 U223 ( .A(inA[15]), .ZN(n154) );
  INV_X1 U224 ( .A(inB[15]), .ZN(n153) );
  INV_X1 U225 ( .A(inB[14]), .ZN(n152) );
  INV_X1 U226 ( .A(inA[14]), .ZN(n151) );
  INV_X1 U227 ( .A(inA[13]), .ZN(n150) );
  INV_X1 U228 ( .A(inB[13]), .ZN(n149) );
  INV_X1 U229 ( .A(inB[12]), .ZN(n148) );
  INV_X1 U230 ( .A(inA[12]), .ZN(n147) );
  INV_X1 U231 ( .A(inA[11]), .ZN(n146) );
  INV_X1 U232 ( .A(inB[11]), .ZN(n145) );
  INV_X1 U233 ( .A(inB[10]), .ZN(n144) );
  INV_X1 U234 ( .A(inA[10]), .ZN(n143) );
  INV_X1 U235 ( .A(inA[9]), .ZN(n142) );
  INV_X1 U236 ( .A(inB[9]), .ZN(n140) );
  INV_X1 U237 ( .A(inB[8]), .ZN(n139) );
  INV_X1 U238 ( .A(inA[8]), .ZN(n137) );
  INV_X1 U239 ( .A(inA[7]), .ZN(n136) );
  INV_X1 U240 ( .A(inB[7]), .ZN(n134) );
  INV_X1 U241 ( .A(inB[6]), .ZN(n133) );
  INV_X1 U242 ( .A(inA[6]), .ZN(n131) );
  INV_X1 U243 ( .A(net36967), .ZN(net27642) );
endmodule


module mux4to1_N32 ( inadd, inlog, insh, incom, .sel({\sel[4] , \sel[3] , 
        \sel[2] , \sel[1] , \sel[0] }), O );
  input [31:0] inadd;
  input [31:0] inlog;
  input [31:0] insh;
  input [31:0] incom;
  output [31:0] O;
  input \sel[4] , \sel[3] , \sel[2] , \sel[1] , \sel[0] ;
  wire   n6, n7, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n28, n29, n50, n51, n68, n69, n70, n71, net27574, net27576, net27607,
         net29471, net29469, net29475, net29479, net29483, net29481, net38998,
         net38995, net39329, net39295, net27572, net39337, net39325, net39320,
         net39318, net39313, net39291, net39286, net39326, net39290, net27618,
         net27616, net27611, net25507, n8, n1, n2, n3, n4, n5, n9, n10, n11,
         n24, n25, n26, n27, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n72, n73,
         n74, n75, n76, n77;
  wire   [4:0] sel;

  NOR2_X1 U2 ( .A1(net39313), .A2(sel[2]), .ZN(net39320) );
  INV_X1 U3 ( .A(sel[3]), .ZN(net39313) );
  INV_X1 U4 ( .A(sel[4]), .ZN(n11) );
  AOI21_X1 U5 ( .B1(net39326), .B2(net25507), .A(sel[4]), .ZN(net39325) );
  AOI21_X1 U6 ( .B1(n33), .B2(net39318), .A(sel[2]), .ZN(n32) );
  INV_X1 U7 ( .A(sel[1]), .ZN(net39318) );
  NOR2_X1 U8 ( .A1(sel[0]), .A2(sel[4]), .ZN(n33) );
  NAND2_X1 U9 ( .A1(sel[1]), .A2(sel[0]), .ZN(net39326) );
  NAND2_X1 U10 ( .A1(sel[3]), .A2(net27611), .ZN(net39290) );
  OAI21_X1 U11 ( .B1(sel[1]), .B2(sel[2]), .A(sel[4]), .ZN(n24) );
  NAND2_X1 U12 ( .A1(inlog[27]), .A2(net29479), .ZN(net38998) );
  NAND2_X1 U13 ( .A1(net39286), .A2(n27), .ZN(n26) );
  NAND2_X1 U14 ( .A1(net39337), .A2(sel[1]), .ZN(n27) );
  OAI21_X1 U15 ( .B1(net39320), .B2(net27611), .A(n11), .ZN(net39337) );
  INV_X1 U16 ( .A(inlog[28]), .ZN(net39329) );
  NAND2_X1 U17 ( .A1(n30), .A2(n31), .ZN(net39291) );
  NOR2_X1 U18 ( .A1(sel[4]), .A2(sel[3]), .ZN(n30) );
  NOR2_X1 U19 ( .A1(net27611), .A2(sel[2]), .ZN(n34) );
  INV_X1 U20 ( .A(sel[2]), .ZN(net25507) );
  AND4_X1 U21 ( .A1(n11), .A2(sel[2]), .A3(sel[1]), .A4(net39290), .ZN(n1) );
  OR2_X1 U22 ( .A1(n37), .A2(net38995), .ZN(n2) );
  AND2_X1 U23 ( .A1(net39326), .A2(n11), .ZN(n3) );
  OR2_X1 U24 ( .A1(net39291), .A2(net39329), .ZN(n4) );
  AND2_X1 U25 ( .A1(net38998), .A2(n26), .ZN(n5) );
  AOI22_X1 U26 ( .A1(incom[0]), .A2(net29471), .B1(insh[0]), .B2(net29483), 
        .ZN(n9) );
  NAND2_X1 U27 ( .A1(n9), .A2(net27607), .ZN(O[0]) );
  BUF_X1 U28 ( .A(n1), .Z(net29483) );
  BUF_X1 U29 ( .A(n1), .Z(net29481) );
  INV_X1 U30 ( .A(sel[0]), .ZN(net27611) );
  BUF_X1 U31 ( .A(n8), .Z(net29471) );
  INV_X1 U32 ( .A(net27616), .ZN(n8) );
  BUF_X1 U33 ( .A(n8), .Z(net29469) );
  MUX2_X1 U34 ( .A(n24), .B(net27618), .S(sel[3]), .Z(net27616) );
  OAI21_X1 U35 ( .B1(n3), .B2(n10), .A(net25507), .ZN(net27618) );
  NOR2_X1 U36 ( .A1(sel[0]), .A2(sel[1]), .ZN(n10) );
  AOI22_X1 U37 ( .A1(inlog[29]), .A2(net29479), .B1(inadd[29]), .B2(net29475), 
        .ZN(n25) );
  NAND2_X1 U38 ( .A1(n25), .A2(net27572), .ZN(O[29]) );
  INV_X2 U39 ( .A(n26), .ZN(net29475) );
  INV_X2 U40 ( .A(net39291), .ZN(net29479) );
  OAI211_X1 U41 ( .C1(n26), .C2(net39295), .A(n4), .B(net27574), .ZN(O[28]) );
  MUX2_X1 U42 ( .A(n32), .B(net39325), .S(sel[3]), .Z(net39286) );
  MUX2_X1 U43 ( .A(sel[2]), .B(n34), .S(sel[1]), .Z(n31) );
  AOI22_X1 U44 ( .A1(incom[29]), .A2(net29471), .B1(insh[29]), .B2(net29483), 
        .ZN(net27572) );
  NOR2_X1 U45 ( .A1(inadd[27]), .A2(n2), .ZN(n36) );
  INV_X1 U46 ( .A(net27576), .ZN(n37) );
  INV_X1 U47 ( .A(net38998), .ZN(net38995) );
  AND2_X1 U48 ( .A1(n5), .A2(net27576), .ZN(n35) );
  NOR2_X1 U49 ( .A1(n35), .A2(n36), .ZN(O[27]) );
  INV_X1 U50 ( .A(inadd[28]), .ZN(net39295) );
  NAND2_X1 U51 ( .A1(n6), .A2(n7), .ZN(O[9]) );
  AOI22_X1 U52 ( .A1(incom[9]), .A2(net29469), .B1(insh[9]), .B2(net29481), 
        .ZN(n7) );
  AOI22_X1 U53 ( .A1(inlog[9]), .A2(net29479), .B1(inadd[9]), .B2(net29475), 
        .ZN(n6) );
  NAND2_X1 U54 ( .A1(n12), .A2(n13), .ZN(O[8]) );
  AOI22_X1 U55 ( .A1(incom[8]), .A2(net29469), .B1(insh[8]), .B2(net29481), 
        .ZN(n13) );
  AOI22_X1 U56 ( .A1(inlog[8]), .A2(net29479), .B1(inadd[8]), .B2(net29475), 
        .ZN(n12) );
  NAND2_X1 U57 ( .A1(n70), .A2(n71), .ZN(O[10]) );
  AOI22_X1 U58 ( .A1(incom[10]), .A2(net29469), .B1(insh[10]), .B2(net29481), 
        .ZN(n71) );
  AOI22_X1 U59 ( .A1(inlog[10]), .A2(net29479), .B1(inadd[10]), .B2(net29475), 
        .ZN(n70) );
  NAND2_X1 U60 ( .A1(n68), .A2(n69), .ZN(O[11]) );
  AOI22_X1 U61 ( .A1(incom[11]), .A2(net29469), .B1(insh[11]), .B2(net29481), 
        .ZN(n69) );
  AOI22_X1 U62 ( .A1(inlog[11]), .A2(net29479), .B1(inadd[11]), .B2(net29475), 
        .ZN(n68) );
  NAND2_X1 U63 ( .A1(n14), .A2(n15), .ZN(O[7]) );
  AOI22_X1 U64 ( .A1(incom[7]), .A2(net29469), .B1(insh[7]), .B2(net29481), 
        .ZN(n15) );
  AOI22_X1 U65 ( .A1(inlog[7]), .A2(net29479), .B1(inadd[7]), .B2(net29475), 
        .ZN(n14) );
  NAND2_X1 U66 ( .A1(n16), .A2(n17), .ZN(O[6]) );
  AOI22_X1 U67 ( .A1(incom[6]), .A2(net29469), .B1(insh[6]), .B2(net29481), 
        .ZN(n17) );
  AOI22_X1 U68 ( .A1(inlog[6]), .A2(net29479), .B1(inadd[6]), .B2(net29475), 
        .ZN(n16) );
  NAND2_X1 U69 ( .A1(n20), .A2(n21), .ZN(O[4]) );
  AOI22_X1 U70 ( .A1(incom[4]), .A2(net29469), .B1(insh[4]), .B2(net29481), 
        .ZN(n21) );
  AOI22_X1 U71 ( .A1(inlog[4]), .A2(net29479), .B1(inadd[4]), .B2(net29475), 
        .ZN(n20) );
  NAND2_X1 U72 ( .A1(n18), .A2(n19), .ZN(O[5]) );
  AOI22_X1 U73 ( .A1(incom[5]), .A2(net29469), .B1(insh[5]), .B2(net29481), 
        .ZN(n19) );
  AOI22_X1 U74 ( .A1(inlog[5]), .A2(net29479), .B1(inadd[5]), .B2(net29475), 
        .ZN(n18) );
  NAND2_X1 U75 ( .A1(n50), .A2(n51), .ZN(O[1]) );
  AOI22_X1 U76 ( .A1(inlog[1]), .A2(net29479), .B1(inadd[1]), .B2(net29475), 
        .ZN(n50) );
  AOI22_X1 U77 ( .A1(incom[1]), .A2(net29469), .B1(insh[1]), .B2(net29481), 
        .ZN(n51) );
  NAND2_X1 U78 ( .A1(n28), .A2(n29), .ZN(O[2]) );
  AOI22_X1 U79 ( .A1(inlog[2]), .A2(net29479), .B1(inadd[2]), .B2(net29475), 
        .ZN(n28) );
  AOI22_X1 U80 ( .A1(incom[2]), .A2(net29469), .B1(insh[2]), .B2(net29481), 
        .ZN(n29) );
  NAND2_X1 U81 ( .A1(n22), .A2(n23), .ZN(O[3]) );
  AOI22_X1 U82 ( .A1(inlog[3]), .A2(net29479), .B1(inadd[3]), .B2(net29475), 
        .ZN(n22) );
  AOI22_X1 U83 ( .A1(incom[3]), .A2(net29469), .B1(insh[3]), .B2(net29481), 
        .ZN(n23) );
  AOI22_X1 U84 ( .A1(inlog[0]), .A2(net29479), .B1(inadd[0]), .B2(net29475), 
        .ZN(net27607) );
  AOI22_X1 U85 ( .A1(inlog[12]), .A2(net29479), .B1(inadd[12]), .B2(net29475), 
        .ZN(n39) );
  AOI22_X1 U86 ( .A1(incom[12]), .A2(net29471), .B1(insh[12]), .B2(net29483), 
        .ZN(n38) );
  NAND2_X1 U87 ( .A1(n39), .A2(n38), .ZN(O[12]) );
  AOI22_X1 U88 ( .A1(inlog[13]), .A2(net29479), .B1(inadd[13]), .B2(net29475), 
        .ZN(n41) );
  AOI22_X1 U89 ( .A1(incom[13]), .A2(net29471), .B1(insh[13]), .B2(net29483), 
        .ZN(n40) );
  NAND2_X1 U90 ( .A1(n41), .A2(n40), .ZN(O[13]) );
  AOI22_X1 U91 ( .A1(inlog[14]), .A2(net29479), .B1(inadd[14]), .B2(net29475), 
        .ZN(n43) );
  AOI22_X1 U92 ( .A1(incom[14]), .A2(net29471), .B1(insh[14]), .B2(net29483), 
        .ZN(n42) );
  NAND2_X1 U93 ( .A1(n43), .A2(n42), .ZN(O[14]) );
  AOI22_X1 U94 ( .A1(inlog[15]), .A2(net29479), .B1(inadd[15]), .B2(net29475), 
        .ZN(n45) );
  AOI22_X1 U95 ( .A1(incom[15]), .A2(net29471), .B1(insh[15]), .B2(net29483), 
        .ZN(n44) );
  NAND2_X1 U96 ( .A1(n45), .A2(n44), .ZN(O[15]) );
  AOI22_X1 U97 ( .A1(inlog[16]), .A2(net29479), .B1(inadd[16]), .B2(net29475), 
        .ZN(n47) );
  AOI22_X1 U98 ( .A1(incom[16]), .A2(net29471), .B1(insh[16]), .B2(net29483), 
        .ZN(n46) );
  NAND2_X1 U99 ( .A1(n47), .A2(n46), .ZN(O[16]) );
  AOI22_X1 U100 ( .A1(inlog[17]), .A2(net29479), .B1(inadd[17]), .B2(net29475), 
        .ZN(n49) );
  AOI22_X1 U101 ( .A1(incom[17]), .A2(net29471), .B1(insh[17]), .B2(net29483), 
        .ZN(n48) );
  NAND2_X1 U102 ( .A1(n49), .A2(n48), .ZN(O[17]) );
  AOI22_X1 U103 ( .A1(inlog[18]), .A2(net29479), .B1(inadd[18]), .B2(net29475), 
        .ZN(n53) );
  AOI22_X1 U104 ( .A1(incom[18]), .A2(net29471), .B1(insh[18]), .B2(net29483), 
        .ZN(n52) );
  NAND2_X1 U105 ( .A1(n53), .A2(n52), .ZN(O[18]) );
  AOI22_X1 U106 ( .A1(inlog[19]), .A2(net29479), .B1(inadd[19]), .B2(net29475), 
        .ZN(n55) );
  AOI22_X1 U107 ( .A1(incom[19]), .A2(net29471), .B1(insh[19]), .B2(net29483), 
        .ZN(n54) );
  NAND2_X1 U108 ( .A1(n55), .A2(n54), .ZN(O[19]) );
  AOI22_X1 U109 ( .A1(inlog[20]), .A2(net29479), .B1(inadd[20]), .B2(net29475), 
        .ZN(n57) );
  AOI22_X1 U110 ( .A1(incom[20]), .A2(net29471), .B1(insh[20]), .B2(net29483), 
        .ZN(n56) );
  NAND2_X1 U111 ( .A1(n57), .A2(n56), .ZN(O[20]) );
  AOI22_X1 U112 ( .A1(inlog[21]), .A2(net29479), .B1(inadd[21]), .B2(net29475), 
        .ZN(n59) );
  AOI22_X1 U113 ( .A1(incom[21]), .A2(net29471), .B1(insh[21]), .B2(net29483), 
        .ZN(n58) );
  NAND2_X1 U114 ( .A1(n59), .A2(n58), .ZN(O[21]) );
  AOI22_X1 U115 ( .A1(inlog[22]), .A2(net29479), .B1(inadd[22]), .B2(net29475), 
        .ZN(n61) );
  AOI22_X1 U116 ( .A1(incom[22]), .A2(net29471), .B1(insh[22]), .B2(net29483), 
        .ZN(n60) );
  NAND2_X1 U117 ( .A1(n61), .A2(n60), .ZN(O[22]) );
  AOI22_X1 U118 ( .A1(inlog[23]), .A2(net29479), .B1(inadd[23]), .B2(net29475), 
        .ZN(n63) );
  AOI22_X1 U119 ( .A1(incom[23]), .A2(net29471), .B1(insh[23]), .B2(net29483), 
        .ZN(n62) );
  NAND2_X1 U120 ( .A1(n63), .A2(n62), .ZN(O[23]) );
  AOI22_X1 U121 ( .A1(inlog[24]), .A2(net29479), .B1(inadd[24]), .B2(net29475), 
        .ZN(n65) );
  AOI22_X1 U122 ( .A1(incom[24]), .A2(net29471), .B1(insh[24]), .B2(net29483), 
        .ZN(n64) );
  NAND2_X1 U123 ( .A1(n65), .A2(n64), .ZN(O[24]) );
  AOI22_X1 U124 ( .A1(inlog[25]), .A2(net29479), .B1(inadd[25]), .B2(net29475), 
        .ZN(n67) );
  AOI22_X1 U125 ( .A1(incom[25]), .A2(net29471), .B1(insh[25]), .B2(net29483), 
        .ZN(n66) );
  NAND2_X1 U126 ( .A1(n67), .A2(n66), .ZN(O[25]) );
  AOI22_X1 U127 ( .A1(inlog[26]), .A2(net29479), .B1(inadd[26]), .B2(net29475), 
        .ZN(n73) );
  AOI22_X1 U128 ( .A1(incom[26]), .A2(net29471), .B1(insh[26]), .B2(net29483), 
        .ZN(n72) );
  NAND2_X1 U129 ( .A1(n73), .A2(n72), .ZN(O[26]) );
  AOI22_X1 U130 ( .A1(incom[27]), .A2(net29471), .B1(insh[27]), .B2(net29483), 
        .ZN(net27576) );
  AOI22_X1 U131 ( .A1(incom[28]), .A2(net29471), .B1(insh[28]), .B2(net29483), 
        .ZN(net27574) );
  AOI22_X1 U132 ( .A1(inlog[30]), .A2(net29479), .B1(inadd[30]), .B2(net29475), 
        .ZN(n75) );
  AOI22_X1 U133 ( .A1(incom[30]), .A2(net29471), .B1(insh[30]), .B2(net29483), 
        .ZN(n74) );
  NAND2_X1 U134 ( .A1(n75), .A2(n74), .ZN(O[30]) );
  AOI22_X1 U135 ( .A1(inlog[31]), .A2(net29479), .B1(inadd[31]), .B2(net29475), 
        .ZN(n77) );
  AOI22_X1 U136 ( .A1(incom[31]), .A2(net29469), .B1(insh[31]), .B2(net29481), 
        .ZN(n76) );
  NAND2_X1 U137 ( .A1(n77), .A2(n76), .ZN(O[31]) );
endmodule


module ALU_N32 ( INA, INB, .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), 
        alu_out );
  input [31:0] INA;
  input [31:0] INB;
  output [31:0] alu_out;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;
  wire   [4:0] OP;
  wire   [31:0] res1;
  wire   [31:0] res2;
  wire   [31:0] res3;
  wire   [31:0] res4;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  add_wrapper_N32 adder ( .A({INA[31], n6, INA[29], n5, INA[27:26], n9, 
        INA[24:22], n12, INA[20:14], n4, n8, n35, n1, INA[9:6], n38, n33, n47, 
        n45, n39, n40}), .B(INB), .SEL({\OP[4] , \OP[3] , \OP[2] , \OP[1] , 
        \OP[0] }), .O(res1) );
  logic_N32 log ( .A({INA[31], n6, INA[29], n5, INA[27:26], n9, INA[24:22], 
        n12, INA[20:14], n4, n8, n35, n1, INA[9:6], n38, n33, n47, n45, n39, 
        n40}), .B({INB[31:22], n15, n13, n29, n32, n30, n10, n21, n18, n2, n23, 
        n28, n25, n20, n41, n27, n42, n22, n26, n31, n44, n19, n43}), .SEL({
        \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), .O(res2) );
  SHIFTER_GENERIC_N32 shifter ( .A({INA[31], n6, INA[29], n5, INA[27:26], n9, 
        INA[24:22], n12, INA[20:14], n4, n8, n35, INA[10:6], n38, n33, n47, 
        n45, n39, n40}), .B({INB[31:22], n15, n13, n29, n32, n30, n10, n21, 
        n18, n2, n23, n28, n25, n20, INB[8], n27, n42, n22, n26, n31, n44, n16, 
        n37}), .sel({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), .OUTPUT(
        res3) );
  comparator_N32 comp ( .inA(INA), .inB({INB[31:22], n15, n13, n29, n32, n30, 
        n10, n21, n18, n2, n23, n28, n25, n20, n41, n27, n42, n22, n26, n3, 
        n24, n16, n17}), .op({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), 
        .res({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, res4[0]}) );
  mux4to1_N32 mux ( .inadd(res1), .inlog(res2), .insh(res3), .incom({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, res4[0]}), .sel({\OP[4] , \OP[3] , 
        \OP[2] , \OP[1] , \OP[0] }), .O(alu_out) );
  BUF_X2 U1 ( .A(INA[1]), .Z(n39) );
  BUF_X2 U2 ( .A(INA[5]), .Z(n38) );
  BUF_X1 U3 ( .A(INA[30]), .Z(n6) );
  BUF_X1 U4 ( .A(INA[4]), .Z(n33) );
  BUF_X1 U5 ( .A(INA[0]), .Z(n40) );
  BUF_X1 U6 ( .A(n24), .Z(n44) );
  CLKBUF_X2 U7 ( .A(INB[1]), .Z(n16) );
  CLKBUF_X1 U8 ( .A(INB[4]), .Z(n26) );
  CLKBUF_X1 U9 ( .A(INA[10]), .Z(n1) );
  CLKBUF_X1 U10 ( .A(INB[13]), .Z(n2) );
  CLKBUF_X1 U11 ( .A(INB[3]), .Z(n3) );
  INV_X2 U12 ( .A(n14), .ZN(n37) );
  BUF_X2 U13 ( .A(INA[13]), .Z(n4) );
  BUF_X2 U14 ( .A(INA[28]), .Z(n5) );
  INV_X1 U15 ( .A(INA[12]), .ZN(n7) );
  INV_X2 U16 ( .A(n7), .ZN(n8) );
  BUF_X2 U17 ( .A(INA[25]), .Z(n9) );
  CLKBUF_X1 U18 ( .A(INB[16]), .Z(n10) );
  INV_X1 U19 ( .A(INA[21]), .ZN(n11) );
  INV_X2 U20 ( .A(n11), .ZN(n12) );
  CLKBUF_X1 U21 ( .A(INB[2]), .Z(n24) );
  CLKBUF_X1 U22 ( .A(INB[20]), .Z(n13) );
  CLKBUF_X1 U23 ( .A(n36), .Z(n14) );
  CLKBUF_X1 U24 ( .A(INB[21]), .Z(n15) );
  CLKBUF_X1 U25 ( .A(INB[5]), .Z(n22) );
  INV_X1 U26 ( .A(n36), .ZN(n17) );
  CLKBUF_X1 U27 ( .A(INB[14]), .Z(n18) );
  CLKBUF_X1 U28 ( .A(n16), .Z(n19) );
  CLKBUF_X1 U29 ( .A(INB[9]), .Z(n20) );
  CLKBUF_X1 U30 ( .A(INB[15]), .Z(n21) );
  CLKBUF_X1 U31 ( .A(INB[12]), .Z(n23) );
  CLKBUF_X1 U32 ( .A(INB[10]), .Z(n25) );
  CLKBUF_X1 U33 ( .A(INB[7]), .Z(n27) );
  CLKBUF_X1 U34 ( .A(INB[11]), .Z(n28) );
  CLKBUF_X1 U35 ( .A(INB[19]), .Z(n29) );
  CLKBUF_X1 U36 ( .A(INB[17]), .Z(n30) );
  CLKBUF_X1 U37 ( .A(n3), .Z(n31) );
  CLKBUF_X1 U38 ( .A(INB[18]), .Z(n32) );
  INV_X1 U39 ( .A(INA[11]), .ZN(n34) );
  INV_X2 U40 ( .A(n34), .ZN(n35) );
  INV_X1 U41 ( .A(INB[0]), .ZN(n36) );
  CLKBUF_X1 U42 ( .A(INB[6]), .Z(n42) );
  CLKBUF_X1 U43 ( .A(INB[8]), .Z(n41) );
  CLKBUF_X1 U44 ( .A(n37), .Z(n43) );
  CLKBUF_X1 U45 ( .A(INA[2]), .Z(n45) );
  INV_X1 U46 ( .A(INA[3]), .ZN(n46) );
  INV_X2 U47 ( .A(n46), .ZN(n47) );
endmodule


module FWD_CAM_1 ( RST, DATA_IN_1, DATA_IN_2, DATA_IN_3, MATCH_1, MATCH_2, 
        MATCH_3 );
  input [5:0] DATA_IN_1;
  input [5:0] DATA_IN_2;
  input [5:0] DATA_IN_3;
  input RST;
  output MATCH_1, MATCH_2, MATCH_3;
  wire   n1, n2, n3, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  NAND3_X1 U27 ( .A1(DATA_IN_3[3]), .A2(n42), .A3(DATA_IN_3[4]), .ZN(n43) );
  NAND3_X1 U28 ( .A1(DATA_IN_2[3]), .A2(n35), .A3(DATA_IN_2[4]), .ZN(n36) );
  NAND3_X1 U29 ( .A1(DATA_IN_1[3]), .A2(n28), .A3(DATA_IN_1[4]), .ZN(n29) );
  AND2_X1 U3 ( .A1(RST), .A2(n31), .ZN(MATCH_1) );
  OAI21_X1 U4 ( .B1(DATA_IN_1[5]), .B2(n30), .A(n29), .ZN(n31) );
  AOI22_X1 U5 ( .A1(n27), .A2(DATA_IN_1[4]), .B1(DATA_IN_1[3]), .B2(n26), .ZN(
        n30) );
  AND2_X1 U6 ( .A1(RST), .A2(n45), .ZN(MATCH_3) );
  OAI21_X1 U7 ( .B1(DATA_IN_3[5]), .B2(n44), .A(n43), .ZN(n45) );
  AND2_X1 U8 ( .A1(RST), .A2(n38), .ZN(MATCH_2) );
  OAI21_X1 U9 ( .B1(DATA_IN_2[5]), .B2(n37), .A(n36), .ZN(n38) );
  AND2_X1 U10 ( .A1(n32), .A2(DATA_IN_2[2]), .ZN(n34) );
  XNOR2_X1 U11 ( .A(DATA_IN_2[2]), .B(n2), .ZN(n35) );
  AND2_X1 U12 ( .A1(n39), .A2(DATA_IN_3[2]), .ZN(n41) );
  XNOR2_X1 U13 ( .A(DATA_IN_3[2]), .B(n1), .ZN(n42) );
  OAI211_X1 U14 ( .C1(DATA_IN_2[4]), .C2(DATA_IN_2[0]), .A(DATA_IN_2[2]), .B(
        DATA_IN_2[1]), .ZN(n33) );
  INV_X1 U15 ( .A(DATA_IN_2[1]), .ZN(n2) );
  OAI211_X1 U16 ( .C1(DATA_IN_3[4]), .C2(DATA_IN_3[0]), .A(DATA_IN_3[2]), .B(
        DATA_IN_3[1]), .ZN(n40) );
  INV_X1 U17 ( .A(DATA_IN_3[1]), .ZN(n1) );
  AOI22_X1 U18 ( .A1(n41), .A2(DATA_IN_3[4]), .B1(DATA_IN_3[3]), .B2(n40), 
        .ZN(n44) );
  OAI22_X1 U19 ( .A1(DATA_IN_3[0]), .A2(DATA_IN_3[1]), .B1(n1), .B2(
        DATA_IN_3[3]), .ZN(n39) );
  INV_X1 U20 ( .A(DATA_IN_1[1]), .ZN(n3) );
  OAI22_X1 U21 ( .A1(DATA_IN_1[0]), .A2(DATA_IN_1[1]), .B1(n3), .B2(
        DATA_IN_1[3]), .ZN(n25) );
  AOI22_X1 U22 ( .A1(n34), .A2(DATA_IN_2[4]), .B1(DATA_IN_2[3]), .B2(n33), 
        .ZN(n37) );
  OAI22_X1 U23 ( .A1(DATA_IN_2[0]), .A2(DATA_IN_2[1]), .B1(n2), .B2(
        DATA_IN_2[3]), .ZN(n32) );
  AND2_X1 U24 ( .A1(n25), .A2(DATA_IN_1[2]), .ZN(n27) );
  OAI211_X1 U25 ( .C1(DATA_IN_1[4]), .C2(DATA_IN_1[0]), .A(DATA_IN_1[2]), .B(
        DATA_IN_1[1]), .ZN(n26) );
  XNOR2_X1 U26 ( .A(DATA_IN_1[2]), .B(n3), .ZN(n28) );
endmodule


module FWD_UNIT_BRANCH ( Rst, Rs1, Rd_M, Rd_W, ICODE, ICODE_M, ICODE_W, SEL );
  input [4:0] Rs1;
  input [4:0] Rd_M;
  input [4:0] Rd_W;
  input [5:0] ICODE;
  input [5:0] ICODE_M;
  input [5:0] ICODE_W;
  output [1:0] SEL;
  input Rst;
  wire   match_op_M, match_op_W, N12, N13, N14, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27;

  DLH_X1 \SEL_reg[1]  ( .G(N12), .D(N14), .Q(SEL[1]) );
  DLH_X1 \SEL_reg[0]  ( .G(N12), .D(N13), .Q(SEL[0]) );
  FWD_CAM_1 CAM ( .RST(Rst), .DATA_IN_1(ICODE), .DATA_IN_2(ICODE_M), 
        .DATA_IN_3(ICODE_W), .MATCH_2(match_op_M), .MATCH_3(match_op_W) );
  INV_X1 U3 ( .A(Rst), .ZN(n1) );
  NOR4_X1 U4 ( .A1(n2), .A2(n3), .A3(n1), .A4(n4), .ZN(N14) );
  XOR2_X1 U5 ( .A(Rs1[3]), .B(Rd_W[3]), .Z(n4) );
  OAI221_X1 U6 ( .B1(match_op_W), .B2(n5), .C1(n6), .C2(n7), .A(n8), .ZN(n3)
         );
  OR2_X1 U7 ( .A1(Rd_W[0]), .A2(Rd_W[1]), .ZN(n7) );
  OR3_X1 U8 ( .A1(Rd_W[3]), .A2(Rd_W[4]), .A3(Rd_W[2]), .ZN(n6) );
  NOR4_X1 U9 ( .A1(n9), .A2(ICODE_W[0]), .A3(ICODE_W[2]), .A4(ICODE_W[1]), 
        .ZN(n5) );
  OR3_X1 U10 ( .A1(ICODE_W[5]), .A2(ICODE_W[4]), .A3(ICODE_W[3]), .ZN(n9) );
  NAND4_X1 U11 ( .A1(n10), .A2(n11), .A3(n12), .A4(n13), .ZN(n2) );
  XNOR2_X1 U12 ( .A(Rd_W[0]), .B(Rs1[0]), .ZN(n13) );
  XNOR2_X1 U13 ( .A(Rd_W[1]), .B(Rs1[1]), .ZN(n12) );
  XNOR2_X1 U14 ( .A(Rd_W[2]), .B(Rs1[2]), .ZN(n11) );
  XOR2_X1 U15 ( .A(Rd_W[4]), .B(n14), .Z(n10) );
  NOR2_X1 U16 ( .A1(n1), .A2(n8), .ZN(N13) );
  OR4_X1 U17 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n8) );
  OAI211_X1 U18 ( .C1(match_op_M), .C2(n19), .A(n20), .B(n21), .ZN(n18) );
  XNOR2_X1 U19 ( .A(Rd_M[0]), .B(Rs1[0]), .ZN(n21) );
  XNOR2_X1 U20 ( .A(Rd_M[1]), .B(Rs1[1]), .ZN(n20) );
  NOR4_X1 U21 ( .A1(n22), .A2(ICODE_M[0]), .A3(ICODE_M[2]), .A4(ICODE_M[1]), 
        .ZN(n19) );
  OR3_X1 U22 ( .A1(ICODE_M[5]), .A2(ICODE_M[4]), .A3(ICODE_M[3]), .ZN(n22) );
  MUX2_X1 U23 ( .A(n23), .B(n14), .S(Rd_M[4]), .Z(n17) );
  NAND2_X1 U24 ( .A1(n14), .A2(n24), .ZN(n23) );
  OR4_X1 U25 ( .A1(Rd_M[0]), .A2(Rd_M[1]), .A3(Rd_M[2]), .A4(Rd_M[3]), .ZN(n24) );
  INV_X1 U26 ( .A(Rs1[4]), .ZN(n14) );
  XOR2_X1 U27 ( .A(Rs1[3]), .B(Rd_M[3]), .Z(n16) );
  XOR2_X1 U28 ( .A(Rs1[2]), .B(Rd_M[2]), .Z(n15) );
  NAND2_X1 U29 ( .A1(Rst), .A2(n25), .ZN(N12) );
  NAND3_X1 U30 ( .A1(ICODE[2]), .A2(n26), .A3(n27), .ZN(n25) );
  NOR3_X1 U31 ( .A1(ICODE[3]), .A2(ICODE[5]), .A3(ICODE[4]), .ZN(n27) );
  INV_X1 U32 ( .A(ICODE[1]), .ZN(n26) );
endmodule


module mux_3to1_N32_2 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;

  BUF_X1 U1 ( .A(n109), .Z(n1) );
  BUF_X1 U2 ( .A(n109), .Z(n2) );
  BUF_X1 U3 ( .A(n109), .Z(n3) );
  NOR2_X1 U4 ( .A1(n6), .A2(n7), .ZN(n109) );
  INV_X1 U5 ( .A(n93), .ZN(Y[23]) );
  INV_X1 U6 ( .A(n92), .ZN(Y[22]) );
  INV_X1 U7 ( .A(n91), .ZN(Y[21]) );
  INV_X1 U8 ( .A(n112), .ZN(Y[9]) );
  INV_X1 U9 ( .A(n108), .ZN(Y[8]) );
  INV_X1 U10 ( .A(n107), .ZN(Y[7]) );
  INV_X1 U11 ( .A(n89), .ZN(Y[1]) );
  INV_X1 U12 ( .A(n88), .ZN(Y[19]) );
  INV_X1 U13 ( .A(n87), .ZN(Y[18]) );
  INV_X1 U14 ( .A(n105), .ZN(Y[5]) );
  INV_X1 U15 ( .A(n104), .ZN(Y[4]) );
  INV_X1 U16 ( .A(n103), .ZN(Y[3]) );
  INV_X1 U17 ( .A(n85), .ZN(Y[16]) );
  INV_X1 U18 ( .A(n84), .ZN(Y[15]) );
  INV_X1 U19 ( .A(n83), .ZN(Y[14]) );
  INV_X1 U20 ( .A(n101), .ZN(Y[30]) );
  INV_X1 U21 ( .A(n100), .ZN(Y[2]) );
  INV_X1 U22 ( .A(n99), .ZN(Y[29]) );
  INV_X1 U23 ( .A(n81), .ZN(Y[12]) );
  INV_X1 U24 ( .A(n80), .ZN(Y[11]) );
  INV_X1 U25 ( .A(n79), .ZN(Y[10]) );
  INV_X1 U26 ( .A(n97), .ZN(Y[27]) );
  INV_X1 U27 ( .A(n96), .ZN(Y[26]) );
  INV_X1 U28 ( .A(n95), .ZN(Y[25]) );
  BUF_X1 U29 ( .A(n110), .Z(n6) );
  BUF_X1 U30 ( .A(n110), .Z(n4) );
  BUF_X1 U31 ( .A(n110), .Z(n5) );
  BUF_X1 U32 ( .A(n111), .Z(n9) );
  BUF_X1 U33 ( .A(n111), .Z(n7) );
  BUF_X1 U34 ( .A(n111), .Z(n8) );
  AOI222_X1 U35 ( .A1(B[14]), .A2(n7), .B1(C[14]), .B2(n6), .C1(A[14]), .C2(n1), .ZN(n83) );
  AOI222_X1 U36 ( .A1(B[15]), .A2(n7), .B1(C[15]), .B2(n6), .C1(A[15]), .C2(n1), .ZN(n84) );
  AOI222_X1 U37 ( .A1(B[16]), .A2(n7), .B1(C[16]), .B2(n6), .C1(A[16]), .C2(n1), .ZN(n85) );
  AOI222_X1 U38 ( .A1(B[10]), .A2(n7), .B1(C[10]), .B2(n6), .C1(A[10]), .C2(n1), .ZN(n79) );
  AOI222_X1 U39 ( .A1(B[11]), .A2(n7), .B1(C[11]), .B2(n6), .C1(A[11]), .C2(n1), .ZN(n80) );
  AOI222_X1 U40 ( .A1(B[12]), .A2(n7), .B1(C[12]), .B2(n6), .C1(A[12]), .C2(n1), .ZN(n81) );
  AOI222_X1 U41 ( .A1(B[21]), .A2(n8), .B1(C[21]), .B2(n5), .C1(A[21]), .C2(n2), .ZN(n91) );
  AOI222_X1 U42 ( .A1(B[22]), .A2(n8), .B1(C[22]), .B2(n5), .C1(A[22]), .C2(n2), .ZN(n92) );
  AOI222_X1 U43 ( .A1(B[23]), .A2(n8), .B1(C[23]), .B2(n5), .C1(A[23]), .C2(n2), .ZN(n93) );
  AOI222_X1 U44 ( .A1(B[18]), .A2(n7), .B1(C[18]), .B2(n5), .C1(A[18]), .C2(n1), .ZN(n87) );
  AOI222_X1 U45 ( .A1(B[19]), .A2(n7), .B1(C[19]), .B2(n5), .C1(A[19]), .C2(n1), .ZN(n88) );
  AOI222_X1 U46 ( .A1(B[1]), .A2(n8), .B1(C[1]), .B2(n5), .C1(A[1]), .C2(n1), 
        .ZN(n89) );
  AOI222_X1 U47 ( .A1(B[7]), .A2(n9), .B1(C[7]), .B2(n4), .C1(A[7]), .C2(n3), 
        .ZN(n107) );
  AOI222_X1 U48 ( .A1(B[8]), .A2(n9), .B1(C[8]), .B2(n4), .C1(A[8]), .C2(n3), 
        .ZN(n108) );
  AOI222_X1 U49 ( .A1(B[9]), .A2(n9), .B1(C[9]), .B2(n4), .C1(A[9]), .C2(n3), 
        .ZN(n112) );
  AOI222_X1 U50 ( .A1(B[3]), .A2(n9), .B1(C[3]), .B2(n4), .C1(A[3]), .C2(n3), 
        .ZN(n103) );
  AOI222_X1 U51 ( .A1(B[4]), .A2(n9), .B1(C[4]), .B2(n4), .C1(A[4]), .C2(n3), 
        .ZN(n104) );
  AOI222_X1 U52 ( .A1(B[5]), .A2(n9), .B1(C[5]), .B2(n4), .C1(A[5]), .C2(n3), 
        .ZN(n105) );
  AOI222_X1 U53 ( .A1(B[29]), .A2(n8), .B1(C[29]), .B2(n4), .C1(A[29]), .C2(n2), .ZN(n99) );
  AOI222_X1 U54 ( .A1(B[2]), .A2(n8), .B1(C[2]), .B2(n4), .C1(A[2]), .C2(n2), 
        .ZN(n100) );
  AOI222_X1 U55 ( .A1(B[30]), .A2(n9), .B1(C[30]), .B2(n4), .C1(A[30]), .C2(n2), .ZN(n101) );
  AOI222_X1 U56 ( .A1(B[25]), .A2(n8), .B1(C[25]), .B2(n5), .C1(A[25]), .C2(n2), .ZN(n95) );
  AOI222_X1 U57 ( .A1(B[26]), .A2(n8), .B1(C[26]), .B2(n5), .C1(A[26]), .C2(n2), .ZN(n96) );
  AOI222_X1 U58 ( .A1(B[27]), .A2(n8), .B1(C[27]), .B2(n5), .C1(A[27]), .C2(n2), .ZN(n97) );
  INV_X1 U59 ( .A(n86), .ZN(Y[17]) );
  AOI222_X1 U60 ( .A1(B[17]), .A2(n7), .B1(C[17]), .B2(n5), .C1(A[17]), .C2(n1), .ZN(n86) );
  INV_X1 U61 ( .A(n98), .ZN(Y[28]) );
  AOI222_X1 U62 ( .A1(B[28]), .A2(n8), .B1(C[28]), .B2(n4), .C1(A[28]), .C2(n2), .ZN(n98) );
  INV_X1 U63 ( .A(n94), .ZN(Y[24]) );
  AOI222_X1 U64 ( .A1(B[24]), .A2(n8), .B1(C[24]), .B2(n5), .C1(A[24]), .C2(n2), .ZN(n94) );
  INV_X1 U65 ( .A(n82), .ZN(Y[13]) );
  AOI222_X1 U66 ( .A1(B[13]), .A2(n7), .B1(C[13]), .B2(n6), .C1(A[13]), .C2(n1), .ZN(n82) );
  INV_X1 U67 ( .A(n78), .ZN(Y[0]) );
  AOI222_X1 U68 ( .A1(B[0]), .A2(n7), .B1(C[0]), .B2(n6), .C1(A[0]), .C2(n1), 
        .ZN(n78) );
  INV_X1 U69 ( .A(n90), .ZN(Y[20]) );
  AOI222_X1 U70 ( .A1(B[20]), .A2(n8), .B1(C[20]), .B2(n5), .C1(A[20]), .C2(n2), .ZN(n90) );
  INV_X1 U71 ( .A(n106), .ZN(Y[6]) );
  AOI222_X1 U72 ( .A1(B[6]), .A2(n9), .B1(C[6]), .B2(n4), .C1(A[6]), .C2(n3), 
        .ZN(n106) );
  INV_X1 U73 ( .A(n102), .ZN(Y[31]) );
  AOI222_X1 U74 ( .A1(B[31]), .A2(n9), .B1(C[31]), .B2(n4), .C1(A[31]), .C2(n3), .ZN(n102) );
  NOR2_X1 U75 ( .A1(n77), .A2(SEL[1]), .ZN(n111) );
  AND2_X1 U76 ( .A1(SEL[1]), .A2(n77), .ZN(n110) );
  INV_X1 U77 ( .A(SEL[0]), .ZN(n77) );
endmodule


module branch_cond_N32 ( A, EN, .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , 
        \OP[0] }), PRE, DISCARD, WRONG, RIGHT, SEL );
  input [31:0] A;
  input EN, \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] , PRE;
  output DISCARD, WRONG, RIGHT, SEL;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n1, n2, n3, n4, n5;
  wire   [4:0] OP;

  NAND3_X1 U29 ( .A1(OP[2]), .A2(n2), .A3(OP[3]), .ZN(n12) );
  NOR2_X1 U3 ( .A1(n5), .A2(n11), .ZN(WRONG) );
  AOI22_X1 U4 ( .A1(n1), .A2(n8), .B1(n9), .B2(n7), .ZN(n11) );
  NOR4_X1 U5 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n19) );
  NOR4_X1 U6 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n23) );
  NOR4_X1 U7 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n18) );
  NOR4_X1 U8 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n22) );
  NOR4_X1 U9 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n17) );
  NOR4_X1 U10 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n21) );
  NOR4_X1 U11 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n16) );
  NOR4_X1 U12 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n20) );
  INV_X1 U13 ( .A(n9), .ZN(n1) );
  OR2_X1 U14 ( .A1(WRONG), .A2(SEL), .ZN(DISCARD) );
  NOR2_X1 U15 ( .A1(n6), .A2(n5), .ZN(RIGHT) );
  AOI22_X1 U16 ( .A1(n7), .A2(n1), .B1(n8), .B2(n9), .ZN(n6) );
  NOR3_X1 U17 ( .A1(n12), .A2(OP[0]), .A3(n3), .ZN(n7) );
  INV_X1 U18 ( .A(OP[4]), .ZN(n2) );
  XNOR2_X1 U19 ( .A(PRE), .B(n13), .ZN(n9) );
  NOR2_X1 U20 ( .A1(n14), .A2(n15), .ZN(n13) );
  NAND4_X1 U21 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n14) );
  NAND4_X1 U22 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n15) );
  INV_X1 U23 ( .A(OP[1]), .ZN(n3) );
  NOR3_X1 U24 ( .A1(n12), .A2(OP[1]), .A3(n4), .ZN(n8) );
  INV_X1 U25 ( .A(OP[0]), .ZN(n4) );
  AND4_X1 U26 ( .A1(OP[4]), .A2(EN), .A3(n10), .A4(n3), .ZN(SEL) );
  NOR2_X1 U27 ( .A1(OP[3]), .A2(OP[2]), .ZN(n10) );
  INV_X1 U28 ( .A(EN), .ZN(n5) );
endmodule


module EX_MEM ( CLK, RST, NPC_IN, NPC_L_IN, ALU_IN, B_IN, RD_IN, OPCODE_IN, 
        NPC_OUT, NPC_L_OUT, ALU_OUT, B_OUT, RD_OUT, OPCODE_OUT );
  input [31:0] NPC_IN;
  input [31:0] NPC_L_IN;
  input [31:0] ALU_IN;
  input [31:0] B_IN;
  input [4:0] RD_IN;
  input [5:0] OPCODE_IN;
  output [31:0] NPC_OUT;
  output [31:0] NPC_L_OUT;
  output [31:0] ALU_OUT;
  output [31:0] B_OUT;
  output [4:0] RD_OUT;
  output [5:0] OPCODE_OUT;
  input CLK, RST;
  wire   n3, n5, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24;

  DFFR_X1 \OPCODE_OUT_reg[5]  ( .D(OPCODE_IN[5]), .CK(CLK), .RN(n13), .Q(
        OPCODE_OUT[5]) );
  DFFR_X1 \OPCODE_OUT_reg[4]  ( .D(OPCODE_IN[4]), .CK(CLK), .RN(n13), .QN(n3)
         );
  DFFR_X1 \OPCODE_OUT_reg[3]  ( .D(OPCODE_IN[3]), .CK(CLK), .RN(n13), .QN(n7)
         );
  DFFR_X1 \OPCODE_OUT_reg[0]  ( .D(OPCODE_IN[0]), .CK(CLK), .RN(n13), .Q(
        OPCODE_OUT[0]) );
  DFFR_X1 \ALU_OUT_reg[31]  ( .D(ALU_IN[31]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[31]) );
  DFFR_X1 \ALU_OUT_reg[30]  ( .D(ALU_IN[30]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[30]) );
  DFFR_X1 \ALU_OUT_reg[29]  ( .D(ALU_IN[29]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[29]) );
  DFFR_X1 \ALU_OUT_reg[28]  ( .D(ALU_IN[28]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[28]) );
  DFFR_X1 \ALU_OUT_reg[27]  ( .D(ALU_IN[27]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[27]) );
  DFFR_X1 \ALU_OUT_reg[26]  ( .D(ALU_IN[26]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[26]) );
  DFFR_X1 \ALU_OUT_reg[25]  ( .D(ALU_IN[25]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[25]) );
  DFFR_X1 \ALU_OUT_reg[24]  ( .D(ALU_IN[24]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[24]) );
  DFFR_X1 \ALU_OUT_reg[23]  ( .D(ALU_IN[23]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[23]) );
  DFFR_X1 \ALU_OUT_reg[22]  ( .D(ALU_IN[22]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[22]) );
  DFFR_X1 \ALU_OUT_reg[21]  ( .D(ALU_IN[21]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[21]) );
  DFFR_X1 \ALU_OUT_reg[20]  ( .D(ALU_IN[20]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[20]) );
  DFFR_X1 \ALU_OUT_reg[19]  ( .D(ALU_IN[19]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[19]) );
  DFFR_X1 \ALU_OUT_reg[18]  ( .D(ALU_IN[18]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[18]) );
  DFFR_X1 \ALU_OUT_reg[17]  ( .D(ALU_IN[17]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[17]) );
  DFFR_X1 \ALU_OUT_reg[16]  ( .D(ALU_IN[16]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[16]) );
  DFFR_X1 \ALU_OUT_reg[15]  ( .D(ALU_IN[15]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[15]) );
  DFFR_X1 \ALU_OUT_reg[14]  ( .D(ALU_IN[14]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[14]) );
  DFFR_X1 \ALU_OUT_reg[13]  ( .D(ALU_IN[13]), .CK(CLK), .RN(n15), .Q(
        ALU_OUT[13]) );
  DFFR_X1 \ALU_OUT_reg[12]  ( .D(ALU_IN[12]), .CK(CLK), .RN(n15), .Q(
        ALU_OUT[12]) );
  DFFR_X1 \ALU_OUT_reg[11]  ( .D(ALU_IN[11]), .CK(CLK), .RN(n15), .Q(
        ALU_OUT[11]) );
  DFFR_X1 \ALU_OUT_reg[10]  ( .D(ALU_IN[10]), .CK(CLK), .RN(n15), .Q(
        ALU_OUT[10]) );
  DFFR_X1 \ALU_OUT_reg[9]  ( .D(ALU_IN[9]), .CK(CLK), .RN(n15), .Q(ALU_OUT[9])
         );
  DFFR_X1 \ALU_OUT_reg[8]  ( .D(ALU_IN[8]), .CK(CLK), .RN(n15), .Q(ALU_OUT[8])
         );
  DFFR_X1 \ALU_OUT_reg[7]  ( .D(ALU_IN[7]), .CK(CLK), .RN(n15), .Q(ALU_OUT[7])
         );
  DFFR_X1 \ALU_OUT_reg[6]  ( .D(ALU_IN[6]), .CK(CLK), .RN(n15), .Q(ALU_OUT[6])
         );
  DFFR_X1 \ALU_OUT_reg[5]  ( .D(ALU_IN[5]), .CK(CLK), .RN(n15), .Q(ALU_OUT[5])
         );
  DFFR_X1 \ALU_OUT_reg[4]  ( .D(ALU_IN[4]), .CK(CLK), .RN(n15), .Q(ALU_OUT[4])
         );
  DFFR_X1 \ALU_OUT_reg[3]  ( .D(ALU_IN[3]), .CK(CLK), .RN(n15), .Q(ALU_OUT[3])
         );
  DFFR_X1 \ALU_OUT_reg[2]  ( .D(ALU_IN[2]), .CK(CLK), .RN(n15), .Q(ALU_OUT[2])
         );
  DFFR_X1 \ALU_OUT_reg[1]  ( .D(ALU_IN[1]), .CK(CLK), .RN(n16), .Q(ALU_OUT[1])
         );
  DFFR_X1 \ALU_OUT_reg[0]  ( .D(ALU_IN[0]), .CK(CLK), .RN(n16), .Q(ALU_OUT[0])
         );
  DFFR_X1 \B_OUT_reg[31]  ( .D(B_IN[31]), .CK(CLK), .RN(n16), .Q(B_OUT[31]) );
  DFFR_X1 \B_OUT_reg[30]  ( .D(B_IN[30]), .CK(CLK), .RN(n16), .Q(B_OUT[30]) );
  DFFR_X1 \B_OUT_reg[29]  ( .D(B_IN[29]), .CK(CLK), .RN(n16), .Q(B_OUT[29]) );
  DFFR_X1 \B_OUT_reg[28]  ( .D(B_IN[28]), .CK(CLK), .RN(n16), .Q(B_OUT[28]) );
  DFFR_X1 \B_OUT_reg[27]  ( .D(B_IN[27]), .CK(CLK), .RN(n16), .Q(B_OUT[27]) );
  DFFR_X1 \B_OUT_reg[26]  ( .D(B_IN[26]), .CK(CLK), .RN(n16), .Q(B_OUT[26]) );
  DFFR_X1 \B_OUT_reg[25]  ( .D(B_IN[25]), .CK(CLK), .RN(n16), .Q(B_OUT[25]) );
  DFFR_X1 \B_OUT_reg[24]  ( .D(B_IN[24]), .CK(CLK), .RN(n16), .Q(B_OUT[24]) );
  DFFR_X1 \B_OUT_reg[23]  ( .D(B_IN[23]), .CK(CLK), .RN(n16), .Q(B_OUT[23]) );
  DFFR_X1 \B_OUT_reg[22]  ( .D(B_IN[22]), .CK(CLK), .RN(n16), .Q(B_OUT[22]) );
  DFFR_X1 \B_OUT_reg[21]  ( .D(B_IN[21]), .CK(CLK), .RN(n17), .Q(B_OUT[21]) );
  DFFR_X1 \B_OUT_reg[20]  ( .D(B_IN[20]), .CK(CLK), .RN(n17), .Q(B_OUT[20]) );
  DFFR_X1 \B_OUT_reg[19]  ( .D(B_IN[19]), .CK(CLK), .RN(n17), .Q(B_OUT[19]) );
  DFFR_X1 \B_OUT_reg[18]  ( .D(B_IN[18]), .CK(CLK), .RN(n17), .Q(B_OUT[18]) );
  DFFR_X1 \B_OUT_reg[17]  ( .D(B_IN[17]), .CK(CLK), .RN(n17), .Q(B_OUT[17]) );
  DFFR_X1 \B_OUT_reg[16]  ( .D(B_IN[16]), .CK(CLK), .RN(n17), .Q(B_OUT[16]) );
  DFFR_X1 \B_OUT_reg[15]  ( .D(B_IN[15]), .CK(CLK), .RN(n17), .Q(B_OUT[15]) );
  DFFR_X1 \B_OUT_reg[14]  ( .D(B_IN[14]), .CK(CLK), .RN(n17), .Q(B_OUT[14]) );
  DFFR_X1 \B_OUT_reg[13]  ( .D(B_IN[13]), .CK(CLK), .RN(n17), .Q(B_OUT[13]) );
  DFFR_X1 \B_OUT_reg[12]  ( .D(B_IN[12]), .CK(CLK), .RN(n17), .Q(B_OUT[12]) );
  DFFR_X1 \B_OUT_reg[11]  ( .D(B_IN[11]), .CK(CLK), .RN(n17), .Q(B_OUT[11]) );
  DFFR_X1 \B_OUT_reg[10]  ( .D(B_IN[10]), .CK(CLK), .RN(n17), .Q(B_OUT[10]) );
  DFFR_X1 \B_OUT_reg[9]  ( .D(B_IN[9]), .CK(CLK), .RN(n18), .Q(B_OUT[9]) );
  DFFR_X1 \B_OUT_reg[8]  ( .D(B_IN[8]), .CK(CLK), .RN(n18), .Q(B_OUT[8]) );
  DFFR_X1 \B_OUT_reg[7]  ( .D(B_IN[7]), .CK(CLK), .RN(n18), .Q(B_OUT[7]) );
  DFFR_X1 \B_OUT_reg[6]  ( .D(B_IN[6]), .CK(CLK), .RN(n18), .Q(B_OUT[6]) );
  DFFR_X1 \B_OUT_reg[5]  ( .D(B_IN[5]), .CK(CLK), .RN(n18), .Q(B_OUT[5]) );
  DFFR_X1 \B_OUT_reg[4]  ( .D(B_IN[4]), .CK(CLK), .RN(n18), .Q(B_OUT[4]) );
  DFFR_X1 \B_OUT_reg[3]  ( .D(B_IN[3]), .CK(CLK), .RN(n18), .Q(B_OUT[3]) );
  DFFR_X1 \B_OUT_reg[2]  ( .D(B_IN[2]), .CK(CLK), .RN(n18), .Q(B_OUT[2]) );
  DFFR_X1 \B_OUT_reg[1]  ( .D(B_IN[1]), .CK(CLK), .RN(n18), .Q(B_OUT[1]) );
  DFFR_X1 \B_OUT_reg[0]  ( .D(B_IN[0]), .CK(CLK), .RN(n18), .Q(B_OUT[0]) );
  DFFR_X1 \NPC_OUT_reg[31]  ( .D(NPC_IN[31]), .CK(CLK), .RN(n18), .Q(
        NPC_OUT[31]) );
  DFFR_X1 \NPC_OUT_reg[30]  ( .D(NPC_IN[30]), .CK(CLK), .RN(n18), .Q(
        NPC_OUT[30]) );
  DFFR_X1 \NPC_OUT_reg[29]  ( .D(NPC_IN[29]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[29]) );
  DFFR_X1 \NPC_OUT_reg[28]  ( .D(NPC_IN[28]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[28]) );
  DFFR_X1 \NPC_OUT_reg[27]  ( .D(NPC_IN[27]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[27]) );
  DFFR_X1 \NPC_OUT_reg[26]  ( .D(NPC_IN[26]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[26]) );
  DFFR_X1 \NPC_OUT_reg[25]  ( .D(NPC_IN[25]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[25]) );
  DFFR_X1 \NPC_OUT_reg[24]  ( .D(NPC_IN[24]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[24]) );
  DFFR_X1 \NPC_OUT_reg[23]  ( .D(NPC_IN[23]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[23]) );
  DFFR_X1 \NPC_OUT_reg[22]  ( .D(NPC_IN[22]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[22]) );
  DFFR_X1 \NPC_OUT_reg[21]  ( .D(NPC_IN[21]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[21]) );
  DFFR_X1 \NPC_OUT_reg[20]  ( .D(NPC_IN[20]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[20]) );
  DFFR_X1 \NPC_OUT_reg[19]  ( .D(NPC_IN[19]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[19]) );
  DFFR_X1 \NPC_OUT_reg[18]  ( .D(NPC_IN[18]), .CK(CLK), .RN(n19), .Q(
        NPC_OUT[18]) );
  DFFR_X1 \NPC_OUT_reg[17]  ( .D(NPC_IN[17]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[17]) );
  DFFR_X1 \NPC_OUT_reg[16]  ( .D(NPC_IN[16]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[16]) );
  DFFR_X1 \NPC_OUT_reg[15]  ( .D(NPC_IN[15]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[15]) );
  DFFR_X1 \NPC_OUT_reg[14]  ( .D(NPC_IN[14]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[14]) );
  DFFR_X1 \NPC_OUT_reg[13]  ( .D(NPC_IN[13]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[13]) );
  DFFR_X1 \NPC_OUT_reg[12]  ( .D(NPC_IN[12]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[12]) );
  DFFR_X1 \NPC_OUT_reg[11]  ( .D(NPC_IN[11]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[11]) );
  DFFR_X1 \NPC_OUT_reg[10]  ( .D(NPC_IN[10]), .CK(CLK), .RN(n20), .Q(
        NPC_OUT[10]) );
  DFFR_X1 \NPC_OUT_reg[9]  ( .D(NPC_IN[9]), .CK(CLK), .RN(n20), .Q(NPC_OUT[9])
         );
  DFFR_X1 \NPC_OUT_reg[8]  ( .D(NPC_IN[8]), .CK(CLK), .RN(n20), .Q(NPC_OUT[8])
         );
  DFFR_X1 \NPC_OUT_reg[7]  ( .D(NPC_IN[7]), .CK(CLK), .RN(n20), .Q(NPC_OUT[7])
         );
  DFFR_X1 \NPC_OUT_reg[6]  ( .D(NPC_IN[6]), .CK(CLK), .RN(n20), .Q(NPC_OUT[6])
         );
  DFFR_X1 \NPC_OUT_reg[5]  ( .D(NPC_IN[5]), .CK(CLK), .RN(n21), .Q(NPC_OUT[5])
         );
  DFFR_X1 \NPC_OUT_reg[4]  ( .D(NPC_IN[4]), .CK(CLK), .RN(n21), .Q(NPC_OUT[4])
         );
  DFFR_X1 \NPC_OUT_reg[3]  ( .D(NPC_IN[3]), .CK(CLK), .RN(n21), .Q(NPC_OUT[3])
         );
  DFFR_X1 \NPC_OUT_reg[2]  ( .D(NPC_IN[2]), .CK(CLK), .RN(n21), .Q(NPC_OUT[2])
         );
  DFFR_X1 \NPC_OUT_reg[1]  ( .D(NPC_IN[1]), .CK(CLK), .RN(n21), .Q(NPC_OUT[1])
         );
  DFFR_X1 \NPC_OUT_reg[0]  ( .D(NPC_IN[0]), .CK(CLK), .RN(n21), .Q(NPC_OUT[0])
         );
  DFFR_X1 \NPC_L_OUT_reg[31]  ( .D(NPC_L_IN[31]), .CK(CLK), .RN(n21), .Q(
        NPC_L_OUT[31]) );
  DFFR_X1 \NPC_L_OUT_reg[30]  ( .D(NPC_L_IN[30]), .CK(CLK), .RN(n21), .Q(
        NPC_L_OUT[30]) );
  DFFR_X1 \NPC_L_OUT_reg[29]  ( .D(NPC_L_IN[29]), .CK(CLK), .RN(n21), .Q(
        NPC_L_OUT[29]) );
  DFFR_X1 \NPC_L_OUT_reg[28]  ( .D(NPC_L_IN[28]), .CK(CLK), .RN(n21), .Q(
        NPC_L_OUT[28]) );
  DFFR_X1 \NPC_L_OUT_reg[27]  ( .D(NPC_L_IN[27]), .CK(CLK), .RN(n21), .Q(
        NPC_L_OUT[27]) );
  DFFR_X1 \NPC_L_OUT_reg[26]  ( .D(NPC_L_IN[26]), .CK(CLK), .RN(n21), .Q(
        NPC_L_OUT[26]) );
  DFFR_X1 \NPC_L_OUT_reg[25]  ( .D(NPC_L_IN[25]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[25]) );
  DFFR_X1 \NPC_L_OUT_reg[24]  ( .D(NPC_L_IN[24]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[24]) );
  DFFR_X1 \NPC_L_OUT_reg[23]  ( .D(NPC_L_IN[23]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[23]) );
  DFFR_X1 \NPC_L_OUT_reg[22]  ( .D(NPC_L_IN[22]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[22]) );
  DFFR_X1 \NPC_L_OUT_reg[21]  ( .D(NPC_L_IN[21]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[21]) );
  DFFR_X1 \NPC_L_OUT_reg[20]  ( .D(NPC_L_IN[20]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[20]) );
  DFFR_X1 \NPC_L_OUT_reg[19]  ( .D(NPC_L_IN[19]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[19]) );
  DFFR_X1 \NPC_L_OUT_reg[18]  ( .D(NPC_L_IN[18]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[18]) );
  DFFR_X1 \NPC_L_OUT_reg[17]  ( .D(NPC_L_IN[17]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[17]) );
  DFFR_X1 \NPC_L_OUT_reg[16]  ( .D(NPC_L_IN[16]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[16]) );
  DFFR_X1 \NPC_L_OUT_reg[15]  ( .D(NPC_L_IN[15]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[15]) );
  DFFR_X1 \NPC_L_OUT_reg[14]  ( .D(NPC_L_IN[14]), .CK(CLK), .RN(n22), .Q(
        NPC_L_OUT[14]) );
  DFFR_X1 \NPC_L_OUT_reg[13]  ( .D(NPC_L_IN[13]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[13]) );
  DFFR_X1 \NPC_L_OUT_reg[12]  ( .D(NPC_L_IN[12]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[12]) );
  DFFR_X1 \NPC_L_OUT_reg[11]  ( .D(NPC_L_IN[11]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[11]) );
  DFFR_X1 \NPC_L_OUT_reg[10]  ( .D(NPC_L_IN[10]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[10]) );
  DFFR_X1 \NPC_L_OUT_reg[9]  ( .D(NPC_L_IN[9]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[9]) );
  DFFR_X1 \NPC_L_OUT_reg[8]  ( .D(NPC_L_IN[8]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[8]) );
  DFFR_X1 \NPC_L_OUT_reg[7]  ( .D(NPC_L_IN[7]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[7]) );
  DFFR_X1 \NPC_L_OUT_reg[6]  ( .D(NPC_L_IN[6]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[6]) );
  DFFR_X1 \NPC_L_OUT_reg[5]  ( .D(NPC_L_IN[5]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[5]) );
  DFFR_X1 \NPC_L_OUT_reg[4]  ( .D(NPC_L_IN[4]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[4]) );
  DFFR_X1 \NPC_L_OUT_reg[3]  ( .D(NPC_L_IN[3]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[3]) );
  DFFR_X1 \NPC_L_OUT_reg[2]  ( .D(NPC_L_IN[2]), .CK(CLK), .RN(n23), .Q(
        NPC_L_OUT[2]) );
  DFFR_X1 \NPC_L_OUT_reg[1]  ( .D(NPC_L_IN[1]), .CK(CLK), .RN(n24), .Q(
        NPC_L_OUT[1]) );
  DFFR_X1 \NPC_L_OUT_reg[0]  ( .D(NPC_L_IN[0]), .CK(CLK), .RN(n24), .Q(
        NPC_L_OUT[0]) );
  DFFR_X1 \RD_OUT_reg[4]  ( .D(RD_IN[4]), .CK(CLK), .RN(n24), .Q(RD_OUT[4]) );
  DFFR_X1 \RD_OUT_reg[3]  ( .D(RD_IN[3]), .CK(CLK), .RN(n24), .Q(RD_OUT[3]) );
  DFFR_X1 \RD_OUT_reg[1]  ( .D(RD_IN[1]), .CK(CLK), .RN(n24), .Q(RD_OUT[1]) );
  DFFR_X1 \RD_OUT_reg[0]  ( .D(RD_IN[0]), .CK(CLK), .RN(n24), .Q(RD_OUT[0]) );
  DFFR_X1 \OPCODE_OUT_reg[1]  ( .D(OPCODE_IN[1]), .CK(CLK), .RN(n13), .QN(n5)
         );
  DFFR_X1 \OPCODE_OUT_reg[2]  ( .D(OPCODE_IN[2]), .CK(CLK), .RN(n13), .QN(n9)
         );
  DFFR_X1 \RD_OUT_reg[2]  ( .D(RD_IN[2]), .CK(CLK), .RN(RST), .Q(RD_OUT[2]) );
  INV_X1 U3 ( .A(n3), .ZN(OPCODE_OUT[4]) );
  INV_X1 U4 ( .A(n5), .ZN(OPCODE_OUT[1]) );
  INV_X1 U5 ( .A(n9), .ZN(OPCODE_OUT[2]) );
  INV_X1 U6 ( .A(n7), .ZN(OPCODE_OUT[3]) );
  BUF_X1 U7 ( .A(RST), .Z(n12) );
  BUF_X1 U8 ( .A(RST), .Z(n11) );
  CLKBUF_X1 U9 ( .A(n11), .Z(n13) );
  CLKBUF_X1 U10 ( .A(n11), .Z(n14) );
  CLKBUF_X1 U11 ( .A(n11), .Z(n15) );
  CLKBUF_X1 U12 ( .A(n11), .Z(n16) );
  CLKBUF_X1 U13 ( .A(n11), .Z(n17) );
  CLKBUF_X1 U14 ( .A(n11), .Z(n18) );
  CLKBUF_X1 U15 ( .A(n12), .Z(n19) );
  CLKBUF_X1 U16 ( .A(n12), .Z(n20) );
  CLKBUF_X1 U17 ( .A(n12), .Z(n21) );
  CLKBUF_X1 U18 ( .A(n12), .Z(n22) );
  CLKBUF_X1 U19 ( .A(n12), .Z(n23) );
  CLKBUF_X1 U20 ( .A(n12), .Z(n24) );
endmodule


module MEM_WB ( CLK, RST, NPC_L_IN, ALU_IN, LMD_IN, RD_IN, OPCODE_IN, 
        NPC_L_OUT, ALU_OUT, LMD_OUT, RD_OUT, OPCODE_OUT );
  input [31:0] NPC_L_IN;
  input [31:0] ALU_IN;
  input [31:0] LMD_IN;
  input [4:0] RD_IN;
  input [5:0] OPCODE_IN;
  output [31:0] NPC_L_OUT;
  output [31:0] ALU_OUT;
  output [31:0] LMD_OUT;
  output [4:0] RD_OUT;
  output [5:0] OPCODE_OUT;
  input CLK, RST;
  wire   n1, n3, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20;

  DFFR_X1 \OPCODE_OUT_reg[5]  ( .D(OPCODE_IN[5]), .CK(CLK), .RN(n12), .Q(
        OPCODE_OUT[5]) );
  DFFR_X1 \OPCODE_OUT_reg[4]  ( .D(OPCODE_IN[4]), .CK(CLK), .RN(n12), .Q(
        OPCODE_OUT[4]) );
  DFFR_X1 \OPCODE_OUT_reg[3]  ( .D(OPCODE_IN[3]), .CK(CLK), .RN(n12), .QN(n7)
         );
  DFFR_X1 \OPCODE_OUT_reg[1]  ( .D(OPCODE_IN[1]), .CK(CLK), .RN(n12), .QN(n1)
         );
  DFFR_X1 \OPCODE_OUT_reg[0]  ( .D(OPCODE_IN[0]), .CK(CLK), .RN(n12), .QN(n3)
         );
  DFFR_X1 \ALU_OUT_reg[31]  ( .D(ALU_IN[31]), .CK(CLK), .RN(n12), .Q(
        ALU_OUT[31]) );
  DFFR_X1 \ALU_OUT_reg[30]  ( .D(ALU_IN[30]), .CK(CLK), .RN(n12), .Q(
        ALU_OUT[30]) );
  DFFR_X1 \ALU_OUT_reg[29]  ( .D(ALU_IN[29]), .CK(CLK), .RN(n12), .Q(
        ALU_OUT[29]) );
  DFFR_X1 \ALU_OUT_reg[28]  ( .D(ALU_IN[28]), .CK(CLK), .RN(n12), .Q(
        ALU_OUT[28]) );
  DFFR_X1 \ALU_OUT_reg[27]  ( .D(ALU_IN[27]), .CK(CLK), .RN(n12), .Q(
        ALU_OUT[27]) );
  DFFR_X1 \ALU_OUT_reg[26]  ( .D(ALU_IN[26]), .CK(CLK), .RN(n12), .Q(
        ALU_OUT[26]) );
  DFFR_X1 \ALU_OUT_reg[25]  ( .D(ALU_IN[25]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[25]) );
  DFFR_X1 \ALU_OUT_reg[24]  ( .D(ALU_IN[24]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[24]) );
  DFFR_X1 \ALU_OUT_reg[23]  ( .D(ALU_IN[23]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[23]) );
  DFFR_X1 \ALU_OUT_reg[22]  ( .D(ALU_IN[22]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[22]) );
  DFFR_X1 \ALU_OUT_reg[21]  ( .D(ALU_IN[21]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[21]) );
  DFFR_X1 \ALU_OUT_reg[20]  ( .D(ALU_IN[20]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[20]) );
  DFFR_X1 \ALU_OUT_reg[19]  ( .D(ALU_IN[19]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[19]) );
  DFFR_X1 \ALU_OUT_reg[18]  ( .D(ALU_IN[18]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[18]) );
  DFFR_X1 \ALU_OUT_reg[17]  ( .D(ALU_IN[17]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[17]) );
  DFFR_X1 \ALU_OUT_reg[16]  ( .D(ALU_IN[16]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[16]) );
  DFFR_X1 \ALU_OUT_reg[15]  ( .D(ALU_IN[15]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[15]) );
  DFFR_X1 \ALU_OUT_reg[14]  ( .D(ALU_IN[14]), .CK(CLK), .RN(n13), .Q(
        ALU_OUT[14]) );
  DFFR_X1 \ALU_OUT_reg[13]  ( .D(ALU_IN[13]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[13]) );
  DFFR_X1 \ALU_OUT_reg[12]  ( .D(ALU_IN[12]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[12]) );
  DFFR_X1 \ALU_OUT_reg[11]  ( .D(ALU_IN[11]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[11]) );
  DFFR_X1 \ALU_OUT_reg[10]  ( .D(ALU_IN[10]), .CK(CLK), .RN(n14), .Q(
        ALU_OUT[10]) );
  DFFR_X1 \ALU_OUT_reg[9]  ( .D(ALU_IN[9]), .CK(CLK), .RN(n14), .Q(ALU_OUT[9])
         );
  DFFR_X1 \ALU_OUT_reg[8]  ( .D(ALU_IN[8]), .CK(CLK), .RN(n14), .Q(ALU_OUT[8])
         );
  DFFR_X1 \ALU_OUT_reg[7]  ( .D(ALU_IN[7]), .CK(CLK), .RN(n14), .Q(ALU_OUT[7])
         );
  DFFR_X1 \ALU_OUT_reg[6]  ( .D(ALU_IN[6]), .CK(CLK), .RN(n14), .Q(ALU_OUT[6])
         );
  DFFR_X1 \ALU_OUT_reg[5]  ( .D(ALU_IN[5]), .CK(CLK), .RN(n14), .Q(ALU_OUT[5])
         );
  DFFR_X1 \ALU_OUT_reg[4]  ( .D(ALU_IN[4]), .CK(CLK), .RN(n14), .Q(ALU_OUT[4])
         );
  DFFR_X1 \ALU_OUT_reg[3]  ( .D(ALU_IN[3]), .CK(CLK), .RN(n14), .Q(ALU_OUT[3])
         );
  DFFR_X1 \ALU_OUT_reg[2]  ( .D(ALU_IN[2]), .CK(CLK), .RN(n14), .Q(ALU_OUT[2])
         );
  DFFR_X1 \ALU_OUT_reg[1]  ( .D(ALU_IN[1]), .CK(CLK), .RN(n15), .Q(ALU_OUT[1])
         );
  DFFR_X1 \ALU_OUT_reg[0]  ( .D(ALU_IN[0]), .CK(CLK), .RN(n15), .Q(ALU_OUT[0])
         );
  DFFR_X1 \LMD_OUT_reg[31]  ( .D(LMD_IN[31]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[31]) );
  DFFR_X1 \LMD_OUT_reg[30]  ( .D(LMD_IN[30]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[30]) );
  DFFR_X1 \LMD_OUT_reg[29]  ( .D(LMD_IN[29]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[29]) );
  DFFR_X1 \LMD_OUT_reg[28]  ( .D(LMD_IN[28]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[28]) );
  DFFR_X1 \LMD_OUT_reg[27]  ( .D(LMD_IN[27]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[27]) );
  DFFR_X1 \LMD_OUT_reg[26]  ( .D(LMD_IN[26]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[26]) );
  DFFR_X1 \LMD_OUT_reg[25]  ( .D(LMD_IN[25]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[25]) );
  DFFR_X1 \LMD_OUT_reg[24]  ( .D(LMD_IN[24]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[24]) );
  DFFR_X1 \LMD_OUT_reg[23]  ( .D(LMD_IN[23]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[23]) );
  DFFR_X1 \LMD_OUT_reg[22]  ( .D(LMD_IN[22]), .CK(CLK), .RN(n15), .Q(
        LMD_OUT[22]) );
  DFFR_X1 \LMD_OUT_reg[21]  ( .D(LMD_IN[21]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[21]) );
  DFFR_X1 \LMD_OUT_reg[20]  ( .D(LMD_IN[20]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[20]) );
  DFFR_X1 \LMD_OUT_reg[19]  ( .D(LMD_IN[19]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[19]) );
  DFFR_X1 \LMD_OUT_reg[18]  ( .D(LMD_IN[18]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[18]) );
  DFFR_X1 \LMD_OUT_reg[17]  ( .D(LMD_IN[17]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[17]) );
  DFFR_X1 \LMD_OUT_reg[16]  ( .D(LMD_IN[16]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[16]) );
  DFFR_X1 \LMD_OUT_reg[15]  ( .D(LMD_IN[15]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[15]) );
  DFFR_X1 \LMD_OUT_reg[14]  ( .D(LMD_IN[14]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[14]) );
  DFFR_X1 \LMD_OUT_reg[13]  ( .D(LMD_IN[13]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[13]) );
  DFFR_X1 \LMD_OUT_reg[12]  ( .D(LMD_IN[12]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[12]) );
  DFFR_X1 \LMD_OUT_reg[11]  ( .D(LMD_IN[11]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[11]) );
  DFFR_X1 \LMD_OUT_reg[10]  ( .D(LMD_IN[10]), .CK(CLK), .RN(n16), .Q(
        LMD_OUT[10]) );
  DFFR_X1 \LMD_OUT_reg[9]  ( .D(LMD_IN[9]), .CK(CLK), .RN(n17), .Q(LMD_OUT[9])
         );
  DFFR_X1 \LMD_OUT_reg[8]  ( .D(LMD_IN[8]), .CK(CLK), .RN(n17), .Q(LMD_OUT[8])
         );
  DFFR_X1 \LMD_OUT_reg[7]  ( .D(LMD_IN[7]), .CK(CLK), .RN(n17), .Q(LMD_OUT[7])
         );
  DFFR_X1 \LMD_OUT_reg[6]  ( .D(LMD_IN[6]), .CK(CLK), .RN(n17), .Q(LMD_OUT[6])
         );
  DFFR_X1 \LMD_OUT_reg[5]  ( .D(LMD_IN[5]), .CK(CLK), .RN(n17), .Q(LMD_OUT[5])
         );
  DFFR_X1 \LMD_OUT_reg[4]  ( .D(LMD_IN[4]), .CK(CLK), .RN(n17), .Q(LMD_OUT[4])
         );
  DFFR_X1 \LMD_OUT_reg[3]  ( .D(LMD_IN[3]), .CK(CLK), .RN(n17), .Q(LMD_OUT[3])
         );
  DFFR_X1 \LMD_OUT_reg[2]  ( .D(LMD_IN[2]), .CK(CLK), .RN(n17), .Q(LMD_OUT[2])
         );
  DFFR_X1 \LMD_OUT_reg[1]  ( .D(LMD_IN[1]), .CK(CLK), .RN(n17), .Q(LMD_OUT[1])
         );
  DFFR_X1 \LMD_OUT_reg[0]  ( .D(LMD_IN[0]), .CK(CLK), .RN(n17), .Q(LMD_OUT[0])
         );
  DFFR_X1 \NPC_L_OUT_reg[31]  ( .D(NPC_L_IN[31]), .CK(CLK), .RN(n17), .Q(
        NPC_L_OUT[31]) );
  DFFR_X1 \NPC_L_OUT_reg[30]  ( .D(NPC_L_IN[30]), .CK(CLK), .RN(n17), .Q(
        NPC_L_OUT[30]) );
  DFFR_X1 \NPC_L_OUT_reg[29]  ( .D(NPC_L_IN[29]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[29]) );
  DFFR_X1 \NPC_L_OUT_reg[28]  ( .D(NPC_L_IN[28]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[28]) );
  DFFR_X1 \NPC_L_OUT_reg[27]  ( .D(NPC_L_IN[27]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[27]) );
  DFFR_X1 \NPC_L_OUT_reg[26]  ( .D(NPC_L_IN[26]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[26]) );
  DFFR_X1 \NPC_L_OUT_reg[25]  ( .D(NPC_L_IN[25]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[25]) );
  DFFR_X1 \NPC_L_OUT_reg[24]  ( .D(NPC_L_IN[24]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[24]) );
  DFFR_X1 \NPC_L_OUT_reg[23]  ( .D(NPC_L_IN[23]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[23]) );
  DFFR_X1 \NPC_L_OUT_reg[22]  ( .D(NPC_L_IN[22]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[22]) );
  DFFR_X1 \NPC_L_OUT_reg[21]  ( .D(NPC_L_IN[21]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[21]) );
  DFFR_X1 \NPC_L_OUT_reg[20]  ( .D(NPC_L_IN[20]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[20]) );
  DFFR_X1 \NPC_L_OUT_reg[19]  ( .D(NPC_L_IN[19]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[19]) );
  DFFR_X1 \NPC_L_OUT_reg[18]  ( .D(NPC_L_IN[18]), .CK(CLK), .RN(n18), .Q(
        NPC_L_OUT[18]) );
  DFFR_X1 \NPC_L_OUT_reg[17]  ( .D(NPC_L_IN[17]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[17]) );
  DFFR_X1 \NPC_L_OUT_reg[16]  ( .D(NPC_L_IN[16]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[16]) );
  DFFR_X1 \NPC_L_OUT_reg[15]  ( .D(NPC_L_IN[15]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[15]) );
  DFFR_X1 \NPC_L_OUT_reg[14]  ( .D(NPC_L_IN[14]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[14]) );
  DFFR_X1 \NPC_L_OUT_reg[13]  ( .D(NPC_L_IN[13]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[13]) );
  DFFR_X1 \NPC_L_OUT_reg[12]  ( .D(NPC_L_IN[12]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[12]) );
  DFFR_X1 \NPC_L_OUT_reg[11]  ( .D(NPC_L_IN[11]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[11]) );
  DFFR_X1 \NPC_L_OUT_reg[10]  ( .D(NPC_L_IN[10]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[10]) );
  DFFR_X1 \NPC_L_OUT_reg[9]  ( .D(NPC_L_IN[9]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[9]) );
  DFFR_X1 \NPC_L_OUT_reg[8]  ( .D(NPC_L_IN[8]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[8]) );
  DFFR_X1 \NPC_L_OUT_reg[7]  ( .D(NPC_L_IN[7]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[7]) );
  DFFR_X1 \NPC_L_OUT_reg[6]  ( .D(NPC_L_IN[6]), .CK(CLK), .RN(n19), .Q(
        NPC_L_OUT[6]) );
  DFFR_X1 \NPC_L_OUT_reg[5]  ( .D(NPC_L_IN[5]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[5]) );
  DFFR_X1 \NPC_L_OUT_reg[4]  ( .D(NPC_L_IN[4]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[4]) );
  DFFR_X1 \NPC_L_OUT_reg[3]  ( .D(NPC_L_IN[3]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[3]) );
  DFFR_X1 \NPC_L_OUT_reg[2]  ( .D(NPC_L_IN[2]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[2]) );
  DFFR_X1 \NPC_L_OUT_reg[1]  ( .D(NPC_L_IN[1]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[1]) );
  DFFR_X1 \NPC_L_OUT_reg[0]  ( .D(NPC_L_IN[0]), .CK(CLK), .RN(n20), .Q(
        NPC_L_OUT[0]) );
  DFFR_X1 \RD_OUT_reg[3]  ( .D(RD_IN[3]), .CK(CLK), .RN(n20), .Q(RD_OUT[3]) );
  DFFR_X1 \RD_OUT_reg[2]  ( .D(RD_IN[2]), .CK(CLK), .RN(n20), .Q(RD_OUT[2]) );
  DFFR_X1 \RD_OUT_reg[0]  ( .D(RD_IN[0]), .CK(CLK), .RN(n20), .Q(RD_OUT[0]) );
  DFFR_X1 \OPCODE_OUT_reg[2]  ( .D(OPCODE_IN[2]), .CK(CLK), .RN(n12), .QN(n5)
         );
  DFFR_X2 \RD_OUT_reg[1]  ( .D(RD_IN[1]), .CK(CLK), .RN(n20), .Q(RD_OUT[1]) );
  DFFR_X2 \RD_OUT_reg[4]  ( .D(RD_IN[4]), .CK(CLK), .RN(n20), .Q(RD_OUT[4]) );
  INV_X1 U3 ( .A(n3), .ZN(OPCODE_OUT[0]) );
  INV_X1 U4 ( .A(n5), .ZN(OPCODE_OUT[2]) );
  INV_X1 U5 ( .A(n1), .ZN(OPCODE_OUT[1]) );
  INV_X1 U6 ( .A(n7), .ZN(OPCODE_OUT[3]) );
  CLKBUF_X1 U7 ( .A(RST), .Z(n9) );
  CLKBUF_X1 U8 ( .A(RST), .Z(n10) );
  CLKBUF_X1 U9 ( .A(RST), .Z(n11) );
  CLKBUF_X1 U10 ( .A(n9), .Z(n12) );
  CLKBUF_X1 U11 ( .A(n9), .Z(n13) );
  CLKBUF_X1 U12 ( .A(n9), .Z(n14) );
  CLKBUF_X1 U13 ( .A(n10), .Z(n15) );
  CLKBUF_X1 U14 ( .A(n10), .Z(n16) );
  CLKBUF_X1 U15 ( .A(n10), .Z(n17) );
  CLKBUF_X1 U16 ( .A(n11), .Z(n18) );
  CLKBUF_X1 U17 ( .A(n11), .Z(n19) );
  CLKBUF_X1 U18 ( .A(n11), .Z(n20) );
endmodule


module mux_3to1_N32_1 ( A, B, C, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;

  BUF_X1 U1 ( .A(n109), .Z(n1) );
  BUF_X1 U2 ( .A(n109), .Z(n2) );
  BUF_X1 U3 ( .A(n109), .Z(n3) );
  NOR2_X1 U4 ( .A1(n6), .A2(n7), .ZN(n109) );
  BUF_X1 U5 ( .A(n110), .Z(n6) );
  BUF_X1 U6 ( .A(n110), .Z(n5) );
  BUF_X1 U7 ( .A(n110), .Z(n4) );
  BUF_X1 U8 ( .A(n111), .Z(n9) );
  BUF_X1 U9 ( .A(n111), .Z(n7) );
  BUF_X1 U10 ( .A(n111), .Z(n8) );
  NOR2_X1 U11 ( .A1(n77), .A2(SEL[1]), .ZN(n111) );
  AND2_X1 U12 ( .A1(SEL[1]), .A2(n77), .ZN(n110) );
  INV_X1 U13 ( .A(n78), .ZN(Y[0]) );
  AOI222_X1 U14 ( .A1(B[0]), .A2(n7), .B1(C[0]), .B2(n6), .C1(A[0]), .C2(n1), 
        .ZN(n78) );
  INV_X1 U15 ( .A(n89), .ZN(Y[1]) );
  AOI222_X1 U16 ( .A1(B[1]), .A2(n8), .B1(C[1]), .B2(n5), .C1(A[1]), .C2(n1), 
        .ZN(n89) );
  INV_X1 U17 ( .A(n100), .ZN(Y[2]) );
  AOI222_X1 U18 ( .A1(B[2]), .A2(n8), .B1(C[2]), .B2(n4), .C1(A[2]), .C2(n2), 
        .ZN(n100) );
  INV_X1 U19 ( .A(n103), .ZN(Y[3]) );
  AOI222_X1 U20 ( .A1(B[3]), .A2(n9), .B1(C[3]), .B2(n4), .C1(A[3]), .C2(n3), 
        .ZN(n103) );
  INV_X1 U21 ( .A(n104), .ZN(Y[4]) );
  AOI222_X1 U22 ( .A1(B[4]), .A2(n9), .B1(C[4]), .B2(n4), .C1(A[4]), .C2(n3), 
        .ZN(n104) );
  INV_X1 U23 ( .A(n105), .ZN(Y[5]) );
  AOI222_X1 U24 ( .A1(B[5]), .A2(n9), .B1(C[5]), .B2(n4), .C1(A[5]), .C2(n3), 
        .ZN(n105) );
  INV_X1 U25 ( .A(n106), .ZN(Y[6]) );
  AOI222_X1 U26 ( .A1(B[6]), .A2(n9), .B1(C[6]), .B2(n4), .C1(A[6]), .C2(n3), 
        .ZN(n106) );
  INV_X1 U27 ( .A(n107), .ZN(Y[7]) );
  AOI222_X1 U28 ( .A1(B[7]), .A2(n9), .B1(C[7]), .B2(n4), .C1(A[7]), .C2(n3), 
        .ZN(n107) );
  INV_X1 U29 ( .A(n108), .ZN(Y[8]) );
  AOI222_X1 U30 ( .A1(B[8]), .A2(n9), .B1(C[8]), .B2(n4), .C1(A[8]), .C2(n3), 
        .ZN(n108) );
  INV_X1 U31 ( .A(n112), .ZN(Y[9]) );
  AOI222_X1 U32 ( .A1(B[9]), .A2(n9), .B1(C[9]), .B2(n4), .C1(A[9]), .C2(n3), 
        .ZN(n112) );
  INV_X1 U33 ( .A(n79), .ZN(Y[10]) );
  AOI222_X1 U34 ( .A1(B[10]), .A2(n7), .B1(C[10]), .B2(n6), .C1(A[10]), .C2(n1), .ZN(n79) );
  INV_X1 U35 ( .A(n80), .ZN(Y[11]) );
  AOI222_X1 U36 ( .A1(B[11]), .A2(n7), .B1(C[11]), .B2(n6), .C1(A[11]), .C2(n1), .ZN(n80) );
  INV_X1 U37 ( .A(n81), .ZN(Y[12]) );
  AOI222_X1 U38 ( .A1(B[12]), .A2(n7), .B1(C[12]), .B2(n6), .C1(A[12]), .C2(n1), .ZN(n81) );
  INV_X1 U39 ( .A(n82), .ZN(Y[13]) );
  AOI222_X1 U40 ( .A1(B[13]), .A2(n7), .B1(C[13]), .B2(n6), .C1(A[13]), .C2(n1), .ZN(n82) );
  INV_X1 U41 ( .A(n83), .ZN(Y[14]) );
  AOI222_X1 U42 ( .A1(B[14]), .A2(n7), .B1(C[14]), .B2(n6), .C1(A[14]), .C2(n1), .ZN(n83) );
  INV_X1 U43 ( .A(n84), .ZN(Y[15]) );
  AOI222_X1 U44 ( .A1(B[15]), .A2(n7), .B1(C[15]), .B2(n6), .C1(A[15]), .C2(n1), .ZN(n84) );
  INV_X1 U45 ( .A(n85), .ZN(Y[16]) );
  AOI222_X1 U46 ( .A1(B[16]), .A2(n7), .B1(C[16]), .B2(n6), .C1(A[16]), .C2(n1), .ZN(n85) );
  INV_X1 U47 ( .A(n86), .ZN(Y[17]) );
  AOI222_X1 U48 ( .A1(B[17]), .A2(n7), .B1(C[17]), .B2(n5), .C1(A[17]), .C2(n1), .ZN(n86) );
  INV_X1 U49 ( .A(n87), .ZN(Y[18]) );
  AOI222_X1 U50 ( .A1(B[18]), .A2(n7), .B1(C[18]), .B2(n5), .C1(A[18]), .C2(n1), .ZN(n87) );
  INV_X1 U51 ( .A(n88), .ZN(Y[19]) );
  AOI222_X1 U52 ( .A1(B[19]), .A2(n7), .B1(C[19]), .B2(n5), .C1(A[19]), .C2(n1), .ZN(n88) );
  INV_X1 U53 ( .A(n90), .ZN(Y[20]) );
  AOI222_X1 U54 ( .A1(B[20]), .A2(n8), .B1(C[20]), .B2(n5), .C1(A[20]), .C2(n2), .ZN(n90) );
  INV_X1 U55 ( .A(n91), .ZN(Y[21]) );
  AOI222_X1 U56 ( .A1(B[21]), .A2(n8), .B1(C[21]), .B2(n5), .C1(A[21]), .C2(n2), .ZN(n91) );
  INV_X1 U57 ( .A(n92), .ZN(Y[22]) );
  AOI222_X1 U58 ( .A1(B[22]), .A2(n8), .B1(C[22]), .B2(n5), .C1(A[22]), .C2(n2), .ZN(n92) );
  INV_X1 U59 ( .A(n93), .ZN(Y[23]) );
  AOI222_X1 U60 ( .A1(B[23]), .A2(n8), .B1(C[23]), .B2(n5), .C1(A[23]), .C2(n2), .ZN(n93) );
  INV_X1 U61 ( .A(n94), .ZN(Y[24]) );
  AOI222_X1 U62 ( .A1(B[24]), .A2(n8), .B1(C[24]), .B2(n5), .C1(A[24]), .C2(n2), .ZN(n94) );
  INV_X1 U63 ( .A(n95), .ZN(Y[25]) );
  AOI222_X1 U64 ( .A1(B[25]), .A2(n8), .B1(C[25]), .B2(n5), .C1(A[25]), .C2(n2), .ZN(n95) );
  INV_X1 U65 ( .A(n96), .ZN(Y[26]) );
  AOI222_X1 U66 ( .A1(B[26]), .A2(n8), .B1(C[26]), .B2(n5), .C1(A[26]), .C2(n2), .ZN(n96) );
  INV_X1 U67 ( .A(n97), .ZN(Y[27]) );
  AOI222_X1 U68 ( .A1(B[27]), .A2(n8), .B1(C[27]), .B2(n5), .C1(A[27]), .C2(n2), .ZN(n97) );
  INV_X1 U69 ( .A(n98), .ZN(Y[28]) );
  AOI222_X1 U70 ( .A1(B[28]), .A2(n8), .B1(C[28]), .B2(n4), .C1(A[28]), .C2(n2), .ZN(n98) );
  INV_X1 U71 ( .A(n99), .ZN(Y[29]) );
  AOI222_X1 U72 ( .A1(B[29]), .A2(n8), .B1(C[29]), .B2(n4), .C1(A[29]), .C2(n2), .ZN(n99) );
  INV_X1 U73 ( .A(n101), .ZN(Y[30]) );
  AOI222_X1 U74 ( .A1(B[30]), .A2(n9), .B1(C[30]), .B2(n4), .C1(A[30]), .C2(n2), .ZN(n101) );
  INV_X1 U75 ( .A(n102), .ZN(Y[31]) );
  AOI222_X1 U76 ( .A1(B[31]), .A2(n9), .B1(C[31]), .B2(n4), .C1(A[31]), .C2(n3), .ZN(n102) );
  INV_X1 U77 ( .A(SEL[0]), .ZN(n77) );
endmodule


module DPATH ( Clk, Rst, MUXA_SEL, MUXB_SEL, BR_EN, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), WB_MUX_SEL, RF_WE, DRAM_OUT, IRAM_OUT, IR1, DRAM_IN, 
        DRAM_ADD, IR_ADD );
  input [1:0] WB_MUX_SEL;
  input [31:0] DRAM_OUT;
  input [31:0] IRAM_OUT;
  output [31:0] IR1;
  output [31:0] DRAM_IN;
  output [11:0] DRAM_ADD;
  output [7:0] IR_ADD;
  input Clk, Rst, MUXA_SEL, MUXB_SEL, BR_EN, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , RF_WE;
  wire   jr_sel, pc_out_1, pc_out_0, wrong_br, right_br, npc_mux_sel,
         prediction, discard_s, pr_D, pr_E, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [4:0] ALU_OPCODE;
  wire   [31:0] alu_out;
  wire   [31:0] npc;
  wire   [31:0] pc_in;
  wire   [31:10] pc_out;
  wire   [31:0] npc_M;
  wire   [15:0] ir_E;
  wire   [31:0] npc_pre;
  wire   [31:0] link_addr_F;
  wire   [31:0] npc_mux_out;
  wire   [31:0] npc_D;
  wire   [31:0] link_addr_D;
  wire   [4:0] add_S1;
  wire   [4:0] add_S2;
  wire   [4:0] dest_D;
  wire   [4:0] add_D;
  wire   [31:0] WB;
  wire   [31:0] a_out;
  wire   [31:0] b_out;
  wire   [31:0] imm_out;
  wire   [31:0] npc_E;
  wire   [31:0] link_addr_E;
  wire   [31:0] A_s;
  wire   [31:0] B_s;
  wire   [31:0] IMM_s;
  wire   [4:0] Rs1;
  wire   [4:0] Rs2;
  wire   [4:0] dest_E;
  wire   [5:0] opcode_E;
  wire   [31:0] mux_a_in;
  wire   [31:0] mux_b_in;
  wire   [4:0] dest_M;
  wire   [5:0] opcode_M;
  wire   [5:0] opcode_W;
  wire   [1:0] FWD_MUX_A_S;
  wire   [1:0] FWD_MUX_B_S;
  wire   [31:12] alu_out_M;
  wire   [31:0] alu_out_W;
  wire   [31:0] alu_a_in;
  wire   [31:0] alu_b_in;
  wire   [1:0] FWD_MUX_BR_S;
  wire   [31:0] br_mux_out;
  wire   [31:0] link_addr_M;
  wire   [31:0] link_addr_W;
  wire   [31:0] LMD_out;

  MUX21_GENERIC_N32_0 NPC_mux ( .A(alu_out), .B(npc), .SEL(jr_sel), .Y(pc_in)
         );
  register_e_N32 PC_reg ( .D(pc_in), .clk(Clk), .rst(n16), .O({pc_out, IR_ADD, 
        pc_out_1, pc_out_0}) );
  branch_predictor BR_pred ( .RST(n16), .PC_IN({pc_out, IR_ADD, pc_out_1, 
        pc_out_0}), .PC_FAIL(npc_M), .IR_IN(IRAM_OUT), .IR_FAIL(ir_E), 
        .WRONG_PRE(wrong_br), .RIGHT_PRE(right_br), .NPC_OUT(npc_pre), 
        .LINK_ADD(link_addr_F), .SEL(npc_mux_sel), .TAKEN(prediction) );
  MUX21_GENERIC_N32_3 NPC_add_mux ( .A(npc_pre), .B({pc_out, IR_ADD, pc_out_1, 
        pc_out_0}), .SEL(npc_mux_sel), .Y(npc_mux_out) );
  NPC_adder NPC_add ( .inPC(npc_mux_out), .outPC(npc) );
  IF_ID IF_IDs ( .CLK(Clk), .RST(n16), .DISCARD(discard_s), .NPC_IN(npc), 
        .NPC_L_IN(link_addr_F), .IR_IN(IRAM_OUT), .PR_IN(prediction), 
        .NPC_OUT(npc_D), .NPC_L_OUT(link_addr_D), .IR_OUT(IR1), .PR_OUT(pr_D)
         );
  IR_decoder dec ( .rst(n16), .IR_OUT(IR1[31:11]), .ADDS1(add_S1), .ADDS2(
        add_S2), .ADDD(dest_D) );
  register_file_N32_addBit5 Reg_F ( .RESET(n16), .RE(1'b1), .WE(RF_WE), 
        .ADD_WR(add_D), .ADD_RDA(add_S1), .ADD_RDB(add_S2), .DATAIN(WB), 
        .OUTA(a_out), .OUTB(b_out) );
  sign_extender sign_ext ( .d_in(IR1), .rst(n16), .d_ext(imm_out) );
  ID_EX ID_EXs ( .CLK(Clk), .RST(n16), .NPC_IN(npc_D), .NPC_L_IN(link_addr_D), 
        .A_IN(a_out), .B_IN(b_out), .IMM_IN(imm_out), .RS1_IN(add_S1), 
        .RS2_IN(add_S2), .RD_IN(dest_D), .OPCODE_IN(IR1[31:26]), .IR_IN(
        IR1[15:0]), .PR_IN(pr_D), .NPC_OUT(npc_E), .NPC_L_OUT(link_addr_E), 
        .A_OUT(A_s), .B_OUT(B_s), .IMM_OUT(IMM_s), .RS1_OUT(Rs1), .RS2_OUT(Rs2), .RD_OUT(dest_E), .OPCODE_OUT(opcode_E), .IR_OUT(ir_E), .PR_OUT(pr_E) );
  MUX21_GENERIC_N32_2 A_mux ( .A(npc_E), .B(A_s), .SEL(MUXA_SEL), .Y(mux_a_in)
         );
  MUX21_GENERIC_N32_1 B_mux ( .A(IMM_s), .B(B_s), .SEL(MUXB_SEL), .Y(mux_b_in)
         );
  FWD_UNIT FORWARDING ( .Rst(n16), .Rs1(Rs1), .Rs2(Rs2), .Rd_M(dest_M), .Rd_W(
        add_D), .ICODE(opcode_E), .ICODE_M(opcode_M), .ICODE_W(opcode_W), 
        .SEL_A(FWD_MUX_A_S), .SEL_B(FWD_MUX_B_S) );
  mux_3to1_N32_0 FWD_MUX_A ( .A(mux_a_in), .B({alu_out_M, DRAM_ADD}), .C(
        alu_out_W), .SEL(FWD_MUX_A_S), .Y(alu_a_in) );
  mux_3to1_N32_3 FWD_MUX_B ( .A(mux_b_in), .B({alu_out_M, DRAM_ADD}), .C(
        alu_out_W), .SEL(FWD_MUX_B_S), .Y(alu_b_in) );
  ALU_N32 ALU_C ( .INA(alu_a_in), .INB(alu_b_in), .OP({\ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), 
        .alu_out(alu_out) );
  FWD_UNIT_BRANCH FORWARDING_BR ( .Rst(n16), .Rs1(Rs1), .Rd_M(dest_M), .Rd_W(
        add_D), .ICODE({opcode_E[5], n9, n3, opcode_E[2], n13, n7}), .ICODE_M(
        {opcode_M[5], n8, n15, n5, n14, n10}), .ICODE_W({opcode_W[5], n11, n6, 
        n4, n12, opcode_W[0]}), .SEL(FWD_MUX_BR_S) );
  mux_3to1_N32_2 FWD_MUX_BRANCH ( .A(A_s), .B({alu_out_M, DRAM_ADD}), .C(
        alu_out_W), .SEL(FWD_MUX_BR_S), .Y(br_mux_out) );
  branch_cond_N32 branch ( .A(br_mux_out), .EN(BR_EN), .OP({\ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , n2, ALU_OPCODE[0]}), .PRE(pr_E), 
        .DISCARD(discard_s), .WRONG(wrong_br), .RIGHT(right_br), .SEL(jr_sel)
         );
  EX_MEM EX_MEM_s ( .CLK(Clk), .RST(n16), .NPC_IN(npc_E), .NPC_L_IN(
        link_addr_E), .ALU_IN({alu_out[31:30], n1, alu_out[28:0]}), .B_IN(B_s), 
        .RD_IN(dest_E), .OPCODE_IN({opcode_E[5], n9, n3, opcode_E[2], n13, n7}), .NPC_OUT(npc_M), .NPC_L_OUT(link_addr_M), .ALU_OUT({alu_out_M, DRAM_ADD}), 
        .B_OUT(DRAM_IN), .RD_OUT(dest_M), .OPCODE_OUT(opcode_M) );
  MEM_WB MEM_WB_s ( .CLK(Clk), .RST(n16), .NPC_L_IN(link_addr_M), .ALU_IN({
        alu_out_M, DRAM_ADD}), .LMD_IN(DRAM_OUT), .RD_IN(dest_M), .OPCODE_IN({
        opcode_M[5:4], n15, n5, n14, n10}), .NPC_L_OUT(link_addr_W), .ALU_OUT(
        alu_out_W), .LMD_OUT(LMD_out), .RD_OUT(add_D), .OPCODE_OUT(opcode_W)
         );
  mux_3to1_N32_1 RF_in_mux ( .A(alu_out_W), .B(LMD_out), .C(link_addr_W), 
        .SEL(WB_MUX_SEL), .Y(WB) );
  CLKBUF_X1 U2 ( .A(alu_out[29]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(ALU_OPCODE[1]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(opcode_E[3]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(opcode_W[2]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(opcode_M[2]), .Z(n5) );
  CLKBUF_X1 U7 ( .A(opcode_W[3]), .Z(n6) );
  CLKBUF_X1 U8 ( .A(opcode_E[0]), .Z(n7) );
  CLKBUF_X1 U9 ( .A(opcode_M[4]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(opcode_E[4]), .Z(n9) );
  BUF_X1 U11 ( .A(Rst), .Z(n16) );
  CLKBUF_X1 U12 ( .A(opcode_M[0]), .Z(n10) );
  CLKBUF_X1 U13 ( .A(opcode_W[4]), .Z(n11) );
  CLKBUF_X1 U14 ( .A(opcode_W[1]), .Z(n12) );
  CLKBUF_X1 U15 ( .A(opcode_E[1]), .Z(n13) );
  CLKBUF_X1 U16 ( .A(opcode_M[1]), .Z(n14) );
  CLKBUF_X1 U17 ( .A(opcode_M[3]), .Z(n15) );
endmodule


module DLX_syn ( Clk, Rst, IRAM_DATA_OUT, DRAM_DATA_OUT, DRAM_DATA_IN, 
        DRAM_ADDRESS, DRAM_ENABLE, DRAM_RW, DRAM_SEL, IRAM_ADDRESS );
  input [31:0] IRAM_DATA_OUT;
  input [31:0] DRAM_DATA_OUT;
  output [31:0] DRAM_DATA_IN;
  output [11:0] DRAM_ADDRESS;
  output [2:0] DRAM_SEL;
  output [7:0] IRAM_ADDRESS;
  input Clk, Rst;
  output DRAM_ENABLE, DRAM_RW;
  wire   IR_CU_31, IR_CU_30, IR_CU_29, IR_CU_28, IR_CU_27, IR_CU_26,
         MUXA_SEL_i, MUXB_SEL_i, BR_EN_i, RF_WE_i;
  wire   [10:0] IR_CU;
  wire   [4:0] ALU_OPCODE_i;
  wire   [1:0] WB_MUX_SEL_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  dlx_cu_MICROCODE_MEM_SIZE63_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE11 CU_I ( 
        .Clk(Clk), .Rst(Rst), .OPCODE_IN({IR_CU_31, IR_CU_30, IR_CU_29, 
        IR_CU_28, IR_CU_27, IR_CU_26}), .FUNC_IN(IR_CU), .MUXA_SEL(MUXA_SEL_i), 
        .MUXB_SEL(MUXB_SEL_i), .BR_EN(BR_EN_i), .ALU_OPCODE(ALU_OPCODE_i), 
        .DRAM_RW(DRAM_RW), .DRAM_EN(DRAM_ENABLE), .DRAM_SEL(DRAM_SEL), 
        .WB_MUX_SEL(WB_MUX_SEL_i), .RF_WE(RF_WE_i) );
  DPATH DataP ( .Clk(Clk), .Rst(Rst), .MUXA_SEL(MUXA_SEL_i), .MUXB_SEL(
        MUXB_SEL_i), .BR_EN(BR_EN_i), .ALU_OPCODE(ALU_OPCODE_i), .WB_MUX_SEL(
        WB_MUX_SEL_i), .RF_WE(RF_WE_i), .DRAM_OUT(DRAM_DATA_OUT), .IRAM_OUT(
        IRAM_DATA_OUT), .IR1({IR_CU_31, IR_CU_30, IR_CU_29, IR_CU_28, IR_CU_27, 
        IR_CU_26, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, IR_CU}), .DRAM_IN(DRAM_DATA_IN), .DRAM_ADD(
        DRAM_ADDRESS), .IR_ADD(IRAM_ADDRESS) );
endmodule

