
module register_file_N32_addBit5 ( RESET, RE, WE, ADD_WR, ADD_RDA, ADD_RDB, 
        DATAIN, OUTA, OUTB );
  input [4:0] ADD_WR;
  input [4:0] ADD_RDA;
  input [4:0] ADD_RDB;
  input [31:0] DATAIN;
  output [31:0] OUTA;
  output [31:0] OUTB;
  input RESET, RE, WE;
  wire   \REGISTERS[1][31] , \REGISTERS[1][30] , \REGISTERS[1][29] ,
         \REGISTERS[1][28] , \REGISTERS[1][27] , \REGISTERS[1][26] ,
         \REGISTERS[1][25] , \REGISTERS[1][24] , \REGISTERS[1][23] ,
         \REGISTERS[1][22] , \REGISTERS[1][21] , \REGISTERS[1][20] ,
         \REGISTERS[1][19] , \REGISTERS[1][18] , \REGISTERS[1][17] ,
         \REGISTERS[1][16] , \REGISTERS[1][15] , \REGISTERS[1][14] ,
         \REGISTERS[1][13] , \REGISTERS[1][12] , \REGISTERS[1][11] ,
         \REGISTERS[1][10] , \REGISTERS[1][9] , \REGISTERS[1][8] ,
         \REGISTERS[1][7] , \REGISTERS[1][6] , \REGISTERS[1][5] ,
         \REGISTERS[1][4] , \REGISTERS[1][3] , \REGISTERS[1][2] ,
         \REGISTERS[1][1] , \REGISTERS[1][0] , \REGISTERS[2][31] ,
         \REGISTERS[2][30] , \REGISTERS[2][29] , \REGISTERS[2][28] ,
         \REGISTERS[2][27] , \REGISTERS[2][26] , \REGISTERS[2][25] ,
         \REGISTERS[2][24] , \REGISTERS[2][23] , \REGISTERS[2][22] ,
         \REGISTERS[2][21] , \REGISTERS[2][20] , \REGISTERS[2][19] ,
         \REGISTERS[2][18] , \REGISTERS[2][17] , \REGISTERS[2][16] ,
         \REGISTERS[2][15] , \REGISTERS[2][14] , \REGISTERS[2][13] ,
         \REGISTERS[2][12] , \REGISTERS[2][11] , \REGISTERS[2][10] ,
         \REGISTERS[2][9] , \REGISTERS[2][8] , \REGISTERS[2][7] ,
         \REGISTERS[2][6] , \REGISTERS[2][5] , \REGISTERS[2][4] ,
         \REGISTERS[2][3] , \REGISTERS[2][2] , \REGISTERS[2][1] ,
         \REGISTERS[2][0] , \REGISTERS[3][31] , \REGISTERS[3][30] ,
         \REGISTERS[3][29] , \REGISTERS[3][28] , \REGISTERS[3][27] ,
         \REGISTERS[3][26] , \REGISTERS[3][25] , \REGISTERS[3][24] ,
         \REGISTERS[3][23] , \REGISTERS[3][22] , \REGISTERS[3][21] ,
         \REGISTERS[3][20] , \REGISTERS[3][19] , \REGISTERS[3][18] ,
         \REGISTERS[3][17] , \REGISTERS[3][16] , \REGISTERS[3][15] ,
         \REGISTERS[3][14] , \REGISTERS[3][13] , \REGISTERS[3][12] ,
         \REGISTERS[3][11] , \REGISTERS[3][10] , \REGISTERS[3][9] ,
         \REGISTERS[3][8] , \REGISTERS[3][7] , \REGISTERS[3][6] ,
         \REGISTERS[3][5] , \REGISTERS[3][4] , \REGISTERS[3][3] ,
         \REGISTERS[3][2] , \REGISTERS[3][1] , \REGISTERS[3][0] ,
         \REGISTERS[4][31] , \REGISTERS[4][30] , \REGISTERS[4][29] ,
         \REGISTERS[4][28] , \REGISTERS[4][27] , \REGISTERS[4][26] ,
         \REGISTERS[4][25] , \REGISTERS[4][24] , \REGISTERS[4][23] ,
         \REGISTERS[4][22] , \REGISTERS[4][21] , \REGISTERS[4][20] ,
         \REGISTERS[4][19] , \REGISTERS[4][18] , \REGISTERS[4][17] ,
         \REGISTERS[4][16] , \REGISTERS[4][15] , \REGISTERS[4][14] ,
         \REGISTERS[4][13] , \REGISTERS[4][12] , \REGISTERS[4][11] ,
         \REGISTERS[4][10] , \REGISTERS[4][9] , \REGISTERS[4][8] ,
         \REGISTERS[4][7] , \REGISTERS[4][6] , \REGISTERS[4][5] ,
         \REGISTERS[4][4] , \REGISTERS[4][3] , \REGISTERS[4][2] ,
         \REGISTERS[4][1] , \REGISTERS[4][0] , \REGISTERS[5][31] ,
         \REGISTERS[5][30] , \REGISTERS[5][29] , \REGISTERS[5][28] ,
         \REGISTERS[5][27] , \REGISTERS[5][26] , \REGISTERS[5][25] ,
         \REGISTERS[5][24] , \REGISTERS[5][23] , \REGISTERS[5][22] ,
         \REGISTERS[5][21] , \REGISTERS[5][20] , \REGISTERS[5][19] ,
         \REGISTERS[5][18] , \REGISTERS[5][17] , \REGISTERS[5][16] ,
         \REGISTERS[5][15] , \REGISTERS[5][14] , \REGISTERS[5][13] ,
         \REGISTERS[5][12] , \REGISTERS[5][11] , \REGISTERS[5][10] ,
         \REGISTERS[5][9] , \REGISTERS[5][8] , \REGISTERS[5][7] ,
         \REGISTERS[5][6] , \REGISTERS[5][5] , \REGISTERS[5][4] ,
         \REGISTERS[5][3] , \REGISTERS[5][2] , \REGISTERS[5][1] ,
         \REGISTERS[5][0] , \REGISTERS[6][31] , \REGISTERS[6][30] ,
         \REGISTERS[6][29] , \REGISTERS[6][28] , \REGISTERS[6][27] ,
         \REGISTERS[6][26] , \REGISTERS[6][25] , \REGISTERS[6][24] ,
         \REGISTERS[6][23] , \REGISTERS[6][22] , \REGISTERS[6][21] ,
         \REGISTERS[6][20] , \REGISTERS[6][19] , \REGISTERS[6][18] ,
         \REGISTERS[6][17] , \REGISTERS[6][16] , \REGISTERS[6][15] ,
         \REGISTERS[6][14] , \REGISTERS[6][13] , \REGISTERS[6][12] ,
         \REGISTERS[6][11] , \REGISTERS[6][10] , \REGISTERS[6][9] ,
         \REGISTERS[6][8] , \REGISTERS[6][7] , \REGISTERS[6][6] ,
         \REGISTERS[6][5] , \REGISTERS[6][4] , \REGISTERS[6][3] ,
         \REGISTERS[6][2] , \REGISTERS[6][1] , \REGISTERS[6][0] ,
         \REGISTERS[7][31] , \REGISTERS[7][30] , \REGISTERS[7][29] ,
         \REGISTERS[7][28] , \REGISTERS[7][27] , \REGISTERS[7][26] ,
         \REGISTERS[7][25] , \REGISTERS[7][24] , \REGISTERS[7][23] ,
         \REGISTERS[7][22] , \REGISTERS[7][21] , \REGISTERS[7][20] ,
         \REGISTERS[7][19] , \REGISTERS[7][18] , \REGISTERS[7][17] ,
         \REGISTERS[7][16] , \REGISTERS[7][15] , \REGISTERS[7][14] ,
         \REGISTERS[7][13] , \REGISTERS[7][12] , \REGISTERS[7][11] ,
         \REGISTERS[7][10] , \REGISTERS[7][9] , \REGISTERS[7][8] ,
         \REGISTERS[7][7] , \REGISTERS[7][6] , \REGISTERS[7][5] ,
         \REGISTERS[7][4] , \REGISTERS[7][3] , \REGISTERS[7][2] ,
         \REGISTERS[7][1] , \REGISTERS[7][0] , \REGISTERS[8][31] ,
         \REGISTERS[8][30] , \REGISTERS[8][29] , \REGISTERS[8][28] ,
         \REGISTERS[8][27] , \REGISTERS[8][26] , \REGISTERS[8][25] ,
         \REGISTERS[8][24] , \REGISTERS[8][23] , \REGISTERS[8][22] ,
         \REGISTERS[8][21] , \REGISTERS[8][20] , \REGISTERS[8][19] ,
         \REGISTERS[8][18] , \REGISTERS[8][17] , \REGISTERS[8][16] ,
         \REGISTERS[8][15] , \REGISTERS[8][14] , \REGISTERS[8][13] ,
         \REGISTERS[8][12] , \REGISTERS[8][11] , \REGISTERS[8][10] ,
         \REGISTERS[8][9] , \REGISTERS[8][8] , \REGISTERS[8][7] ,
         \REGISTERS[8][6] , \REGISTERS[8][5] , \REGISTERS[8][4] ,
         \REGISTERS[8][3] , \REGISTERS[8][2] , \REGISTERS[8][1] ,
         \REGISTERS[8][0] , \REGISTERS[9][31] , \REGISTERS[9][30] ,
         \REGISTERS[9][29] , \REGISTERS[9][28] , \REGISTERS[9][27] ,
         \REGISTERS[9][26] , \REGISTERS[9][25] , \REGISTERS[9][24] ,
         \REGISTERS[9][23] , \REGISTERS[9][22] , \REGISTERS[9][21] ,
         \REGISTERS[9][20] , \REGISTERS[9][19] , \REGISTERS[9][18] ,
         \REGISTERS[9][17] , \REGISTERS[9][16] , \REGISTERS[9][15] ,
         \REGISTERS[9][14] , \REGISTERS[9][13] , \REGISTERS[9][12] ,
         \REGISTERS[9][11] , \REGISTERS[9][10] , \REGISTERS[9][9] ,
         \REGISTERS[9][8] , \REGISTERS[9][7] , \REGISTERS[9][6] ,
         \REGISTERS[9][5] , \REGISTERS[9][4] , \REGISTERS[9][3] ,
         \REGISTERS[9][2] , \REGISTERS[9][1] , \REGISTERS[9][0] ,
         \REGISTERS[10][31] , \REGISTERS[10][30] , \REGISTERS[10][29] ,
         \REGISTERS[10][28] , \REGISTERS[10][27] , \REGISTERS[10][26] ,
         \REGISTERS[10][25] , \REGISTERS[10][24] , \REGISTERS[10][23] ,
         \REGISTERS[10][22] , \REGISTERS[10][21] , \REGISTERS[10][20] ,
         \REGISTERS[10][19] , \REGISTERS[10][18] , \REGISTERS[10][17] ,
         \REGISTERS[10][16] , \REGISTERS[10][15] , \REGISTERS[10][14] ,
         \REGISTERS[10][13] , \REGISTERS[10][12] , \REGISTERS[10][11] ,
         \REGISTERS[10][10] , \REGISTERS[10][9] , \REGISTERS[10][8] ,
         \REGISTERS[10][7] , \REGISTERS[10][6] , \REGISTERS[10][5] ,
         \REGISTERS[10][4] , \REGISTERS[10][3] , \REGISTERS[10][2] ,
         \REGISTERS[10][1] , \REGISTERS[10][0] , \REGISTERS[11][31] ,
         \REGISTERS[11][30] , \REGISTERS[11][29] , \REGISTERS[11][28] ,
         \REGISTERS[11][27] , \REGISTERS[11][26] , \REGISTERS[11][25] ,
         \REGISTERS[11][24] , \REGISTERS[11][23] , \REGISTERS[11][22] ,
         \REGISTERS[11][21] , \REGISTERS[11][20] , \REGISTERS[11][19] ,
         \REGISTERS[11][18] , \REGISTERS[11][17] , \REGISTERS[11][16] ,
         \REGISTERS[11][15] , \REGISTERS[11][14] , \REGISTERS[11][13] ,
         \REGISTERS[11][12] , \REGISTERS[11][11] , \REGISTERS[11][10] ,
         \REGISTERS[11][9] , \REGISTERS[11][8] , \REGISTERS[11][7] ,
         \REGISTERS[11][6] , \REGISTERS[11][5] , \REGISTERS[11][4] ,
         \REGISTERS[11][3] , \REGISTERS[11][2] , \REGISTERS[11][1] ,
         \REGISTERS[11][0] , \REGISTERS[12][31] , \REGISTERS[12][30] ,
         \REGISTERS[12][29] , \REGISTERS[12][28] , \REGISTERS[12][27] ,
         \REGISTERS[12][26] , \REGISTERS[12][25] , \REGISTERS[12][24] ,
         \REGISTERS[12][23] , \REGISTERS[12][22] , \REGISTERS[12][21] ,
         \REGISTERS[12][20] , \REGISTERS[12][19] , \REGISTERS[12][18] ,
         \REGISTERS[12][17] , \REGISTERS[12][16] , \REGISTERS[12][15] ,
         \REGISTERS[12][14] , \REGISTERS[12][13] , \REGISTERS[12][12] ,
         \REGISTERS[12][11] , \REGISTERS[12][10] , \REGISTERS[12][9] ,
         \REGISTERS[12][8] , \REGISTERS[12][7] , \REGISTERS[12][6] ,
         \REGISTERS[12][5] , \REGISTERS[12][4] , \REGISTERS[12][3] ,
         \REGISTERS[12][2] , \REGISTERS[12][1] , \REGISTERS[12][0] ,
         \REGISTERS[13][31] , \REGISTERS[13][30] , \REGISTERS[13][29] ,
         \REGISTERS[13][28] , \REGISTERS[13][27] , \REGISTERS[13][26] ,
         \REGISTERS[13][25] , \REGISTERS[13][24] , \REGISTERS[13][23] ,
         \REGISTERS[13][22] , \REGISTERS[13][21] , \REGISTERS[13][20] ,
         \REGISTERS[13][19] , \REGISTERS[13][18] , \REGISTERS[13][17] ,
         \REGISTERS[13][16] , \REGISTERS[13][15] , \REGISTERS[13][14] ,
         \REGISTERS[13][13] , \REGISTERS[13][12] , \REGISTERS[13][11] ,
         \REGISTERS[13][10] , \REGISTERS[13][9] , \REGISTERS[13][8] ,
         \REGISTERS[13][7] , \REGISTERS[13][6] , \REGISTERS[13][5] ,
         \REGISTERS[13][4] , \REGISTERS[13][3] , \REGISTERS[13][2] ,
         \REGISTERS[13][1] , \REGISTERS[13][0] , \REGISTERS[14][31] ,
         \REGISTERS[14][30] , \REGISTERS[14][29] , \REGISTERS[14][28] ,
         \REGISTERS[14][27] , \REGISTERS[14][26] , \REGISTERS[14][25] ,
         \REGISTERS[14][24] , \REGISTERS[14][23] , \REGISTERS[14][22] ,
         \REGISTERS[14][21] , \REGISTERS[14][20] , \REGISTERS[14][19] ,
         \REGISTERS[14][18] , \REGISTERS[14][17] , \REGISTERS[14][16] ,
         \REGISTERS[14][15] , \REGISTERS[14][14] , \REGISTERS[14][13] ,
         \REGISTERS[14][12] , \REGISTERS[14][11] , \REGISTERS[14][10] ,
         \REGISTERS[14][9] , \REGISTERS[14][8] , \REGISTERS[14][7] ,
         \REGISTERS[14][6] , \REGISTERS[14][5] , \REGISTERS[14][4] ,
         \REGISTERS[14][3] , \REGISTERS[14][2] , \REGISTERS[14][1] ,
         \REGISTERS[14][0] , \REGISTERS[15][31] , \REGISTERS[15][30] ,
         \REGISTERS[15][29] , \REGISTERS[15][28] , \REGISTERS[15][27] ,
         \REGISTERS[15][26] , \REGISTERS[15][25] , \REGISTERS[15][24] ,
         \REGISTERS[15][23] , \REGISTERS[15][22] , \REGISTERS[15][21] ,
         \REGISTERS[15][20] , \REGISTERS[15][19] , \REGISTERS[15][18] ,
         \REGISTERS[15][17] , \REGISTERS[15][16] , \REGISTERS[15][15] ,
         \REGISTERS[15][14] , \REGISTERS[15][13] , \REGISTERS[15][12] ,
         \REGISTERS[15][11] , \REGISTERS[15][10] , \REGISTERS[15][9] ,
         \REGISTERS[15][8] , \REGISTERS[15][7] , \REGISTERS[15][6] ,
         \REGISTERS[15][5] , \REGISTERS[15][4] , \REGISTERS[15][3] ,
         \REGISTERS[15][2] , \REGISTERS[15][1] , \REGISTERS[15][0] ,
         \REGISTERS[16][31] , \REGISTERS[16][30] , \REGISTERS[16][29] ,
         \REGISTERS[16][28] , \REGISTERS[16][27] , \REGISTERS[16][26] ,
         \REGISTERS[16][25] , \REGISTERS[16][24] , \REGISTERS[16][23] ,
         \REGISTERS[16][22] , \REGISTERS[16][21] , \REGISTERS[16][20] ,
         \REGISTERS[16][19] , \REGISTERS[16][18] , \REGISTERS[16][17] ,
         \REGISTERS[16][16] , \REGISTERS[16][15] , \REGISTERS[16][14] ,
         \REGISTERS[16][13] , \REGISTERS[16][12] , \REGISTERS[16][11] ,
         \REGISTERS[16][10] , \REGISTERS[16][9] , \REGISTERS[16][8] ,
         \REGISTERS[16][7] , \REGISTERS[16][6] , \REGISTERS[16][5] ,
         \REGISTERS[16][4] , \REGISTERS[16][3] , \REGISTERS[16][2] ,
         \REGISTERS[16][1] , \REGISTERS[16][0] , \REGISTERS[17][31] ,
         \REGISTERS[17][30] , \REGISTERS[17][29] , \REGISTERS[17][28] ,
         \REGISTERS[17][27] , \REGISTERS[17][26] , \REGISTERS[17][25] ,
         \REGISTERS[17][24] , \REGISTERS[17][23] , \REGISTERS[17][22] ,
         \REGISTERS[17][21] , \REGISTERS[17][20] , \REGISTERS[17][19] ,
         \REGISTERS[17][18] , \REGISTERS[17][17] , \REGISTERS[17][16] ,
         \REGISTERS[17][15] , \REGISTERS[17][14] , \REGISTERS[17][13] ,
         \REGISTERS[17][12] , \REGISTERS[17][11] , \REGISTERS[17][10] ,
         \REGISTERS[17][9] , \REGISTERS[17][8] , \REGISTERS[17][7] ,
         \REGISTERS[17][6] , \REGISTERS[17][5] , \REGISTERS[17][4] ,
         \REGISTERS[17][3] , \REGISTERS[17][2] , \REGISTERS[17][1] ,
         \REGISTERS[17][0] , \REGISTERS[18][31] , \REGISTERS[18][30] ,
         \REGISTERS[18][29] , \REGISTERS[18][28] , \REGISTERS[18][27] ,
         \REGISTERS[18][26] , \REGISTERS[18][25] , \REGISTERS[18][24] ,
         \REGISTERS[18][23] , \REGISTERS[18][22] , \REGISTERS[18][21] ,
         \REGISTERS[18][20] , \REGISTERS[18][19] , \REGISTERS[18][18] ,
         \REGISTERS[18][17] , \REGISTERS[18][16] , \REGISTERS[18][15] ,
         \REGISTERS[18][14] , \REGISTERS[18][13] , \REGISTERS[18][12] ,
         \REGISTERS[18][11] , \REGISTERS[18][10] , \REGISTERS[18][9] ,
         \REGISTERS[18][8] , \REGISTERS[18][7] , \REGISTERS[18][6] ,
         \REGISTERS[18][5] , \REGISTERS[18][4] , \REGISTERS[18][3] ,
         \REGISTERS[18][2] , \REGISTERS[18][1] , \REGISTERS[18][0] ,
         \REGISTERS[19][31] , \REGISTERS[19][30] , \REGISTERS[19][29] ,
         \REGISTERS[19][28] , \REGISTERS[19][27] , \REGISTERS[19][26] ,
         \REGISTERS[19][25] , \REGISTERS[19][24] , \REGISTERS[19][23] ,
         \REGISTERS[19][22] , \REGISTERS[19][21] , \REGISTERS[19][20] ,
         \REGISTERS[19][19] , \REGISTERS[19][18] , \REGISTERS[19][17] ,
         \REGISTERS[19][16] , \REGISTERS[19][15] , \REGISTERS[19][14] ,
         \REGISTERS[19][13] , \REGISTERS[19][12] , \REGISTERS[19][11] ,
         \REGISTERS[19][10] , \REGISTERS[19][9] , \REGISTERS[19][8] ,
         \REGISTERS[19][7] , \REGISTERS[19][6] , \REGISTERS[19][5] ,
         \REGISTERS[19][4] , \REGISTERS[19][3] , \REGISTERS[19][2] ,
         \REGISTERS[19][1] , \REGISTERS[19][0] , \REGISTERS[20][31] ,
         \REGISTERS[20][30] , \REGISTERS[20][29] , \REGISTERS[20][28] ,
         \REGISTERS[20][27] , \REGISTERS[20][26] , \REGISTERS[20][25] ,
         \REGISTERS[20][24] , \REGISTERS[20][23] , \REGISTERS[20][22] ,
         \REGISTERS[20][21] , \REGISTERS[20][20] , \REGISTERS[20][19] ,
         \REGISTERS[20][18] , \REGISTERS[20][17] , \REGISTERS[20][16] ,
         \REGISTERS[20][15] , \REGISTERS[20][14] , \REGISTERS[20][13] ,
         \REGISTERS[20][12] , \REGISTERS[20][11] , \REGISTERS[20][10] ,
         \REGISTERS[20][9] , \REGISTERS[20][8] , \REGISTERS[20][7] ,
         \REGISTERS[20][6] , \REGISTERS[20][5] , \REGISTERS[20][4] ,
         \REGISTERS[20][3] , \REGISTERS[20][2] , \REGISTERS[20][1] ,
         \REGISTERS[20][0] , \REGISTERS[21][31] , \REGISTERS[21][30] ,
         \REGISTERS[21][29] , \REGISTERS[21][28] , \REGISTERS[21][27] ,
         \REGISTERS[21][26] , \REGISTERS[21][25] , \REGISTERS[21][24] ,
         \REGISTERS[21][23] , \REGISTERS[21][22] , \REGISTERS[21][21] ,
         \REGISTERS[21][20] , \REGISTERS[21][19] , \REGISTERS[21][18] ,
         \REGISTERS[21][17] , \REGISTERS[21][16] , \REGISTERS[21][15] ,
         \REGISTERS[21][14] , \REGISTERS[21][13] , \REGISTERS[21][12] ,
         \REGISTERS[21][11] , \REGISTERS[21][10] , \REGISTERS[21][9] ,
         \REGISTERS[21][8] , \REGISTERS[21][7] , \REGISTERS[21][6] ,
         \REGISTERS[21][5] , \REGISTERS[21][4] , \REGISTERS[21][3] ,
         \REGISTERS[21][2] , \REGISTERS[21][1] , \REGISTERS[21][0] ,
         \REGISTERS[22][31] , \REGISTERS[22][30] , \REGISTERS[22][29] ,
         \REGISTERS[22][28] , \REGISTERS[22][27] , \REGISTERS[22][26] ,
         \REGISTERS[22][25] , \REGISTERS[22][24] , \REGISTERS[22][23] ,
         \REGISTERS[22][22] , \REGISTERS[22][21] , \REGISTERS[22][20] ,
         \REGISTERS[22][19] , \REGISTERS[22][18] , \REGISTERS[22][17] ,
         \REGISTERS[22][16] , \REGISTERS[22][15] , \REGISTERS[22][14] ,
         \REGISTERS[22][13] , \REGISTERS[22][12] , \REGISTERS[22][11] ,
         \REGISTERS[22][10] , \REGISTERS[22][9] , \REGISTERS[22][8] ,
         \REGISTERS[22][7] , \REGISTERS[22][6] , \REGISTERS[22][5] ,
         \REGISTERS[22][4] , \REGISTERS[22][3] , \REGISTERS[22][2] ,
         \REGISTERS[22][1] , \REGISTERS[22][0] , \REGISTERS[23][31] ,
         \REGISTERS[23][30] , \REGISTERS[23][29] , \REGISTERS[23][28] ,
         \REGISTERS[23][27] , \REGISTERS[23][26] , \REGISTERS[23][25] ,
         \REGISTERS[23][24] , \REGISTERS[23][23] , \REGISTERS[23][22] ,
         \REGISTERS[23][21] , \REGISTERS[23][20] , \REGISTERS[23][19] ,
         \REGISTERS[23][18] , \REGISTERS[23][17] , \REGISTERS[23][16] ,
         \REGISTERS[23][15] , \REGISTERS[23][14] , \REGISTERS[23][13] ,
         \REGISTERS[23][12] , \REGISTERS[23][11] , \REGISTERS[23][10] ,
         \REGISTERS[23][9] , \REGISTERS[23][8] , \REGISTERS[23][7] ,
         \REGISTERS[23][6] , \REGISTERS[23][5] , \REGISTERS[23][4] ,
         \REGISTERS[23][3] , \REGISTERS[23][2] , \REGISTERS[23][1] ,
         \REGISTERS[23][0] , \REGISTERS[24][31] , \REGISTERS[24][30] ,
         \REGISTERS[24][29] , \REGISTERS[24][28] , \REGISTERS[24][27] ,
         \REGISTERS[24][26] , \REGISTERS[24][25] , \REGISTERS[24][24] ,
         \REGISTERS[24][23] , \REGISTERS[24][22] , \REGISTERS[24][21] ,
         \REGISTERS[24][20] , \REGISTERS[24][19] , \REGISTERS[24][18] ,
         \REGISTERS[24][17] , \REGISTERS[24][16] , \REGISTERS[24][15] ,
         \REGISTERS[24][14] , \REGISTERS[24][13] , \REGISTERS[24][12] ,
         \REGISTERS[24][11] , \REGISTERS[24][10] , \REGISTERS[24][9] ,
         \REGISTERS[24][8] , \REGISTERS[24][7] , \REGISTERS[24][6] ,
         \REGISTERS[24][5] , \REGISTERS[24][4] , \REGISTERS[24][3] ,
         \REGISTERS[24][2] , \REGISTERS[24][1] , \REGISTERS[24][0] ,
         \REGISTERS[25][31] , \REGISTERS[25][30] , \REGISTERS[25][29] ,
         \REGISTERS[25][28] , \REGISTERS[25][27] , \REGISTERS[25][26] ,
         \REGISTERS[25][25] , \REGISTERS[25][24] , \REGISTERS[25][23] ,
         \REGISTERS[25][22] , \REGISTERS[25][21] , \REGISTERS[25][20] ,
         \REGISTERS[25][19] , \REGISTERS[25][18] , \REGISTERS[25][17] ,
         \REGISTERS[25][16] , \REGISTERS[25][15] , \REGISTERS[25][14] ,
         \REGISTERS[25][13] , \REGISTERS[25][12] , \REGISTERS[25][11] ,
         \REGISTERS[25][10] , \REGISTERS[25][9] , \REGISTERS[25][8] ,
         \REGISTERS[25][7] , \REGISTERS[25][6] , \REGISTERS[25][5] ,
         \REGISTERS[25][4] , \REGISTERS[25][3] , \REGISTERS[25][2] ,
         \REGISTERS[25][1] , \REGISTERS[25][0] , \REGISTERS[26][31] ,
         \REGISTERS[26][30] , \REGISTERS[26][29] , \REGISTERS[26][28] ,
         \REGISTERS[26][27] , \REGISTERS[26][26] , \REGISTERS[26][25] ,
         \REGISTERS[26][24] , \REGISTERS[26][23] , \REGISTERS[26][22] ,
         \REGISTERS[26][21] , \REGISTERS[26][20] , \REGISTERS[26][19] ,
         \REGISTERS[26][18] , \REGISTERS[26][17] , \REGISTERS[26][16] ,
         \REGISTERS[26][15] , \REGISTERS[26][14] , \REGISTERS[26][13] ,
         \REGISTERS[26][12] , \REGISTERS[26][11] , \REGISTERS[26][10] ,
         \REGISTERS[26][9] , \REGISTERS[26][8] , \REGISTERS[26][7] ,
         \REGISTERS[26][6] , \REGISTERS[26][5] , \REGISTERS[26][4] ,
         \REGISTERS[26][3] , \REGISTERS[26][2] , \REGISTERS[26][1] ,
         \REGISTERS[26][0] , \REGISTERS[27][31] , \REGISTERS[27][30] ,
         \REGISTERS[27][29] , \REGISTERS[27][28] , \REGISTERS[27][27] ,
         \REGISTERS[27][26] , \REGISTERS[27][25] , \REGISTERS[27][24] ,
         \REGISTERS[27][23] , \REGISTERS[27][22] , \REGISTERS[27][21] ,
         \REGISTERS[27][20] , \REGISTERS[27][19] , \REGISTERS[27][18] ,
         \REGISTERS[27][17] , \REGISTERS[27][16] , \REGISTERS[27][15] ,
         \REGISTERS[27][14] , \REGISTERS[27][13] , \REGISTERS[27][12] ,
         \REGISTERS[27][11] , \REGISTERS[27][10] , \REGISTERS[27][9] ,
         \REGISTERS[27][8] , \REGISTERS[27][7] , \REGISTERS[27][6] ,
         \REGISTERS[27][5] , \REGISTERS[27][4] , \REGISTERS[27][3] ,
         \REGISTERS[27][2] , \REGISTERS[27][1] , \REGISTERS[27][0] ,
         \REGISTERS[28][31] , \REGISTERS[28][30] , \REGISTERS[28][29] ,
         \REGISTERS[28][28] , \REGISTERS[28][27] , \REGISTERS[28][26] ,
         \REGISTERS[28][25] , \REGISTERS[28][24] , \REGISTERS[28][23] ,
         \REGISTERS[28][22] , \REGISTERS[28][21] , \REGISTERS[28][20] ,
         \REGISTERS[28][19] , \REGISTERS[28][18] , \REGISTERS[28][17] ,
         \REGISTERS[28][16] , \REGISTERS[28][15] , \REGISTERS[28][14] ,
         \REGISTERS[28][13] , \REGISTERS[28][12] , \REGISTERS[28][11] ,
         \REGISTERS[28][10] , \REGISTERS[28][9] , \REGISTERS[28][8] ,
         \REGISTERS[28][7] , \REGISTERS[28][6] , \REGISTERS[28][5] ,
         \REGISTERS[28][4] , \REGISTERS[28][3] , \REGISTERS[28][2] ,
         \REGISTERS[28][1] , \REGISTERS[28][0] , \REGISTERS[29][31] ,
         \REGISTERS[29][30] , \REGISTERS[29][29] , \REGISTERS[29][28] ,
         \REGISTERS[29][27] , \REGISTERS[29][26] , \REGISTERS[29][25] ,
         \REGISTERS[29][24] , \REGISTERS[29][23] , \REGISTERS[29][22] ,
         \REGISTERS[29][21] , \REGISTERS[29][20] , \REGISTERS[29][19] ,
         \REGISTERS[29][18] , \REGISTERS[29][17] , \REGISTERS[29][16] ,
         \REGISTERS[29][15] , \REGISTERS[29][14] , \REGISTERS[29][13] ,
         \REGISTERS[29][12] , \REGISTERS[29][11] , \REGISTERS[29][10] ,
         \REGISTERS[29][9] , \REGISTERS[29][8] , \REGISTERS[29][7] ,
         \REGISTERS[29][6] , \REGISTERS[29][5] , \REGISTERS[29][4] ,
         \REGISTERS[29][3] , \REGISTERS[29][2] , \REGISTERS[29][1] ,
         \REGISTERS[29][0] , \REGISTERS[30][31] , \REGISTERS[30][30] ,
         \REGISTERS[30][29] , \REGISTERS[30][28] , \REGISTERS[30][27] ,
         \REGISTERS[30][26] , \REGISTERS[30][25] , \REGISTERS[30][24] ,
         \REGISTERS[30][23] , \REGISTERS[30][22] , \REGISTERS[30][21] ,
         \REGISTERS[30][20] , \REGISTERS[30][19] , \REGISTERS[30][18] ,
         \REGISTERS[30][17] , \REGISTERS[30][16] , \REGISTERS[30][15] ,
         \REGISTERS[30][14] , \REGISTERS[30][13] , \REGISTERS[30][12] ,
         \REGISTERS[30][11] , \REGISTERS[30][10] , \REGISTERS[30][9] ,
         \REGISTERS[30][8] , \REGISTERS[30][7] , \REGISTERS[30][6] ,
         \REGISTERS[30][5] , \REGISTERS[30][4] , \REGISTERS[30][3] ,
         \REGISTERS[30][2] , \REGISTERS[30][1] , \REGISTERS[30][0] ,
         \REGISTERS[31][31] , \REGISTERS[31][30] , \REGISTERS[31][29] ,
         \REGISTERS[31][28] , \REGISTERS[31][27] , \REGISTERS[31][26] ,
         \REGISTERS[31][25] , \REGISTERS[31][24] , \REGISTERS[31][23] ,
         \REGISTERS[31][22] , \REGISTERS[31][21] , \REGISTERS[31][20] ,
         \REGISTERS[31][19] , \REGISTERS[31][18] , \REGISTERS[31][17] ,
         \REGISTERS[31][16] , \REGISTERS[31][15] , \REGISTERS[31][14] ,
         \REGISTERS[31][13] , \REGISTERS[31][12] , \REGISTERS[31][11] ,
         \REGISTERS[31][10] , \REGISTERS[31][9] , \REGISTERS[31][8] ,
         \REGISTERS[31][7] , \REGISTERS[31][6] , \REGISTERS[31][5] ,
         \REGISTERS[31][4] , \REGISTERS[31][3] , \REGISTERS[31][2] ,
         \REGISTERS[31][1] , \REGISTERS[31][0] , N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858;

  DLH_X1 \REGISTERS_reg[1][31]  ( .G(N305), .D(N275), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(N305), .D(N274), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(N305), .D(N273), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(n36299), .D(N272), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(N305), .D(N271), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(N305), .D(N270), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(N305), .D(N269), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(N305), .D(N268), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(N305), .D(N267), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(N305), .D(N266), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(n36299), .D(N265), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n36299), .D(N264), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n36299), .D(N263), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(n36299), .D(N262), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(n36299), .D(N261), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(N305), .D(N260), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(N305), .D(N259), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(n36299), .D(N258), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(N305), .D(N257), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(N305), .D(N256), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n36299), .D(N255), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(n36299), .D(N254), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(n36299), .D(N253), .Q(\REGISTERS[1][9] )
         );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(n36299), .D(N252), .Q(\REGISTERS[1][8] )
         );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n36299), .D(N251), .Q(\REGISTERS[1][7] )
         );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(N305), .D(N250), .Q(\REGISTERS[1][6] ) );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n36299), .D(N249), .Q(\REGISTERS[1][5] )
         );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(n36299), .D(N248), .Q(\REGISTERS[1][4] )
         );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(n36299), .D(N247), .Q(\REGISTERS[1][3] )
         );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(n36299), .D(N246), .Q(\REGISTERS[1][2] )
         );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(N305), .D(N245), .Q(\REGISTERS[1][1] ) );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n36299), .D(N244), .Q(\REGISTERS[1][0] )
         );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(N304), .D(N275), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(N304), .D(N274), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(N304), .D(N273), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(N304), .D(N272), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(N304), .D(N271), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(N304), .D(N270), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(n36300), .D(N269), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(n36300), .D(N268), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n36300), .D(N267), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n36300), .D(N266), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(N304), .D(N265), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(N304), .D(N264), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n36300), .D(N263), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(n36300), .D(N262), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n36300), .D(N261), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(N304), .D(N260), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(N304), .D(N259), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(N304), .D(N258), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(N304), .D(N257), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(N304), .D(N256), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(n36300), .D(N255), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n36300), .D(N254), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(n36300), .D(N253), .Q(\REGISTERS[2][9] )
         );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(n36300), .D(N252), .Q(\REGISTERS[2][8] )
         );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n36300), .D(N251), .Q(\REGISTERS[2][7] )
         );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(N304), .D(N250), .Q(\REGISTERS[2][6] ) );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(n36300), .D(N249), .Q(\REGISTERS[2][5] )
         );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(n36300), .D(N248), .Q(\REGISTERS[2][4] )
         );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(n36300), .D(N247), .Q(\REGISTERS[2][3] )
         );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(n36300), .D(N246), .Q(\REGISTERS[2][2] )
         );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(N304), .D(N245), .Q(\REGISTERS[2][1] ) );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(n36300), .D(N244), .Q(\REGISTERS[2][0] )
         );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(N303), .D(N275), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(N303), .D(N274), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(N303), .D(N273), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(N303), .D(N272), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(N303), .D(N271), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(N303), .D(N270), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(n36301), .D(N269), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(n36301), .D(N268), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n36301), .D(N267), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n36301), .D(N266), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(N303), .D(N265), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(N303), .D(N264), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n36301), .D(N263), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(n36301), .D(N262), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n36301), .D(N261), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(N303), .D(N260), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(N303), .D(N259), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(N303), .D(N258), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(N303), .D(N257), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(N303), .D(N256), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(n36301), .D(N255), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n36301), .D(N254), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(n36301), .D(N253), .Q(\REGISTERS[3][9] )
         );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(n36301), .D(N252), .Q(\REGISTERS[3][8] )
         );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n36301), .D(N251), .Q(\REGISTERS[3][7] )
         );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(N303), .D(N250), .Q(\REGISTERS[3][6] ) );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(n36301), .D(N249), .Q(\REGISTERS[3][5] )
         );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(n36301), .D(N248), .Q(\REGISTERS[3][4] )
         );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(n36301), .D(N247), .Q(\REGISTERS[3][3] )
         );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(n36301), .D(N246), .Q(\REGISTERS[3][2] )
         );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(N303), .D(N245), .Q(\REGISTERS[3][1] ) );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(n36301), .D(N244), .Q(\REGISTERS[3][0] )
         );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(N302), .D(N275), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(N302), .D(N274), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(N302), .D(N273), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(N302), .D(N272), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(N302), .D(N271), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(N302), .D(N270), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(n36302), .D(N269), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(n36302), .D(N268), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n36302), .D(N267), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n36302), .D(N266), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(N302), .D(N265), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(N302), .D(N264), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n36302), .D(N263), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(n36302), .D(N262), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n36302), .D(N261), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(N302), .D(N260), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(N302), .D(N259), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(N302), .D(N258), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(N302), .D(N257), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(N302), .D(N256), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(n36302), .D(N255), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n36302), .D(N254), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(n36302), .D(N253), .Q(\REGISTERS[4][9] )
         );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(n36302), .D(N252), .Q(\REGISTERS[4][8] )
         );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(n36302), .D(N251), .Q(\REGISTERS[4][7] )
         );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(N302), .D(N250), .Q(\REGISTERS[4][6] ) );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(n36302), .D(N249), .Q(\REGISTERS[4][5] )
         );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(n36302), .D(N248), .Q(\REGISTERS[4][4] )
         );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(n36302), .D(N247), .Q(\REGISTERS[4][3] )
         );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(n36302), .D(N246), .Q(\REGISTERS[4][2] )
         );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(N302), .D(N245), .Q(\REGISTERS[4][1] ) );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n36302), .D(N244), .Q(\REGISTERS[4][0] )
         );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(N301), .D(N275), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(N301), .D(N274), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(N301), .D(N273), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(N301), .D(N272), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(N301), .D(N271), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(N301), .D(N270), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(n36303), .D(N269), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(n36303), .D(N268), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n36303), .D(N267), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n36303), .D(N266), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(N301), .D(N265), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(N301), .D(N264), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n36303), .D(N263), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(n36303), .D(N262), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n36303), .D(N261), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(N301), .D(N260), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(N301), .D(N259), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(N301), .D(N258), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(N301), .D(N257), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(N301), .D(N256), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(n36303), .D(N255), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n36303), .D(N254), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(n36303), .D(N253), .Q(\REGISTERS[5][9] )
         );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(n36303), .D(N252), .Q(\REGISTERS[5][8] )
         );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n36303), .D(N251), .Q(\REGISTERS[5][7] )
         );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(N301), .D(N250), .Q(\REGISTERS[5][6] ) );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(n36303), .D(N249), .Q(\REGISTERS[5][5] )
         );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(n36303), .D(N248), .Q(\REGISTERS[5][4] )
         );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(n36303), .D(N247), .Q(\REGISTERS[5][3] )
         );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(n36303), .D(N246), .Q(\REGISTERS[5][2] )
         );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(N301), .D(N245), .Q(\REGISTERS[5][1] ) );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(n36303), .D(N244), .Q(\REGISTERS[5][0] )
         );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(N300), .D(N275), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(N300), .D(N274), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(N300), .D(N273), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(N300), .D(N272), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(N300), .D(N271), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(N300), .D(N270), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(n36304), .D(N269), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(n36304), .D(N268), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n36304), .D(N267), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n36304), .D(N266), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(N300), .D(N265), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(N300), .D(N264), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n36304), .D(N263), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(n36304), .D(N262), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n36304), .D(N261), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(N300), .D(N260), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(N300), .D(N259), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(N300), .D(N258), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(N300), .D(N257), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(N300), .D(N256), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(n36304), .D(N255), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n36304), .D(N254), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(n36304), .D(N253), .Q(\REGISTERS[6][9] )
         );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(n36304), .D(N252), .Q(\REGISTERS[6][8] )
         );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(n36304), .D(N251), .Q(\REGISTERS[6][7] )
         );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(N300), .D(N250), .Q(\REGISTERS[6][6] ) );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(n36304), .D(N249), .Q(\REGISTERS[6][5] )
         );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(n36304), .D(N248), .Q(\REGISTERS[6][4] )
         );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(n36304), .D(N247), .Q(\REGISTERS[6][3] )
         );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(n36304), .D(N246), .Q(\REGISTERS[6][2] )
         );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(N300), .D(N245), .Q(\REGISTERS[6][1] ) );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n36304), .D(N244), .Q(\REGISTERS[6][0] )
         );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(N299), .D(N275), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(N299), .D(N274), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(N299), .D(N273), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(N299), .D(N272), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(N299), .D(N271), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(N299), .D(N270), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(n36305), .D(N269), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(n36305), .D(N268), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n36305), .D(N267), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n36305), .D(N266), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(N299), .D(N265), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(N299), .D(N264), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n36305), .D(N263), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(n36305), .D(N262), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n36305), .D(N261), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(N299), .D(N260), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(N299), .D(N259), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(N299), .D(N258), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(N299), .D(N257), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(N299), .D(N256), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(n36305), .D(N255), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n36305), .D(N254), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(n36305), .D(N253), .Q(\REGISTERS[7][9] )
         );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(n36305), .D(N252), .Q(\REGISTERS[7][8] )
         );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n36305), .D(N251), .Q(\REGISTERS[7][7] )
         );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(N299), .D(N250), .Q(\REGISTERS[7][6] ) );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(n36305), .D(N249), .Q(\REGISTERS[7][5] )
         );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(n36305), .D(N248), .Q(\REGISTERS[7][4] )
         );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(n36305), .D(N247), .Q(\REGISTERS[7][3] )
         );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(n36305), .D(N246), .Q(\REGISTERS[7][2] )
         );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(N299), .D(N245), .Q(\REGISTERS[7][1] ) );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(n36305), .D(N244), .Q(\REGISTERS[7][0] )
         );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(N298), .D(N275), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(N298), .D(N274), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(N298), .D(N273), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(N298), .D(N272), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(N298), .D(N271), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(N298), .D(N270), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(n36306), .D(N269), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(n36306), .D(N268), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n36306), .D(N267), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n36306), .D(N266), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(N298), .D(N265), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(N298), .D(N264), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n36306), .D(N263), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(n36306), .D(N262), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n36306), .D(N261), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(n36306), .D(N260), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(N298), .D(N259), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(N298), .D(N258), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(N298), .D(N257), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(N298), .D(N256), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(n36306), .D(N255), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n36306), .D(N254), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(n36306), .D(N253), .Q(\REGISTERS[8][9] )
         );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(n36306), .D(N252), .Q(\REGISTERS[8][8] )
         );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n36306), .D(N251), .Q(\REGISTERS[8][7] )
         );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(N298), .D(N250), .Q(\REGISTERS[8][6] ) );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(n36306), .D(N249), .Q(\REGISTERS[8][5] )
         );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(n36306), .D(N248), .Q(\REGISTERS[8][4] )
         );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(n36306), .D(N247), .Q(\REGISTERS[8][3] )
         );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(n36306), .D(N246), .Q(\REGISTERS[8][2] )
         );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(N298), .D(N245), .Q(\REGISTERS[8][1] ) );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(N298), .D(N244), .Q(\REGISTERS[8][0] ) );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(N297), .D(N275), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(N297), .D(N274), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(N297), .D(N273), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(N297), .D(N272), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(N297), .D(N271), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(N297), .D(N270), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(n36307), .D(N269), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(n36307), .D(N268), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n36307), .D(N267), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n36307), .D(N266), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(N297), .D(N265), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(N297), .D(N264), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n36307), .D(N263), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(n36307), .D(N262), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n36307), .D(N261), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(N297), .D(N260), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(N297), .D(N259), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(N297), .D(N258), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(N297), .D(N257), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(N297), .D(N256), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(n36307), .D(N255), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n36307), .D(N254), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(n36307), .D(N253), .Q(\REGISTERS[9][9] )
         );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(n36307), .D(N252), .Q(\REGISTERS[9][8] )
         );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n36307), .D(N251), .Q(\REGISTERS[9][7] )
         );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(N297), .D(N250), .Q(\REGISTERS[9][6] ) );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(n36307), .D(N249), .Q(\REGISTERS[9][5] )
         );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(n36307), .D(N248), .Q(\REGISTERS[9][4] )
         );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(n36307), .D(N247), .Q(\REGISTERS[9][3] )
         );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(n36307), .D(N246), .Q(\REGISTERS[9][2] )
         );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(N297), .D(N245), .Q(\REGISTERS[9][1] ) );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(n36307), .D(N244), .Q(\REGISTERS[9][0] )
         );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(N296), .D(N275), .Q(\REGISTERS[10][31] )
         );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(N296), .D(N274), .Q(\REGISTERS[10][30] )
         );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(N296), .D(N273), .Q(\REGISTERS[10][29] )
         );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(N296), .D(N272), .Q(\REGISTERS[10][28] )
         );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(N296), .D(N271), .Q(\REGISTERS[10][27] )
         );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(N296), .D(N270), .Q(\REGISTERS[10][26] )
         );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(n36308), .D(N269), .Q(
        \REGISTERS[10][25] ) );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(n36308), .D(N268), .Q(
        \REGISTERS[10][24] ) );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n36308), .D(N267), .Q(
        \REGISTERS[10][23] ) );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(n36308), .D(N266), .Q(
        \REGISTERS[10][22] ) );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(N296), .D(N265), .Q(\REGISTERS[10][21] )
         );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(N296), .D(N264), .Q(\REGISTERS[10][20] )
         );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n36308), .D(N263), .Q(
        \REGISTERS[10][19] ) );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(n36308), .D(N262), .Q(
        \REGISTERS[10][18] ) );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(N296), .D(N261), .Q(\REGISTERS[10][17] )
         );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n36308), .D(N260), .Q(
        \REGISTERS[10][16] ) );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(N296), .D(N259), .Q(\REGISTERS[10][15] )
         );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(N296), .D(N258), .Q(\REGISTERS[10][14] )
         );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n36308), .D(N257), .Q(
        \REGISTERS[10][13] ) );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(N296), .D(N256), .Q(\REGISTERS[10][12] )
         );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n36308), .D(N255), .Q(
        \REGISTERS[10][11] ) );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n36308), .D(N254), .Q(
        \REGISTERS[10][10] ) );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(n36308), .D(N253), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(n36308), .D(N252), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(n36308), .D(N251), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(N296), .D(N250), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(n36308), .D(N249), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(n36308), .D(N248), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(n36308), .D(N247), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(n36308), .D(N246), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(N296), .D(N245), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(N296), .D(N244), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(N295), .D(N275), .Q(\REGISTERS[11][31] )
         );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(N295), .D(N274), .Q(\REGISTERS[11][30] )
         );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(N295), .D(N273), .Q(\REGISTERS[11][29] )
         );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(N295), .D(N272), .Q(\REGISTERS[11][28] )
         );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(N295), .D(N271), .Q(\REGISTERS[11][27] )
         );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(N295), .D(N270), .Q(\REGISTERS[11][26] )
         );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(n36309), .D(N269), .Q(
        \REGISTERS[11][25] ) );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(n36309), .D(N268), .Q(
        \REGISTERS[11][24] ) );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n36309), .D(N267), .Q(
        \REGISTERS[11][23] ) );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n36309), .D(N266), .Q(
        \REGISTERS[11][22] ) );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(N295), .D(N265), .Q(\REGISTERS[11][21] )
         );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(N295), .D(N264), .Q(\REGISTERS[11][20] )
         );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n36309), .D(N263), .Q(
        \REGISTERS[11][19] ) );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(n36309), .D(N262), .Q(
        \REGISTERS[11][18] ) );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n36309), .D(N261), .Q(
        \REGISTERS[11][17] ) );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(N295), .D(N260), .Q(\REGISTERS[11][16] )
         );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(N295), .D(N259), .Q(\REGISTERS[11][15] )
         );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(N295), .D(N258), .Q(\REGISTERS[11][14] )
         );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(N295), .D(N257), .Q(\REGISTERS[11][13] )
         );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(N295), .D(N256), .Q(\REGISTERS[11][12] )
         );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(n36309), .D(N255), .Q(
        \REGISTERS[11][11] ) );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n36309), .D(N254), .Q(
        \REGISTERS[11][10] ) );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(n36309), .D(N253), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(n36309), .D(N252), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n36309), .D(N251), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(N295), .D(N250), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(n36309), .D(N249), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(n36309), .D(N248), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(n36309), .D(N247), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(n36309), .D(N246), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(N295), .D(N245), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(n36309), .D(N244), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(N294), .D(N275), .Q(\REGISTERS[12][31] )
         );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(N294), .D(N274), .Q(\REGISTERS[12][30] )
         );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(N294), .D(N273), .Q(\REGISTERS[12][29] )
         );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(N294), .D(N272), .Q(\REGISTERS[12][28] )
         );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(N294), .D(N271), .Q(\REGISTERS[12][27] )
         );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(N294), .D(N270), .Q(\REGISTERS[12][26] )
         );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(n36310), .D(N269), .Q(
        \REGISTERS[12][25] ) );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(n36310), .D(N268), .Q(
        \REGISTERS[12][24] ) );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n36310), .D(N267), .Q(
        \REGISTERS[12][23] ) );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n36310), .D(N266), .Q(
        \REGISTERS[12][22] ) );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(N294), .D(N265), .Q(\REGISTERS[12][21] )
         );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(N294), .D(N264), .Q(\REGISTERS[12][20] )
         );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n36310), .D(N263), .Q(
        \REGISTERS[12][19] ) );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(n36310), .D(N262), .Q(
        \REGISTERS[12][18] ) );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n36310), .D(N261), .Q(
        \REGISTERS[12][17] ) );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(N294), .D(N260), .Q(\REGISTERS[12][16] )
         );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(N294), .D(N259), .Q(\REGISTERS[12][15] )
         );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(N294), .D(N258), .Q(\REGISTERS[12][14] )
         );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(N294), .D(N257), .Q(\REGISTERS[12][13] )
         );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(N294), .D(N256), .Q(\REGISTERS[12][12] )
         );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n36310), .D(N255), .Q(
        \REGISTERS[12][11] ) );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n36310), .D(N254), .Q(
        \REGISTERS[12][10] ) );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(n36310), .D(N253), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(n36310), .D(N252), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(n36310), .D(N251), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(N294), .D(N250), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(n36310), .D(N249), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(n36310), .D(N248), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(n36310), .D(N247), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(n36310), .D(N246), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(N294), .D(N245), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(n36310), .D(N244), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(N293), .D(N275), .Q(\REGISTERS[13][31] )
         );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(N293), .D(N274), .Q(\REGISTERS[13][30] )
         );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(N293), .D(N273), .Q(\REGISTERS[13][29] )
         );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(N293), .D(N272), .Q(\REGISTERS[13][28] )
         );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(N293), .D(N271), .Q(\REGISTERS[13][27] )
         );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(N293), .D(N270), .Q(\REGISTERS[13][26] )
         );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(n36311), .D(N269), .Q(
        \REGISTERS[13][25] ) );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(n36311), .D(N268), .Q(
        \REGISTERS[13][24] ) );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n36311), .D(N267), .Q(
        \REGISTERS[13][23] ) );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n36311), .D(N266), .Q(
        \REGISTERS[13][22] ) );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(N293), .D(N265), .Q(\REGISTERS[13][21] )
         );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(N293), .D(N264), .Q(\REGISTERS[13][20] )
         );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n36311), .D(N263), .Q(
        \REGISTERS[13][19] ) );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(n36311), .D(N262), .Q(
        \REGISTERS[13][18] ) );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n36311), .D(N261), .Q(
        \REGISTERS[13][17] ) );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(N293), .D(N260), .Q(\REGISTERS[13][16] )
         );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(N293), .D(N259), .Q(\REGISTERS[13][15] )
         );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(N293), .D(N258), .Q(\REGISTERS[13][14] )
         );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(N293), .D(N257), .Q(\REGISTERS[13][13] )
         );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(N293), .D(N256), .Q(\REGISTERS[13][12] )
         );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(n36311), .D(N255), .Q(
        \REGISTERS[13][11] ) );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n36311), .D(N254), .Q(
        \REGISTERS[13][10] ) );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(n36311), .D(N253), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(n36311), .D(N252), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n36311), .D(N251), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(N293), .D(N250), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(n36311), .D(N249), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(n36311), .D(N248), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(n36311), .D(N247), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(n36311), .D(N246), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(N293), .D(N245), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(n36311), .D(N244), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(N292), .D(N275), .Q(\REGISTERS[14][31] )
         );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(N292), .D(N274), .Q(\REGISTERS[14][30] )
         );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(N292), .D(N273), .Q(\REGISTERS[14][29] )
         );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(N292), .D(N272), .Q(\REGISTERS[14][28] )
         );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(N292), .D(N271), .Q(\REGISTERS[14][27] )
         );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(N292), .D(N270), .Q(\REGISTERS[14][26] )
         );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(n36312), .D(N269), .Q(
        \REGISTERS[14][25] ) );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(n36312), .D(N268), .Q(
        \REGISTERS[14][24] ) );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n36312), .D(N267), .Q(
        \REGISTERS[14][23] ) );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n36312), .D(N266), .Q(
        \REGISTERS[14][22] ) );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(N292), .D(N265), .Q(\REGISTERS[14][21] )
         );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(N292), .D(N264), .Q(\REGISTERS[14][20] )
         );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n36312), .D(N263), .Q(
        \REGISTERS[14][19] ) );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(n36312), .D(N262), .Q(
        \REGISTERS[14][18] ) );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n36312), .D(N261), .Q(
        \REGISTERS[14][17] ) );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(N292), .D(N260), .Q(\REGISTERS[14][16] )
         );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(N292), .D(N259), .Q(\REGISTERS[14][15] )
         );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(N292), .D(N258), .Q(\REGISTERS[14][14] )
         );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(N292), .D(N257), .Q(\REGISTERS[14][13] )
         );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(N292), .D(N256), .Q(\REGISTERS[14][12] )
         );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(n36312), .D(N255), .Q(
        \REGISTERS[14][11] ) );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n36312), .D(N254), .Q(
        \REGISTERS[14][10] ) );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(n36312), .D(N253), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(n36312), .D(N252), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n36312), .D(N251), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(N292), .D(N250), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(n36312), .D(N249), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(n36312), .D(N248), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(n36312), .D(N247), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(n36312), .D(N246), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(N292), .D(N245), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(n36312), .D(N244), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(N291), .D(N275), .Q(\REGISTERS[15][31] )
         );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(N291), .D(N274), .Q(\REGISTERS[15][30] )
         );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(N291), .D(N273), .Q(\REGISTERS[15][29] )
         );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(N291), .D(N272), .Q(\REGISTERS[15][28] )
         );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(N291), .D(N271), .Q(\REGISTERS[15][27] )
         );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(N291), .D(N270), .Q(\REGISTERS[15][26] )
         );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(n36313), .D(N269), .Q(
        \REGISTERS[15][25] ) );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(n36313), .D(N268), .Q(
        \REGISTERS[15][24] ) );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n36313), .D(N267), .Q(
        \REGISTERS[15][23] ) );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n36313), .D(N266), .Q(
        \REGISTERS[15][22] ) );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(N291), .D(N265), .Q(\REGISTERS[15][21] )
         );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(N291), .D(N264), .Q(\REGISTERS[15][20] )
         );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n36313), .D(N263), .Q(
        \REGISTERS[15][19] ) );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(n36313), .D(N262), .Q(
        \REGISTERS[15][18] ) );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n36313), .D(N261), .Q(
        \REGISTERS[15][17] ) );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(N291), .D(N260), .Q(\REGISTERS[15][16] )
         );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(N291), .D(N259), .Q(\REGISTERS[15][15] )
         );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(N291), .D(N258), .Q(\REGISTERS[15][14] )
         );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(N291), .D(N257), .Q(\REGISTERS[15][13] )
         );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(N291), .D(N256), .Q(\REGISTERS[15][12] )
         );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(n36313), .D(N255), .Q(
        \REGISTERS[15][11] ) );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n36313), .D(N254), .Q(
        \REGISTERS[15][10] ) );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(n36313), .D(N253), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(n36313), .D(N252), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n36313), .D(N251), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(N291), .D(N250), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(n36313), .D(N249), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(n36313), .D(N248), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(n36313), .D(N247), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(n36313), .D(N246), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(N291), .D(N245), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(n36313), .D(N244), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(N290), .D(N275), .Q(\REGISTERS[16][31] )
         );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(N290), .D(N274), .Q(\REGISTERS[16][30] )
         );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(N290), .D(N273), .Q(\REGISTERS[16][29] )
         );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(N290), .D(N272), .Q(\REGISTERS[16][28] )
         );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(N290), .D(N271), .Q(\REGISTERS[16][27] )
         );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(N290), .D(N270), .Q(\REGISTERS[16][26] )
         );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(n36314), .D(N269), .Q(
        \REGISTERS[16][25] ) );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(n36314), .D(N268), .Q(
        \REGISTERS[16][24] ) );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n36314), .D(N267), .Q(
        \REGISTERS[16][23] ) );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n36314), .D(N266), .Q(
        \REGISTERS[16][22] ) );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(N290), .D(N265), .Q(\REGISTERS[16][21] )
         );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(N290), .D(N264), .Q(\REGISTERS[16][20] )
         );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n36314), .D(N263), .Q(
        \REGISTERS[16][19] ) );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(n36314), .D(N262), .Q(
        \REGISTERS[16][18] ) );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n36314), .D(N261), .Q(
        \REGISTERS[16][17] ) );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(N290), .D(N260), .Q(\REGISTERS[16][16] )
         );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(N290), .D(N259), .Q(\REGISTERS[16][15] )
         );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(N290), .D(N258), .Q(\REGISTERS[16][14] )
         );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(N290), .D(N257), .Q(\REGISTERS[16][13] )
         );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(N290), .D(N256), .Q(\REGISTERS[16][12] )
         );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(n36314), .D(N255), .Q(
        \REGISTERS[16][11] ) );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n36314), .D(N254), .Q(
        \REGISTERS[16][10] ) );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(n36314), .D(N253), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(n36314), .D(N252), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n36314), .D(N251), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(N290), .D(N250), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(n36314), .D(N249), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(n36314), .D(N248), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(n36314), .D(N247), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(n36314), .D(N246), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(N290), .D(N245), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(n36314), .D(N244), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(N289), .D(N275), .Q(\REGISTERS[17][31] )
         );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(N289), .D(N274), .Q(\REGISTERS[17][30] )
         );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(N289), .D(N273), .Q(\REGISTERS[17][29] )
         );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(N289), .D(N272), .Q(\REGISTERS[17][28] )
         );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(N289), .D(N271), .Q(\REGISTERS[17][27] )
         );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(N289), .D(N270), .Q(\REGISTERS[17][26] )
         );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(n36315), .D(N269), .Q(
        \REGISTERS[17][25] ) );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(n36315), .D(N268), .Q(
        \REGISTERS[17][24] ) );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n36315), .D(N267), .Q(
        \REGISTERS[17][23] ) );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n36315), .D(N266), .Q(
        \REGISTERS[17][22] ) );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(N289), .D(N265), .Q(\REGISTERS[17][21] )
         );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(N289), .D(N264), .Q(\REGISTERS[17][20] )
         );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n36315), .D(N263), .Q(
        \REGISTERS[17][19] ) );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(n36315), .D(N262), .Q(
        \REGISTERS[17][18] ) );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n36315), .D(N261), .Q(
        \REGISTERS[17][17] ) );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(N289), .D(N260), .Q(\REGISTERS[17][16] )
         );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(N289), .D(N259), .Q(\REGISTERS[17][15] )
         );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(N289), .D(N258), .Q(\REGISTERS[17][14] )
         );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(N289), .D(N257), .Q(\REGISTERS[17][13] )
         );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(N289), .D(N256), .Q(\REGISTERS[17][12] )
         );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(n36315), .D(N255), .Q(
        \REGISTERS[17][11] ) );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n36315), .D(N254), .Q(
        \REGISTERS[17][10] ) );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(n36315), .D(N253), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(n36315), .D(N252), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n36315), .D(N251), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(N289), .D(N250), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(n36315), .D(N249), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(n36315), .D(N248), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(n36315), .D(N247), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(n36315), .D(N246), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(N289), .D(N245), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(n36315), .D(N244), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(N288), .D(N275), .Q(\REGISTERS[18][31] )
         );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(N288), .D(N274), .Q(\REGISTERS[18][30] )
         );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(N288), .D(N273), .Q(\REGISTERS[18][29] )
         );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(N288), .D(N272), .Q(\REGISTERS[18][28] )
         );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(N288), .D(N271), .Q(\REGISTERS[18][27] )
         );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(N288), .D(N270), .Q(\REGISTERS[18][26] )
         );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(n36316), .D(N269), .Q(
        \REGISTERS[18][25] ) );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(n36316), .D(N268), .Q(
        \REGISTERS[18][24] ) );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n36316), .D(N267), .Q(
        \REGISTERS[18][23] ) );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n36316), .D(N266), .Q(
        \REGISTERS[18][22] ) );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(N288), .D(N265), .Q(\REGISTERS[18][21] )
         );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(N288), .D(N264), .Q(\REGISTERS[18][20] )
         );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n36316), .D(N263), .Q(
        \REGISTERS[18][19] ) );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(n36316), .D(N262), .Q(
        \REGISTERS[18][18] ) );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n36316), .D(N261), .Q(
        \REGISTERS[18][17] ) );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(N288), .D(N260), .Q(\REGISTERS[18][16] )
         );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(N288), .D(N259), .Q(\REGISTERS[18][15] )
         );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(N288), .D(N258), .Q(\REGISTERS[18][14] )
         );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(N288), .D(N257), .Q(\REGISTERS[18][13] )
         );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(N288), .D(N256), .Q(\REGISTERS[18][12] )
         );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(n36316), .D(N255), .Q(
        \REGISTERS[18][11] ) );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n36316), .D(N254), .Q(
        \REGISTERS[18][10] ) );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(n36316), .D(N253), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(n36316), .D(N252), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n36316), .D(N251), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(N288), .D(N250), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(n36316), .D(N249), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(n36316), .D(N248), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(n36316), .D(N247), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(n36316), .D(N246), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(N288), .D(N245), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(n36316), .D(N244), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(N287), .D(N275), .Q(\REGISTERS[19][31] )
         );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(N287), .D(N274), .Q(\REGISTERS[19][30] )
         );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(N287), .D(N273), .Q(\REGISTERS[19][29] )
         );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(N287), .D(N272), .Q(\REGISTERS[19][28] )
         );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(N287), .D(N271), .Q(\REGISTERS[19][27] )
         );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(N287), .D(N270), .Q(\REGISTERS[19][26] )
         );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(n36317), .D(N269), .Q(
        \REGISTERS[19][25] ) );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(n36317), .D(N268), .Q(
        \REGISTERS[19][24] ) );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n36317), .D(N267), .Q(
        \REGISTERS[19][23] ) );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n36317), .D(N266), .Q(
        \REGISTERS[19][22] ) );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(N287), .D(N265), .Q(\REGISTERS[19][21] )
         );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(N287), .D(N264), .Q(\REGISTERS[19][20] )
         );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n36317), .D(N263), .Q(
        \REGISTERS[19][19] ) );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(n36317), .D(N262), .Q(
        \REGISTERS[19][18] ) );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n36317), .D(N261), .Q(
        \REGISTERS[19][17] ) );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(N287), .D(N260), .Q(\REGISTERS[19][16] )
         );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(N287), .D(N259), .Q(\REGISTERS[19][15] )
         );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(N287), .D(N258), .Q(\REGISTERS[19][14] )
         );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(N287), .D(N257), .Q(\REGISTERS[19][13] )
         );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(N287), .D(N256), .Q(\REGISTERS[19][12] )
         );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(n36317), .D(N255), .Q(
        \REGISTERS[19][11] ) );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n36317), .D(N254), .Q(
        \REGISTERS[19][10] ) );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(n36317), .D(N253), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(n36317), .D(N252), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n36317), .D(N251), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(N287), .D(N250), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(n36317), .D(N249), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(n36317), .D(N248), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(n36317), .D(N247), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(n36317), .D(N246), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(N287), .D(N245), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(n36317), .D(N244), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(N286), .D(N275), .Q(\REGISTERS[20][31] )
         );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(N286), .D(N274), .Q(\REGISTERS[20][30] )
         );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(N286), .D(N273), .Q(\REGISTERS[20][29] )
         );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(N286), .D(N272), .Q(\REGISTERS[20][28] )
         );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(N286), .D(N271), .Q(\REGISTERS[20][27] )
         );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(N286), .D(N270), .Q(\REGISTERS[20][26] )
         );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(n36318), .D(N269), .Q(
        \REGISTERS[20][25] ) );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(n36318), .D(N268), .Q(
        \REGISTERS[20][24] ) );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n36318), .D(N267), .Q(
        \REGISTERS[20][23] ) );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n36318), .D(N266), .Q(
        \REGISTERS[20][22] ) );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(N286), .D(N265), .Q(\REGISTERS[20][21] )
         );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(N286), .D(N264), .Q(\REGISTERS[20][20] )
         );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n36318), .D(N263), .Q(
        \REGISTERS[20][19] ) );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(n36318), .D(N262), .Q(
        \REGISTERS[20][18] ) );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n36318), .D(N261), .Q(
        \REGISTERS[20][17] ) );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(N286), .D(N260), .Q(\REGISTERS[20][16] )
         );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(N286), .D(N259), .Q(\REGISTERS[20][15] )
         );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(N286), .D(N258), .Q(\REGISTERS[20][14] )
         );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(N286), .D(N257), .Q(\REGISTERS[20][13] )
         );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(N286), .D(N256), .Q(\REGISTERS[20][12] )
         );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(n36318), .D(N255), .Q(
        \REGISTERS[20][11] ) );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n36318), .D(N254), .Q(
        \REGISTERS[20][10] ) );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(n36318), .D(N253), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(n36318), .D(N252), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n36318), .D(N251), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(N286), .D(N250), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(n36318), .D(N249), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(n36318), .D(N248), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(n36318), .D(N247), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(n36318), .D(N246), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(N286), .D(N245), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(n36318), .D(N244), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(N285), .D(N275), .Q(\REGISTERS[21][31] )
         );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(N285), .D(N274), .Q(\REGISTERS[21][30] )
         );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(N285), .D(N273), .Q(\REGISTERS[21][29] )
         );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(N285), .D(N272), .Q(\REGISTERS[21][28] )
         );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(N285), .D(N271), .Q(\REGISTERS[21][27] )
         );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(N285), .D(N270), .Q(\REGISTERS[21][26] )
         );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(n36319), .D(N269), .Q(
        \REGISTERS[21][25] ) );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(n36319), .D(N268), .Q(
        \REGISTERS[21][24] ) );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n36319), .D(N267), .Q(
        \REGISTERS[21][23] ) );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n36319), .D(N266), .Q(
        \REGISTERS[21][22] ) );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(N285), .D(N265), .Q(\REGISTERS[21][21] )
         );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(N285), .D(N264), .Q(\REGISTERS[21][20] )
         );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n36319), .D(N263), .Q(
        \REGISTERS[21][19] ) );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(n36319), .D(N262), .Q(
        \REGISTERS[21][18] ) );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n36319), .D(N261), .Q(
        \REGISTERS[21][17] ) );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(N285), .D(N260), .Q(\REGISTERS[21][16] )
         );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(N285), .D(N259), .Q(\REGISTERS[21][15] )
         );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(N285), .D(N258), .Q(\REGISTERS[21][14] )
         );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(N285), .D(N257), .Q(\REGISTERS[21][13] )
         );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(N285), .D(N256), .Q(\REGISTERS[21][12] )
         );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(n36319), .D(N255), .Q(
        \REGISTERS[21][11] ) );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n36319), .D(N254), .Q(
        \REGISTERS[21][10] ) );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(n36319), .D(N253), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(n36319), .D(N252), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n36319), .D(N251), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(N285), .D(N250), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(n36319), .D(N249), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(n36319), .D(N248), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(n36319), .D(N247), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(n36319), .D(N246), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(N285), .D(N245), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(n36319), .D(N244), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(N284), .D(N275), .Q(\REGISTERS[22][31] )
         );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(N284), .D(N274), .Q(\REGISTERS[22][30] )
         );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(N284), .D(N273), .Q(\REGISTERS[22][29] )
         );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(N284), .D(N272), .Q(\REGISTERS[22][28] )
         );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(N284), .D(N271), .Q(\REGISTERS[22][27] )
         );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(N284), .D(N270), .Q(\REGISTERS[22][26] )
         );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(n36320), .D(N269), .Q(
        \REGISTERS[22][25] ) );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(n36320), .D(N268), .Q(
        \REGISTERS[22][24] ) );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n36320), .D(N267), .Q(
        \REGISTERS[22][23] ) );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n36320), .D(N266), .Q(
        \REGISTERS[22][22] ) );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(N284), .D(N265), .Q(\REGISTERS[22][21] )
         );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(N284), .D(N264), .Q(\REGISTERS[22][20] )
         );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n36320), .D(N263), .Q(
        \REGISTERS[22][19] ) );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(n36320), .D(N262), .Q(
        \REGISTERS[22][18] ) );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n36320), .D(N261), .Q(
        \REGISTERS[22][17] ) );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(N284), .D(N260), .Q(\REGISTERS[22][16] )
         );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(N284), .D(N259), .Q(\REGISTERS[22][15] )
         );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(N284), .D(N258), .Q(\REGISTERS[22][14] )
         );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(N284), .D(N257), .Q(\REGISTERS[22][13] )
         );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(N284), .D(N256), .Q(\REGISTERS[22][12] )
         );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(n36320), .D(N255), .Q(
        \REGISTERS[22][11] ) );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n36320), .D(N254), .Q(
        \REGISTERS[22][10] ) );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(n36320), .D(N253), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(n36320), .D(N252), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n36320), .D(N251), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(N284), .D(N250), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(n36320), .D(N249), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(n36320), .D(N248), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(n36320), .D(N247), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(n36320), .D(N246), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(N284), .D(N245), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(n36320), .D(N244), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(N283), .D(N275), .Q(\REGISTERS[23][31] )
         );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(N283), .D(N274), .Q(\REGISTERS[23][30] )
         );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(N283), .D(N273), .Q(\REGISTERS[23][29] )
         );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(N283), .D(N272), .Q(\REGISTERS[23][28] )
         );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(N283), .D(N271), .Q(\REGISTERS[23][27] )
         );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(N283), .D(N270), .Q(\REGISTERS[23][26] )
         );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(n36321), .D(N269), .Q(
        \REGISTERS[23][25] ) );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(n36321), .D(N268), .Q(
        \REGISTERS[23][24] ) );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n36321), .D(N267), .Q(
        \REGISTERS[23][23] ) );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n36321), .D(N266), .Q(
        \REGISTERS[23][22] ) );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(N283), .D(N265), .Q(\REGISTERS[23][21] )
         );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(N283), .D(N264), .Q(\REGISTERS[23][20] )
         );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n36321), .D(N263), .Q(
        \REGISTERS[23][19] ) );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(n36321), .D(N262), .Q(
        \REGISTERS[23][18] ) );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n36321), .D(N261), .Q(
        \REGISTERS[23][17] ) );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(N283), .D(N260), .Q(\REGISTERS[23][16] )
         );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(N283), .D(N259), .Q(\REGISTERS[23][15] )
         );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(N283), .D(N258), .Q(\REGISTERS[23][14] )
         );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(N283), .D(N257), .Q(\REGISTERS[23][13] )
         );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(N283), .D(N256), .Q(\REGISTERS[23][12] )
         );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(n36321), .D(N255), .Q(
        \REGISTERS[23][11] ) );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n36321), .D(N254), .Q(
        \REGISTERS[23][10] ) );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(n36321), .D(N253), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(n36321), .D(N252), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n36321), .D(N251), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(N283), .D(N250), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(n36321), .D(N249), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(n36321), .D(N248), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(n36321), .D(N247), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(n36321), .D(N246), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(N283), .D(N245), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(n36321), .D(N244), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(N282), .D(N275), .Q(\REGISTERS[24][31] )
         );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(N282), .D(N274), .Q(\REGISTERS[24][30] )
         );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(N282), .D(N273), .Q(\REGISTERS[24][29] )
         );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(N282), .D(N272), .Q(\REGISTERS[24][28] )
         );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(N282), .D(N271), .Q(\REGISTERS[24][27] )
         );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(N282), .D(N270), .Q(\REGISTERS[24][26] )
         );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(N282), .D(N269), .Q(\REGISTERS[24][25] )
         );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n36322), .D(N268), .Q(
        \REGISTERS[24][24] ) );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n36322), .D(N267), .Q(
        \REGISTERS[24][23] ) );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(n36322), .D(N266), .Q(
        \REGISTERS[24][22] ) );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n36322), .D(N265), .Q(
        \REGISTERS[24][21] ) );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n36322), .D(N264), .Q(
        \REGISTERS[24][20] ) );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(N282), .D(N263), .Q(\REGISTERS[24][19] )
         );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(n36322), .D(N262), .Q(
        \REGISTERS[24][18] ) );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(N282), .D(N261), .Q(\REGISTERS[24][17] )
         );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(N282), .D(N260), .Q(\REGISTERS[24][16] )
         );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n36322), .D(N259), .Q(
        \REGISTERS[24][15] ) );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(N282), .D(N258), .Q(\REGISTERS[24][14] )
         );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(N282), .D(N257), .Q(\REGISTERS[24][13] )
         );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(n36322), .D(N256), .Q(
        \REGISTERS[24][12] ) );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(N282), .D(N255), .Q(\REGISTERS[24][11] )
         );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(N282), .D(N254), .Q(\REGISTERS[24][10] )
         );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(n36322), .D(N253), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(n36322), .D(N252), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(N282), .D(N251), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n36322), .D(N250), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(n36322), .D(N249), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(n36322), .D(N248), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(n36322), .D(N247), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(n36322), .D(N246), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(n36322), .D(N245), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(n36322), .D(N244), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(N281), .D(N275), .Q(\REGISTERS[25][31] )
         );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(N281), .D(N274), .Q(\REGISTERS[25][30] )
         );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(N281), .D(N273), .Q(\REGISTERS[25][29] )
         );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(N281), .D(N272), .Q(\REGISTERS[25][28] )
         );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(N281), .D(N271), .Q(\REGISTERS[25][27] )
         );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(N281), .D(N270), .Q(\REGISTERS[25][26] )
         );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(n36323), .D(N269), .Q(
        \REGISTERS[25][25] ) );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(n36323), .D(N268), .Q(
        \REGISTERS[25][24] ) );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n36323), .D(N267), .Q(
        \REGISTERS[25][23] ) );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n36323), .D(N266), .Q(
        \REGISTERS[25][22] ) );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(N281), .D(N265), .Q(\REGISTERS[25][21] )
         );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(N281), .D(N264), .Q(\REGISTERS[25][20] )
         );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n36323), .D(N263), .Q(
        \REGISTERS[25][19] ) );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(n36323), .D(N262), .Q(
        \REGISTERS[25][18] ) );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n36323), .D(N261), .Q(
        \REGISTERS[25][17] ) );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(N281), .D(N260), .Q(\REGISTERS[25][16] )
         );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(N281), .D(N259), .Q(\REGISTERS[25][15] )
         );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(N281), .D(N258), .Q(\REGISTERS[25][14] )
         );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(N281), .D(N257), .Q(\REGISTERS[25][13] )
         );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(N281), .D(N256), .Q(\REGISTERS[25][12] )
         );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(n36323), .D(N255), .Q(
        \REGISTERS[25][11] ) );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n36323), .D(N254), .Q(
        \REGISTERS[25][10] ) );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(n36323), .D(N253), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(n36323), .D(N252), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n36323), .D(N251), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(N281), .D(N250), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(n36323), .D(N249), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(n36323), .D(N248), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(n36323), .D(N247), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(n36323), .D(N246), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(N281), .D(N245), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(n36323), .D(N244), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(N280), .D(N275), .Q(\REGISTERS[26][31] )
         );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(N280), .D(N274), .Q(\REGISTERS[26][30] )
         );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(N280), .D(N273), .Q(\REGISTERS[26][29] )
         );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(N280), .D(N272), .Q(\REGISTERS[26][28] )
         );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(N280), .D(N271), .Q(\REGISTERS[26][27] )
         );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(N280), .D(N270), .Q(\REGISTERS[26][26] )
         );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(n36324), .D(N269), .Q(
        \REGISTERS[26][25] ) );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(n36324), .D(N268), .Q(
        \REGISTERS[26][24] ) );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n36324), .D(N267), .Q(
        \REGISTERS[26][23] ) );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n36324), .D(N266), .Q(
        \REGISTERS[26][22] ) );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(N280), .D(N265), .Q(\REGISTERS[26][21] )
         );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(N280), .D(N264), .Q(\REGISTERS[26][20] )
         );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n36324), .D(N263), .Q(
        \REGISTERS[26][19] ) );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(n36324), .D(N262), .Q(
        \REGISTERS[26][18] ) );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n36324), .D(N261), .Q(
        \REGISTERS[26][17] ) );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(N280), .D(N260), .Q(\REGISTERS[26][16] )
         );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(N280), .D(N259), .Q(\REGISTERS[26][15] )
         );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(N280), .D(N258), .Q(\REGISTERS[26][14] )
         );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(N280), .D(N257), .Q(\REGISTERS[26][13] )
         );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(N280), .D(N256), .Q(\REGISTERS[26][12] )
         );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(n36324), .D(N255), .Q(
        \REGISTERS[26][11] ) );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n36324), .D(N254), .Q(
        \REGISTERS[26][10] ) );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(n36324), .D(N253), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(n36324), .D(N252), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n36324), .D(N251), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(N280), .D(N250), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(n36324), .D(N249), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(n36324), .D(N248), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(n36324), .D(N247), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(n36324), .D(N246), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(N280), .D(N245), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(n36324), .D(N244), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(N279), .D(N275), .Q(\REGISTERS[27][31] )
         );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(N279), .D(N274), .Q(\REGISTERS[27][30] )
         );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(N279), .D(N273), .Q(\REGISTERS[27][29] )
         );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(N279), .D(N272), .Q(\REGISTERS[27][28] )
         );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(N279), .D(N271), .Q(\REGISTERS[27][27] )
         );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(N279), .D(N270), .Q(\REGISTERS[27][26] )
         );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(n36325), .D(N269), .Q(
        \REGISTERS[27][25] ) );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(n36325), .D(N268), .Q(
        \REGISTERS[27][24] ) );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n36325), .D(N267), .Q(
        \REGISTERS[27][23] ) );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n36325), .D(N266), .Q(
        \REGISTERS[27][22] ) );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(N279), .D(N265), .Q(\REGISTERS[27][21] )
         );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(N279), .D(N264), .Q(\REGISTERS[27][20] )
         );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n36325), .D(N263), .Q(
        \REGISTERS[27][19] ) );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(n36325), .D(N262), .Q(
        \REGISTERS[27][18] ) );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n36325), .D(N261), .Q(
        \REGISTERS[27][17] ) );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(N279), .D(N260), .Q(\REGISTERS[27][16] )
         );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(N279), .D(N259), .Q(\REGISTERS[27][15] )
         );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(N279), .D(N258), .Q(\REGISTERS[27][14] )
         );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(N279), .D(N257), .Q(\REGISTERS[27][13] )
         );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(N279), .D(N256), .Q(\REGISTERS[27][12] )
         );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(n36325), .D(N255), .Q(
        \REGISTERS[27][11] ) );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n36325), .D(N254), .Q(
        \REGISTERS[27][10] ) );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(n36325), .D(N253), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(n36325), .D(N252), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n36325), .D(N251), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(N279), .D(N250), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(n36325), .D(N249), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(n36325), .D(N248), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(n36325), .D(N247), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(n36325), .D(N246), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(N279), .D(N245), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(n36325), .D(N244), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(N278), .D(N275), .Q(\REGISTERS[28][31] )
         );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(N278), .D(N274), .Q(\REGISTERS[28][30] )
         );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(N278), .D(N273), .Q(\REGISTERS[28][29] )
         );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(N278), .D(N272), .Q(\REGISTERS[28][28] )
         );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(N278), .D(N271), .Q(\REGISTERS[28][27] )
         );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(N278), .D(N270), .Q(\REGISTERS[28][26] )
         );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(n36326), .D(N269), .Q(
        \REGISTERS[28][25] ) );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(n36326), .D(N268), .Q(
        \REGISTERS[28][24] ) );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n36326), .D(N267), .Q(
        \REGISTERS[28][23] ) );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n36326), .D(N266), .Q(
        \REGISTERS[28][22] ) );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(N278), .D(N265), .Q(\REGISTERS[28][21] )
         );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(N278), .D(N264), .Q(\REGISTERS[28][20] )
         );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n36326), .D(N263), .Q(
        \REGISTERS[28][19] ) );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(n36326), .D(N262), .Q(
        \REGISTERS[28][18] ) );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n36326), .D(N261), .Q(
        \REGISTERS[28][17] ) );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(N278), .D(N260), .Q(\REGISTERS[28][16] )
         );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(N278), .D(N259), .Q(\REGISTERS[28][15] )
         );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(N278), .D(N258), .Q(\REGISTERS[28][14] )
         );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(N278), .D(N257), .Q(\REGISTERS[28][13] )
         );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(N278), .D(N256), .Q(\REGISTERS[28][12] )
         );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(n36326), .D(N255), .Q(
        \REGISTERS[28][11] ) );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n36326), .D(N254), .Q(
        \REGISTERS[28][10] ) );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(n36326), .D(N253), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(n36326), .D(N252), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n36326), .D(N251), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(N278), .D(N250), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(n36326), .D(N249), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(n36326), .D(N248), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(n36326), .D(N247), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(n36326), .D(N246), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(N278), .D(N245), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(n36326), .D(N244), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(N277), .D(N275), .Q(\REGISTERS[29][31] )
         );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(N277), .D(N274), .Q(\REGISTERS[29][30] )
         );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(N277), .D(N273), .Q(\REGISTERS[29][29] )
         );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(N277), .D(N272), .Q(\REGISTERS[29][28] )
         );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(N277), .D(N271), .Q(\REGISTERS[29][27] )
         );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(N277), .D(N270), .Q(\REGISTERS[29][26] )
         );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(n36327), .D(N269), .Q(
        \REGISTERS[29][25] ) );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(n36327), .D(N268), .Q(
        \REGISTERS[29][24] ) );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n36327), .D(N267), .Q(
        \REGISTERS[29][23] ) );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n36327), .D(N266), .Q(
        \REGISTERS[29][22] ) );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(N277), .D(N265), .Q(\REGISTERS[29][21] )
         );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(N277), .D(N264), .Q(\REGISTERS[29][20] )
         );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n36327), .D(N263), .Q(
        \REGISTERS[29][19] ) );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(n36327), .D(N262), .Q(
        \REGISTERS[29][18] ) );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n36327), .D(N261), .Q(
        \REGISTERS[29][17] ) );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(N277), .D(N260), .Q(\REGISTERS[29][16] )
         );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(N277), .D(N259), .Q(\REGISTERS[29][15] )
         );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(N277), .D(N258), .Q(\REGISTERS[29][14] )
         );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(N277), .D(N257), .Q(\REGISTERS[29][13] )
         );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(N277), .D(N256), .Q(\REGISTERS[29][12] )
         );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(n36327), .D(N255), .Q(
        \REGISTERS[29][11] ) );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n36327), .D(N254), .Q(
        \REGISTERS[29][10] ) );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(n36327), .D(N253), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(n36327), .D(N252), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n36327), .D(N251), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(N277), .D(N250), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(n36327), .D(N249), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(n36327), .D(N248), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(n36327), .D(N247), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(n36327), .D(N246), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(N277), .D(N245), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(n36327), .D(N244), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(N276), .D(N275), .Q(\REGISTERS[30][31] )
         );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(N276), .D(N274), .Q(\REGISTERS[30][30] )
         );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(N276), .D(N273), .Q(\REGISTERS[30][29] )
         );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(N276), .D(N272), .Q(\REGISTERS[30][28] )
         );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(N276), .D(N271), .Q(\REGISTERS[30][27] )
         );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(N276), .D(N270), .Q(\REGISTERS[30][26] )
         );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(n36328), .D(N269), .Q(
        \REGISTERS[30][25] ) );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(n36328), .D(N268), .Q(
        \REGISTERS[30][24] ) );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n36328), .D(N267), .Q(
        \REGISTERS[30][23] ) );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n36328), .D(N266), .Q(
        \REGISTERS[30][22] ) );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(N276), .D(N265), .Q(\REGISTERS[30][21] )
         );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(N276), .D(N264), .Q(\REGISTERS[30][20] )
         );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n36328), .D(N263), .Q(
        \REGISTERS[30][19] ) );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(n36328), .D(N262), .Q(
        \REGISTERS[30][18] ) );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n36328), .D(N261), .Q(
        \REGISTERS[30][17] ) );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(N276), .D(N260), .Q(\REGISTERS[30][16] )
         );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(N276), .D(N259), .Q(\REGISTERS[30][15] )
         );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(N276), .D(N258), .Q(\REGISTERS[30][14] )
         );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(N276), .D(N257), .Q(\REGISTERS[30][13] )
         );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(N276), .D(N256), .Q(\REGISTERS[30][12] )
         );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(n36328), .D(N255), .Q(
        \REGISTERS[30][11] ) );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n36328), .D(N254), .Q(
        \REGISTERS[30][10] ) );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(n36328), .D(N253), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(n36328), .D(N252), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n36328), .D(N251), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(N276), .D(N250), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(n36328), .D(N249), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(n36328), .D(N248), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(n36328), .D(N247), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(n36328), .D(N246), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(N276), .D(N245), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(n36328), .D(N244), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(N243), .D(N275), .Q(\REGISTERS[31][31] )
         );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(N243), .D(N274), .Q(\REGISTERS[31][30] )
         );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(N243), .D(N273), .Q(\REGISTERS[31][29] )
         );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(N243), .D(N272), .Q(\REGISTERS[31][28] )
         );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(N243), .D(N271), .Q(\REGISTERS[31][27] )
         );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(N243), .D(N270), .Q(\REGISTERS[31][26] )
         );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(N243), .D(N269), .Q(\REGISTERS[31][25] )
         );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(N243), .D(N268), .Q(\REGISTERS[31][24] )
         );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(N243), .D(N267), .Q(\REGISTERS[31][23] )
         );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(N243), .D(N266), .Q(\REGISTERS[31][22] )
         );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n36329), .D(N265), .Q(
        \REGISTERS[31][21] ) );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(n36329), .D(N264), .Q(
        \REGISTERS[31][20] ) );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n36329), .D(N263), .Q(
        \REGISTERS[31][19] ) );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(n36329), .D(N262), .Q(
        \REGISTERS[31][18] ) );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n36329), .D(N261), .Q(
        \REGISTERS[31][17] ) );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(N243), .D(N260), .Q(\REGISTERS[31][16] )
         );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(N243), .D(N259), .Q(\REGISTERS[31][15] )
         );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(N243), .D(N258), .Q(\REGISTERS[31][14] )
         );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(N243), .D(N257), .Q(\REGISTERS[31][13] )
         );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(N243), .D(N256), .Q(\REGISTERS[31][12] )
         );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n36329), .D(N255), .Q(
        \REGISTERS[31][11] ) );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n36329), .D(N254), .Q(
        \REGISTERS[31][10] ) );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(n36329), .D(N253), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(n36329), .D(N252), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(n36329), .D(N251), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(n36329), .D(N250), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(n36329), .D(N249), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(n36329), .D(N248), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(n36329), .D(N247), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(n36329), .D(N246), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(n36329), .D(N245), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n36329), .D(N244), .Q(\REGISTERS[31][0] )
         );
  AOI22_X1 U3 ( .A1(\REGISTERS[9][16] ), .A2(n36283), .B1(\REGISTERS[10][16] ), 
        .B2(n36284), .ZN(n35412) );
  AOI22_X1 U4 ( .A1(\REGISTERS[18][16] ), .A2(n36285), .B1(\REGISTERS[2][16] ), 
        .B2(n36286), .ZN(n35413) );
  AOI22_X1 U5 ( .A1(\REGISTERS[31][16] ), .A2(n36287), .B1(\REGISTERS[3][16] ), 
        .B2(n36288), .ZN(n35414) );
  AOI22_X1 U6 ( .A1(\REGISTERS[8][16] ), .A2(n36289), .B1(\REGISTERS[30][16] ), 
        .B2(n36290), .ZN(n35415) );
  NAND4_X1 U7 ( .A1(n35412), .A2(n35413), .A3(n35414), .A4(n35415), .ZN(n35416) );
  AOI22_X1 U8 ( .A1(\REGISTERS[29][16] ), .A2(n36291), .B1(\REGISTERS[11][16] ), .B2(n36292), .ZN(n35417) );
  AOI22_X1 U9 ( .A1(\REGISTERS[16][16] ), .A2(n36293), .B1(\REGISTERS[1][16] ), 
        .B2(n36294), .ZN(n35418) );
  AOI22_X1 U10 ( .A1(\REGISTERS[24][16] ), .A2(n36295), .B1(
        \REGISTERS[12][16] ), .B2(n36296), .ZN(n35419) );
  AOI22_X1 U11 ( .A1(\REGISTERS[15][16] ), .A2(n36297), .B1(
        \REGISTERS[20][16] ), .B2(n36298), .ZN(n35420) );
  NAND4_X1 U12 ( .A1(n35417), .A2(n35418), .A3(n35419), .A4(n35420), .ZN(
        n35421) );
  AOI22_X1 U13 ( .A1(\REGISTERS[22][16] ), .A2(n36268), .B1(\REGISTERS[5][16] ), .B2(n36269), .ZN(n35422) );
  AOI22_X1 U14 ( .A1(\REGISTERS[21][16] ), .A2(n36270), .B1(
        \REGISTERS[25][16] ), .B2(n36271), .ZN(n35423) );
  AOI222_X1 U15 ( .A1(\REGISTERS[23][16] ), .A2(n36272), .B1(
        \REGISTERS[17][16] ), .B2(n36273), .C1(\REGISTERS[19][16] ), .C2(
        n36274), .ZN(n35424) );
  NAND3_X1 U16 ( .A1(n35422), .A2(n35423), .A3(n35424), .ZN(n35425) );
  AOI22_X1 U17 ( .A1(\REGISTERS[13][16] ), .A2(n36275), .B1(
        \REGISTERS[14][16] ), .B2(n36276), .ZN(n35426) );
  AOI22_X1 U18 ( .A1(\REGISTERS[28][16] ), .A2(n36279), .B1(\REGISTERS[6][16] ), .B2(n36280), .ZN(n35427) );
  AOI22_X1 U19 ( .A1(\REGISTERS[7][16] ), .A2(n36281), .B1(\REGISTERS[26][16] ), .B2(n36282), .ZN(n35428) );
  NAND4_X1 U20 ( .A1(n35426), .A2(n36488), .A3(n35427), .A4(n35428), .ZN(
        n35429) );
  OR4_X1 U21 ( .A1(n35416), .A2(n35421), .A3(n35425), .A4(n35429), .ZN(
        OUTA[16]) );
  AOI22_X1 U22 ( .A1(\REGISTERS[9][17] ), .A2(n36283), .B1(\REGISTERS[10][17] ), .B2(n36284), .ZN(n35430) );
  AOI22_X1 U23 ( .A1(\REGISTERS[18][17] ), .A2(n36285), .B1(\REGISTERS[2][17] ), .B2(n36286), .ZN(n35431) );
  AOI22_X1 U24 ( .A1(\REGISTERS[31][17] ), .A2(n36287), .B1(\REGISTERS[3][17] ), .B2(n36288), .ZN(n35432) );
  AOI22_X1 U25 ( .A1(\REGISTERS[8][17] ), .A2(n36289), .B1(\REGISTERS[30][17] ), .B2(n36290), .ZN(n35433) );
  NAND4_X1 U26 ( .A1(n35430), .A2(n35431), .A3(n35432), .A4(n35433), .ZN(
        n35434) );
  AOI22_X1 U27 ( .A1(\REGISTERS[29][17] ), .A2(n36291), .B1(
        \REGISTERS[11][17] ), .B2(n36292), .ZN(n35435) );
  AOI22_X1 U28 ( .A1(\REGISTERS[16][17] ), .A2(n36293), .B1(\REGISTERS[1][17] ), .B2(n36294), .ZN(n35436) );
  AOI22_X1 U29 ( .A1(\REGISTERS[24][17] ), .A2(n36295), .B1(
        \REGISTERS[12][17] ), .B2(n36296), .ZN(n35437) );
  AOI22_X1 U30 ( .A1(\REGISTERS[15][17] ), .A2(n36297), .B1(
        \REGISTERS[20][17] ), .B2(n36298), .ZN(n35438) );
  NAND4_X1 U31 ( .A1(n35435), .A2(n35436), .A3(n35437), .A4(n35438), .ZN(
        n35439) );
  AOI22_X1 U32 ( .A1(\REGISTERS[22][17] ), .A2(n36268), .B1(\REGISTERS[5][17] ), .B2(n36269), .ZN(n35440) );
  AOI22_X1 U33 ( .A1(\REGISTERS[21][17] ), .A2(n36270), .B1(
        \REGISTERS[25][17] ), .B2(n36271), .ZN(n35441) );
  AOI222_X1 U34 ( .A1(\REGISTERS[23][17] ), .A2(n36272), .B1(
        \REGISTERS[17][17] ), .B2(n36273), .C1(\REGISTERS[19][17] ), .C2(
        n36274), .ZN(n35442) );
  NAND3_X1 U35 ( .A1(n35440), .A2(n35441), .A3(n35442), .ZN(n35443) );
  AOI22_X1 U36 ( .A1(\REGISTERS[13][17] ), .A2(n36275), .B1(
        \REGISTERS[14][17] ), .B2(n36276), .ZN(n35444) );
  AOI22_X1 U37 ( .A1(\REGISTERS[28][17] ), .A2(n36279), .B1(\REGISTERS[6][17] ), .B2(n36280), .ZN(n35445) );
  AOI22_X1 U38 ( .A1(\REGISTERS[7][17] ), .A2(n36281), .B1(\REGISTERS[26][17] ), .B2(n36282), .ZN(n35446) );
  NAND4_X1 U39 ( .A1(n35444), .A2(n36489), .A3(n35445), .A4(n35446), .ZN(
        n35447) );
  OR4_X1 U40 ( .A1(n35434), .A2(n35439), .A3(n35443), .A4(n35447), .ZN(
        OUTA[17]) );
  AOI22_X1 U41 ( .A1(\REGISTERS[9][18] ), .A2(n36283), .B1(\REGISTERS[10][18] ), .B2(n36284), .ZN(n35448) );
  AOI22_X1 U42 ( .A1(\REGISTERS[18][18] ), .A2(n36285), .B1(\REGISTERS[2][18] ), .B2(n36286), .ZN(n35449) );
  AOI22_X1 U43 ( .A1(\REGISTERS[31][18] ), .A2(n36287), .B1(\REGISTERS[3][18] ), .B2(n36288), .ZN(n35450) );
  AOI22_X1 U44 ( .A1(\REGISTERS[8][18] ), .A2(n36289), .B1(\REGISTERS[30][18] ), .B2(n36290), .ZN(n35451) );
  NAND4_X1 U45 ( .A1(n35448), .A2(n35449), .A3(n35450), .A4(n35451), .ZN(
        n35452) );
  AOI22_X1 U46 ( .A1(\REGISTERS[29][18] ), .A2(n36291), .B1(
        \REGISTERS[11][18] ), .B2(n36292), .ZN(n35453) );
  AOI22_X1 U47 ( .A1(\REGISTERS[16][18] ), .A2(n36293), .B1(\REGISTERS[1][18] ), .B2(n36294), .ZN(n35454) );
  AOI22_X1 U48 ( .A1(\REGISTERS[24][18] ), .A2(n36295), .B1(
        \REGISTERS[12][18] ), .B2(n36296), .ZN(n35455) );
  AOI22_X1 U49 ( .A1(\REGISTERS[15][18] ), .A2(n36297), .B1(
        \REGISTERS[20][18] ), .B2(n36298), .ZN(n35456) );
  NAND4_X1 U50 ( .A1(n35453), .A2(n35454), .A3(n35455), .A4(n35456), .ZN(
        n35457) );
  AOI22_X1 U51 ( .A1(\REGISTERS[22][18] ), .A2(n36268), .B1(\REGISTERS[5][18] ), .B2(n36269), .ZN(n35458) );
  AOI22_X1 U52 ( .A1(\REGISTERS[21][18] ), .A2(n36270), .B1(
        \REGISTERS[25][18] ), .B2(n36271), .ZN(n35459) );
  AOI222_X1 U53 ( .A1(\REGISTERS[23][18] ), .A2(n36272), .B1(
        \REGISTERS[17][18] ), .B2(n36273), .C1(\REGISTERS[19][18] ), .C2(
        n36274), .ZN(n35460) );
  NAND3_X1 U54 ( .A1(n35458), .A2(n35459), .A3(n35460), .ZN(n35461) );
  AOI22_X1 U55 ( .A1(\REGISTERS[13][18] ), .A2(n36275), .B1(
        \REGISTERS[14][18] ), .B2(n36276), .ZN(n35462) );
  AOI22_X1 U56 ( .A1(\REGISTERS[28][18] ), .A2(n36279), .B1(\REGISTERS[6][18] ), .B2(n36280), .ZN(n35463) );
  AOI22_X1 U57 ( .A1(\REGISTERS[7][18] ), .A2(n36281), .B1(\REGISTERS[26][18] ), .B2(n36282), .ZN(n35464) );
  NAND4_X1 U58 ( .A1(n35462), .A2(n36490), .A3(n35463), .A4(n35464), .ZN(
        n35465) );
  OR4_X1 U59 ( .A1(n35452), .A2(n35457), .A3(n35461), .A4(n35465), .ZN(
        OUTA[18]) );
  AOI22_X1 U60 ( .A1(\REGISTERS[9][19] ), .A2(n36283), .B1(\REGISTERS[10][19] ), .B2(n36284), .ZN(n35466) );
  AOI22_X1 U61 ( .A1(\REGISTERS[18][19] ), .A2(n36285), .B1(\REGISTERS[2][19] ), .B2(n36286), .ZN(n35467) );
  AOI22_X1 U62 ( .A1(\REGISTERS[31][19] ), .A2(n36287), .B1(\REGISTERS[3][19] ), .B2(n36288), .ZN(n35468) );
  AOI22_X1 U63 ( .A1(\REGISTERS[8][19] ), .A2(n36289), .B1(\REGISTERS[30][19] ), .B2(n36290), .ZN(n35469) );
  NAND4_X1 U64 ( .A1(n35466), .A2(n35467), .A3(n35468), .A4(n35469), .ZN(
        n35470) );
  AOI22_X1 U65 ( .A1(\REGISTERS[29][19] ), .A2(n36291), .B1(
        \REGISTERS[11][19] ), .B2(n36292), .ZN(n35471) );
  AOI22_X1 U66 ( .A1(\REGISTERS[16][19] ), .A2(n36293), .B1(\REGISTERS[1][19] ), .B2(n36294), .ZN(n35472) );
  AOI22_X1 U67 ( .A1(\REGISTERS[24][19] ), .A2(n36295), .B1(
        \REGISTERS[12][19] ), .B2(n36296), .ZN(n35473) );
  AOI22_X1 U68 ( .A1(\REGISTERS[15][19] ), .A2(n36297), .B1(
        \REGISTERS[20][19] ), .B2(n36298), .ZN(n35474) );
  NAND4_X1 U69 ( .A1(n35471), .A2(n35472), .A3(n35473), .A4(n35474), .ZN(
        n35475) );
  AOI22_X1 U70 ( .A1(\REGISTERS[22][19] ), .A2(n36268), .B1(\REGISTERS[5][19] ), .B2(n36269), .ZN(n35476) );
  AOI22_X1 U71 ( .A1(\REGISTERS[21][19] ), .A2(n36270), .B1(
        \REGISTERS[25][19] ), .B2(n36271), .ZN(n35477) );
  AOI222_X1 U72 ( .A1(\REGISTERS[23][19] ), .A2(n36272), .B1(
        \REGISTERS[17][19] ), .B2(n36273), .C1(\REGISTERS[19][19] ), .C2(
        n36274), .ZN(n35478) );
  NAND3_X1 U73 ( .A1(n35476), .A2(n35477), .A3(n35478), .ZN(n35479) );
  AOI22_X1 U74 ( .A1(\REGISTERS[13][19] ), .A2(n36275), .B1(
        \REGISTERS[14][19] ), .B2(n36276), .ZN(n35480) );
  AOI22_X1 U75 ( .A1(\REGISTERS[28][19] ), .A2(n36279), .B1(\REGISTERS[6][19] ), .B2(n36280), .ZN(n35481) );
  AOI22_X1 U76 ( .A1(\REGISTERS[7][19] ), .A2(n36281), .B1(\REGISTERS[26][19] ), .B2(n36282), .ZN(n35482) );
  NAND4_X1 U77 ( .A1(n35480), .A2(n36491), .A3(n35481), .A4(n35482), .ZN(
        n35483) );
  OR4_X1 U78 ( .A1(n35470), .A2(n35475), .A3(n35479), .A4(n35483), .ZN(
        OUTA[19]) );
  AOI22_X1 U79 ( .A1(\REGISTERS[9][20] ), .A2(n36283), .B1(\REGISTERS[10][20] ), .B2(n36284), .ZN(n35484) );
  AOI22_X1 U80 ( .A1(\REGISTERS[18][20] ), .A2(n36285), .B1(\REGISTERS[2][20] ), .B2(n36784), .ZN(n35485) );
  AOI22_X1 U81 ( .A1(\REGISTERS[31][20] ), .A2(n36287), .B1(\REGISTERS[3][20] ), .B2(n36288), .ZN(n35486) );
  AOI22_X1 U82 ( .A1(\REGISTERS[8][20] ), .A2(n36289), .B1(\REGISTERS[30][20] ), .B2(n36290), .ZN(n35487) );
  NAND4_X1 U83 ( .A1(n35484), .A2(n35485), .A3(n35486), .A4(n35487), .ZN(
        n35488) );
  AOI22_X1 U84 ( .A1(\REGISTERS[29][20] ), .A2(n36291), .B1(
        \REGISTERS[11][20] ), .B2(n36292), .ZN(n35489) );
  AOI22_X1 U85 ( .A1(\REGISTERS[16][20] ), .A2(n36293), .B1(\REGISTERS[1][20] ), .B2(n36294), .ZN(n35490) );
  AOI22_X1 U86 ( .A1(\REGISTERS[24][20] ), .A2(n36295), .B1(
        \REGISTERS[12][20] ), .B2(n36296), .ZN(n35491) );
  AOI22_X1 U87 ( .A1(\REGISTERS[15][20] ), .A2(n36297), .B1(
        \REGISTERS[20][20] ), .B2(n36298), .ZN(n35492) );
  NAND4_X1 U88 ( .A1(n35489), .A2(n35490), .A3(n35491), .A4(n35492), .ZN(
        n35493) );
  AOI22_X1 U89 ( .A1(\REGISTERS[22][20] ), .A2(n36268), .B1(\REGISTERS[5][20] ), .B2(n36269), .ZN(n35494) );
  AOI22_X1 U90 ( .A1(\REGISTERS[21][20] ), .A2(n36270), .B1(
        \REGISTERS[25][20] ), .B2(n36271), .ZN(n35495) );
  AOI222_X1 U91 ( .A1(\REGISTERS[23][20] ), .A2(n36272), .B1(
        \REGISTERS[17][20] ), .B2(n36273), .C1(\REGISTERS[19][20] ), .C2(
        n36274), .ZN(n35496) );
  NAND3_X1 U92 ( .A1(n35494), .A2(n35495), .A3(n35496), .ZN(n35497) );
  AOI22_X1 U93 ( .A1(\REGISTERS[13][20] ), .A2(n36275), .B1(
        \REGISTERS[14][20] ), .B2(n36276), .ZN(n35498) );
  AOI22_X1 U94 ( .A1(\REGISTERS[28][20] ), .A2(n36279), .B1(\REGISTERS[6][20] ), .B2(n36280), .ZN(n35499) );
  AOI22_X1 U95 ( .A1(\REGISTERS[7][20] ), .A2(n36281), .B1(\REGISTERS[26][20] ), .B2(n36282), .ZN(n35500) );
  NAND4_X1 U96 ( .A1(n35498), .A2(n36512), .A3(n35499), .A4(n35500), .ZN(
        n35501) );
  OR4_X1 U97 ( .A1(n35488), .A2(n35493), .A3(n35497), .A4(n35501), .ZN(
        OUTA[20]) );
  AOI22_X1 U98 ( .A1(\REGISTERS[9][21] ), .A2(n36283), .B1(\REGISTERS[10][21] ), .B2(n36284), .ZN(n35502) );
  AOI22_X1 U99 ( .A1(\REGISTERS[18][21] ), .A2(n36285), .B1(\REGISTERS[2][21] ), .B2(n36286), .ZN(n35503) );
  AOI22_X1 U100 ( .A1(\REGISTERS[31][21] ), .A2(n36287), .B1(
        \REGISTERS[3][21] ), .B2(n36288), .ZN(n35504) );
  AOI22_X1 U101 ( .A1(\REGISTERS[8][21] ), .A2(n36289), .B1(
        \REGISTERS[30][21] ), .B2(n36290), .ZN(n35505) );
  NAND4_X1 U102 ( .A1(n35502), .A2(n35503), .A3(n35504), .A4(n35505), .ZN(
        n35506) );
  AOI22_X1 U103 ( .A1(\REGISTERS[29][21] ), .A2(n36291), .B1(
        \REGISTERS[11][21] ), .B2(n36292), .ZN(n35507) );
  AOI22_X1 U104 ( .A1(\REGISTERS[16][21] ), .A2(n36293), .B1(
        \REGISTERS[1][21] ), .B2(n36294), .ZN(n35508) );
  AOI22_X1 U105 ( .A1(\REGISTERS[24][21] ), .A2(n36295), .B1(
        \REGISTERS[12][21] ), .B2(n36296), .ZN(n35509) );
  AOI22_X1 U106 ( .A1(\REGISTERS[15][21] ), .A2(n36297), .B1(
        \REGISTERS[20][21] ), .B2(n36298), .ZN(n35510) );
  NAND4_X1 U107 ( .A1(n35507), .A2(n35508), .A3(n35509), .A4(n35510), .ZN(
        n35511) );
  AOI22_X1 U108 ( .A1(\REGISTERS[22][21] ), .A2(n36268), .B1(
        \REGISTERS[5][21] ), .B2(n36269), .ZN(n35512) );
  AOI22_X1 U109 ( .A1(\REGISTERS[21][21] ), .A2(n36270), .B1(
        \REGISTERS[25][21] ), .B2(n36271), .ZN(n35513) );
  AOI222_X1 U110 ( .A1(\REGISTERS[23][21] ), .A2(n36272), .B1(
        \REGISTERS[17][21] ), .B2(n36273), .C1(\REGISTERS[19][21] ), .C2(
        n36274), .ZN(n35514) );
  NAND3_X1 U111 ( .A1(n35512), .A2(n35513), .A3(n35514), .ZN(n35515) );
  AOI22_X1 U112 ( .A1(\REGISTERS[13][21] ), .A2(n36275), .B1(
        \REGISTERS[14][21] ), .B2(n36276), .ZN(n35516) );
  AOI22_X1 U113 ( .A1(\REGISTERS[28][21] ), .A2(n36279), .B1(
        \REGISTERS[6][21] ), .B2(n36280), .ZN(n35517) );
  AOI22_X1 U114 ( .A1(\REGISTERS[7][21] ), .A2(n36281), .B1(
        \REGISTERS[26][21] ), .B2(n36282), .ZN(n35518) );
  NAND4_X1 U115 ( .A1(n35516), .A2(n36513), .A3(n35517), .A4(n35518), .ZN(
        n35519) );
  OR4_X1 U116 ( .A1(n35506), .A2(n35511), .A3(n35515), .A4(n35519), .ZN(
        OUTA[21]) );
  AOI22_X1 U117 ( .A1(\REGISTERS[9][22] ), .A2(n36283), .B1(
        \REGISTERS[10][22] ), .B2(n36284), .ZN(n35520) );
  AOI22_X1 U118 ( .A1(\REGISTERS[18][22] ), .A2(n36285), .B1(
        \REGISTERS[2][22] ), .B2(n36286), .ZN(n35521) );
  AOI22_X1 U119 ( .A1(\REGISTERS[31][22] ), .A2(n36287), .B1(
        \REGISTERS[3][22] ), .B2(n36288), .ZN(n35522) );
  AOI22_X1 U120 ( .A1(\REGISTERS[8][22] ), .A2(n36289), .B1(
        \REGISTERS[30][22] ), .B2(n36290), .ZN(n35523) );
  NAND4_X1 U121 ( .A1(n35520), .A2(n35521), .A3(n35522), .A4(n35523), .ZN(
        n35524) );
  AOI22_X1 U122 ( .A1(\REGISTERS[29][22] ), .A2(n36291), .B1(
        \REGISTERS[11][22] ), .B2(n36292), .ZN(n35525) );
  AOI22_X1 U123 ( .A1(\REGISTERS[16][22] ), .A2(n36293), .B1(
        \REGISTERS[1][22] ), .B2(n36294), .ZN(n35526) );
  AOI22_X1 U124 ( .A1(\REGISTERS[24][22] ), .A2(n36295), .B1(
        \REGISTERS[12][22] ), .B2(n36296), .ZN(n35527) );
  AOI22_X1 U125 ( .A1(\REGISTERS[15][22] ), .A2(n36297), .B1(
        \REGISTERS[20][22] ), .B2(n36298), .ZN(n35528) );
  NAND4_X1 U126 ( .A1(n35525), .A2(n35526), .A3(n35527), .A4(n35528), .ZN(
        n35529) );
  AOI22_X1 U127 ( .A1(\REGISTERS[22][22] ), .A2(n36268), .B1(
        \REGISTERS[5][22] ), .B2(n36269), .ZN(n35530) );
  AOI22_X1 U128 ( .A1(\REGISTERS[21][22] ), .A2(n36270), .B1(
        \REGISTERS[25][22] ), .B2(n36271), .ZN(n35531) );
  AOI222_X1 U129 ( .A1(\REGISTERS[23][22] ), .A2(n36272), .B1(
        \REGISTERS[17][22] ), .B2(n36273), .C1(\REGISTERS[19][22] ), .C2(
        n36274), .ZN(n35532) );
  NAND3_X1 U130 ( .A1(n35530), .A2(n35531), .A3(n35532), .ZN(n35533) );
  AOI22_X1 U131 ( .A1(\REGISTERS[13][22] ), .A2(n36275), .B1(
        \REGISTERS[14][22] ), .B2(n36276), .ZN(n35534) );
  AOI22_X1 U132 ( .A1(\REGISTERS[28][22] ), .A2(n36279), .B1(
        \REGISTERS[6][22] ), .B2(n36280), .ZN(n35535) );
  AOI22_X1 U133 ( .A1(\REGISTERS[7][22] ), .A2(n36281), .B1(
        \REGISTERS[26][22] ), .B2(n36282), .ZN(n35536) );
  NAND4_X1 U134 ( .A1(n35534), .A2(n36514), .A3(n35535), .A4(n35536), .ZN(
        n35537) );
  OR4_X1 U135 ( .A1(n35524), .A2(n35529), .A3(n35533), .A4(n35537), .ZN(
        OUTA[22]) );
  AOI22_X1 U136 ( .A1(\REGISTERS[9][23] ), .A2(n36283), .B1(
        \REGISTERS[10][23] ), .B2(n36284), .ZN(n35538) );
  AOI22_X1 U137 ( .A1(\REGISTERS[18][23] ), .A2(n36285), .B1(
        \REGISTERS[2][23] ), .B2(n36286), .ZN(n35539) );
  AOI22_X1 U138 ( .A1(\REGISTERS[31][23] ), .A2(n36287), .B1(
        \REGISTERS[3][23] ), .B2(n36288), .ZN(n35540) );
  AOI22_X1 U139 ( .A1(\REGISTERS[8][23] ), .A2(n36289), .B1(
        \REGISTERS[30][23] ), .B2(n36290), .ZN(n35541) );
  NAND4_X1 U140 ( .A1(n35538), .A2(n35539), .A3(n35540), .A4(n35541), .ZN(
        n35542) );
  AOI22_X1 U141 ( .A1(\REGISTERS[29][23] ), .A2(n36291), .B1(
        \REGISTERS[11][23] ), .B2(n36292), .ZN(n35543) );
  AOI22_X1 U142 ( .A1(\REGISTERS[16][23] ), .A2(n36293), .B1(
        \REGISTERS[1][23] ), .B2(n36294), .ZN(n35544) );
  AOI22_X1 U143 ( .A1(\REGISTERS[24][23] ), .A2(n36295), .B1(
        \REGISTERS[12][23] ), .B2(n36296), .ZN(n35545) );
  AOI22_X1 U144 ( .A1(\REGISTERS[15][23] ), .A2(n36297), .B1(
        \REGISTERS[20][23] ), .B2(n36298), .ZN(n35546) );
  NAND4_X1 U145 ( .A1(n35543), .A2(n35544), .A3(n35545), .A4(n35546), .ZN(
        n35547) );
  AOI22_X1 U146 ( .A1(\REGISTERS[22][23] ), .A2(n36268), .B1(
        \REGISTERS[5][23] ), .B2(n36269), .ZN(n35548) );
  AOI22_X1 U147 ( .A1(\REGISTERS[21][23] ), .A2(n36270), .B1(
        \REGISTERS[25][23] ), .B2(n36271), .ZN(n35549) );
  AOI222_X1 U148 ( .A1(\REGISTERS[23][23] ), .A2(n36272), .B1(
        \REGISTERS[17][23] ), .B2(n36273), .C1(\REGISTERS[19][23] ), .C2(
        n36274), .ZN(n35550) );
  NAND3_X1 U149 ( .A1(n35548), .A2(n35549), .A3(n35550), .ZN(n35551) );
  AOI22_X1 U150 ( .A1(\REGISTERS[13][23] ), .A2(n36275), .B1(
        \REGISTERS[14][23] ), .B2(n36276), .ZN(n35552) );
  AOI22_X1 U151 ( .A1(\REGISTERS[28][23] ), .A2(n36279), .B1(
        \REGISTERS[6][23] ), .B2(n36280), .ZN(n35553) );
  AOI22_X1 U152 ( .A1(\REGISTERS[7][23] ), .A2(n36281), .B1(
        \REGISTERS[26][23] ), .B2(n36282), .ZN(n35554) );
  NAND4_X1 U153 ( .A1(n35552), .A2(n36515), .A3(n35553), .A4(n35554), .ZN(
        n35555) );
  OR4_X1 U154 ( .A1(n35542), .A2(n35547), .A3(n35551), .A4(n35555), .ZN(
        OUTA[23]) );
  AOI22_X1 U155 ( .A1(\REGISTERS[9][24] ), .A2(n36283), .B1(
        \REGISTERS[10][24] ), .B2(n36284), .ZN(n35556) );
  AOI22_X1 U156 ( .A1(\REGISTERS[18][24] ), .A2(n36285), .B1(
        \REGISTERS[2][24] ), .B2(n36286), .ZN(n35557) );
  AOI22_X1 U157 ( .A1(\REGISTERS[31][24] ), .A2(n36287), .B1(
        \REGISTERS[3][24] ), .B2(n36288), .ZN(n35558) );
  AOI22_X1 U158 ( .A1(\REGISTERS[8][24] ), .A2(n36289), .B1(
        \REGISTERS[30][24] ), .B2(n36290), .ZN(n35559) );
  NAND4_X1 U159 ( .A1(n35556), .A2(n35557), .A3(n35558), .A4(n35559), .ZN(
        n35560) );
  AOI22_X1 U160 ( .A1(\REGISTERS[29][24] ), .A2(n36291), .B1(
        \REGISTERS[11][24] ), .B2(n36292), .ZN(n35561) );
  AOI22_X1 U161 ( .A1(\REGISTERS[16][24] ), .A2(n36293), .B1(
        \REGISTERS[1][24] ), .B2(n36294), .ZN(n35562) );
  AOI22_X1 U162 ( .A1(\REGISTERS[24][24] ), .A2(n36295), .B1(
        \REGISTERS[12][24] ), .B2(n36296), .ZN(n35563) );
  AOI22_X1 U163 ( .A1(\REGISTERS[15][24] ), .A2(n36297), .B1(
        \REGISTERS[20][24] ), .B2(n36298), .ZN(n35564) );
  NAND4_X1 U164 ( .A1(n35561), .A2(n35562), .A3(n35563), .A4(n35564), .ZN(
        n35565) );
  AOI22_X1 U165 ( .A1(\REGISTERS[22][24] ), .A2(n36268), .B1(
        \REGISTERS[5][24] ), .B2(n36269), .ZN(n35566) );
  AOI22_X1 U166 ( .A1(\REGISTERS[21][24] ), .A2(n36270), .B1(
        \REGISTERS[25][24] ), .B2(n36271), .ZN(n35567) );
  AOI222_X1 U167 ( .A1(\REGISTERS[23][24] ), .A2(n36272), .B1(
        \REGISTERS[17][24] ), .B2(n36273), .C1(\REGISTERS[19][24] ), .C2(
        n36274), .ZN(n35568) );
  NAND3_X1 U168 ( .A1(n35566), .A2(n35567), .A3(n35568), .ZN(n35569) );
  AOI22_X1 U169 ( .A1(\REGISTERS[13][24] ), .A2(n36275), .B1(
        \REGISTERS[14][24] ), .B2(n36276), .ZN(n35570) );
  AOI22_X1 U170 ( .A1(\REGISTERS[28][24] ), .A2(n36279), .B1(
        \REGISTERS[6][24] ), .B2(n36280), .ZN(n35571) );
  AOI22_X1 U171 ( .A1(\REGISTERS[7][24] ), .A2(n36281), .B1(
        \REGISTERS[26][24] ), .B2(n36282), .ZN(n35572) );
  NAND4_X1 U172 ( .A1(n35570), .A2(n36516), .A3(n35571), .A4(n35572), .ZN(
        n35573) );
  OR4_X1 U173 ( .A1(n35560), .A2(n35565), .A3(n35569), .A4(n35573), .ZN(
        OUTA[24]) );
  AOI22_X1 U174 ( .A1(\REGISTERS[9][25] ), .A2(n36283), .B1(
        \REGISTERS[10][25] ), .B2(n36284), .ZN(n35574) );
  AOI22_X1 U175 ( .A1(\REGISTERS[18][25] ), .A2(n36285), .B1(
        \REGISTERS[2][25] ), .B2(n36286), .ZN(n35575) );
  AOI22_X1 U176 ( .A1(\REGISTERS[31][25] ), .A2(n36287), .B1(
        \REGISTERS[3][25] ), .B2(n36288), .ZN(n35576) );
  AOI22_X1 U177 ( .A1(\REGISTERS[8][25] ), .A2(n36289), .B1(
        \REGISTERS[30][25] ), .B2(n36290), .ZN(n35577) );
  NAND4_X1 U178 ( .A1(n35574), .A2(n35575), .A3(n35576), .A4(n35577), .ZN(
        n35578) );
  AOI22_X1 U179 ( .A1(\REGISTERS[29][25] ), .A2(n36291), .B1(
        \REGISTERS[11][25] ), .B2(n36292), .ZN(n35579) );
  AOI22_X1 U180 ( .A1(\REGISTERS[16][25] ), .A2(n36293), .B1(
        \REGISTERS[1][25] ), .B2(n36294), .ZN(n35580) );
  AOI22_X1 U181 ( .A1(\REGISTERS[24][25] ), .A2(n36295), .B1(
        \REGISTERS[12][25] ), .B2(n36296), .ZN(n35581) );
  AOI22_X1 U182 ( .A1(\REGISTERS[15][25] ), .A2(n36297), .B1(
        \REGISTERS[20][25] ), .B2(n36298), .ZN(n35582) );
  NAND4_X1 U183 ( .A1(n35579), .A2(n35580), .A3(n35581), .A4(n35582), .ZN(
        n35583) );
  AOI22_X1 U184 ( .A1(\REGISTERS[22][25] ), .A2(n36268), .B1(
        \REGISTERS[5][25] ), .B2(n36269), .ZN(n35584) );
  AOI22_X1 U185 ( .A1(\REGISTERS[21][25] ), .A2(n36270), .B1(
        \REGISTERS[25][25] ), .B2(n36271), .ZN(n35585) );
  AOI222_X1 U186 ( .A1(\REGISTERS[23][25] ), .A2(n36272), .B1(
        \REGISTERS[17][25] ), .B2(n36273), .C1(\REGISTERS[19][25] ), .C2(
        n36274), .ZN(n35586) );
  NAND3_X1 U187 ( .A1(n35584), .A2(n35585), .A3(n35586), .ZN(n35587) );
  AOI22_X1 U188 ( .A1(\REGISTERS[13][25] ), .A2(n36275), .B1(
        \REGISTERS[14][25] ), .B2(n36276), .ZN(n35588) );
  AOI22_X1 U189 ( .A1(\REGISTERS[28][25] ), .A2(n36279), .B1(
        \REGISTERS[6][25] ), .B2(n36280), .ZN(n35589) );
  AOI22_X1 U190 ( .A1(\REGISTERS[7][25] ), .A2(n36281), .B1(
        \REGISTERS[26][25] ), .B2(n36282), .ZN(n35590) );
  NAND4_X1 U191 ( .A1(n35588), .A2(n36517), .A3(n35589), .A4(n35590), .ZN(
        n35591) );
  OR4_X1 U192 ( .A1(n35578), .A2(n35583), .A3(n35587), .A4(n35591), .ZN(
        OUTA[25]) );
  AOI22_X1 U193 ( .A1(n36283), .A2(\REGISTERS[9][0] ), .B1(n36284), .B2(
        \REGISTERS[10][0] ), .ZN(n35592) );
  AOI22_X1 U194 ( .A1(n36285), .A2(\REGISTERS[18][0] ), .B1(n36286), .B2(
        \REGISTERS[2][0] ), .ZN(n35593) );
  AOI22_X1 U195 ( .A1(n36287), .A2(\REGISTERS[31][0] ), .B1(n36288), .B2(
        \REGISTERS[3][0] ), .ZN(n35594) );
  AOI22_X1 U196 ( .A1(n36289), .A2(\REGISTERS[8][0] ), .B1(n36290), .B2(
        \REGISTERS[30][0] ), .ZN(n35595) );
  NAND4_X1 U197 ( .A1(n35592), .A2(n35593), .A3(n35594), .A4(n35595), .ZN(
        n35596) );
  AOI22_X1 U198 ( .A1(n36291), .A2(\REGISTERS[29][0] ), .B1(n36292), .B2(
        \REGISTERS[11][0] ), .ZN(n35597) );
  AOI22_X1 U199 ( .A1(n36293), .A2(\REGISTERS[16][0] ), .B1(n36294), .B2(
        \REGISTERS[1][0] ), .ZN(n35598) );
  AOI22_X1 U200 ( .A1(n36295), .A2(\REGISTERS[24][0] ), .B1(n36296), .B2(
        \REGISTERS[12][0] ), .ZN(n35599) );
  AOI22_X1 U201 ( .A1(n36297), .A2(\REGISTERS[15][0] ), .B1(n36298), .B2(
        \REGISTERS[20][0] ), .ZN(n35600) );
  NAND4_X1 U202 ( .A1(n35597), .A2(n35598), .A3(n35599), .A4(n35600), .ZN(
        n35601) );
  AOI22_X1 U203 ( .A1(n36268), .A2(\REGISTERS[22][0] ), .B1(n36269), .B2(
        \REGISTERS[5][0] ), .ZN(n35602) );
  AOI22_X1 U204 ( .A1(n36270), .A2(\REGISTERS[21][0] ), .B1(n36271), .B2(
        \REGISTERS[25][0] ), .ZN(n35603) );
  AOI222_X1 U205 ( .A1(n36272), .A2(\REGISTERS[23][0] ), .B1(n36273), .B2(
        \REGISTERS[17][0] ), .C1(n36274), .C2(\REGISTERS[19][0] ), .ZN(n35604)
         );
  NAND3_X1 U206 ( .A1(n35602), .A2(n35603), .A3(n35604), .ZN(n35605) );
  AOI22_X1 U207 ( .A1(n36275), .A2(\REGISTERS[13][0] ), .B1(n36276), .B2(
        \REGISTERS[14][0] ), .ZN(n35606) );
  AOI22_X1 U208 ( .A1(n36279), .A2(\REGISTERS[28][0] ), .B1(n36280), .B2(
        \REGISTERS[6][0] ), .ZN(n35607) );
  AOI22_X1 U209 ( .A1(n36281), .A2(\REGISTERS[7][0] ), .B1(n36282), .B2(
        \REGISTERS[26][0] ), .ZN(n35608) );
  NAND4_X1 U210 ( .A1(n35606), .A2(n36355), .A3(n35607), .A4(n35608), .ZN(
        n35609) );
  OR4_X1 U211 ( .A1(n35596), .A2(n35601), .A3(n35605), .A4(n35609), .ZN(
        OUTA[0]) );
  AOI22_X1 U212 ( .A1(n36240), .A2(\REGISTERS[30][31] ), .B1(n36237), .B2(
        \REGISTERS[14][31] ), .ZN(n35610) );
  AOI22_X1 U213 ( .A1(n36238), .A2(\REGISTERS[3][31] ), .B1(n36242), .B2(
        \REGISTERS[4][31] ), .ZN(n35611) );
  AOI22_X1 U214 ( .A1(n36250), .A2(\REGISTERS[17][31] ), .B1(n36245), .B2(
        \REGISTERS[22][31] ), .ZN(n35612) );
  AOI22_X1 U215 ( .A1(n36260), .A2(\REGISTERS[15][31] ), .B1(n36258), .B2(
        \REGISTERS[9][31] ), .ZN(n35613) );
  NAND4_X1 U216 ( .A1(n35610), .A2(n35611), .A3(n35612), .A4(n35613), .ZN(
        n35614) );
  AOI22_X1 U217 ( .A1(n36262), .A2(\REGISTERS[16][31] ), .B1(n36263), .B2(
        \REGISTERS[25][31] ), .ZN(n35615) );
  AOI22_X1 U218 ( .A1(n36265), .A2(\REGISTERS[11][31] ), .B1(n36264), .B2(
        \REGISTERS[2][31] ), .ZN(n35616) );
  AOI22_X1 U219 ( .A1(n36855), .A2(\REGISTERS[31][31] ), .B1(n36261), .B2(
        \REGISTERS[13][31] ), .ZN(n35617) );
  AOI22_X1 U220 ( .A1(n36255), .A2(\REGISTERS[29][31] ), .B1(n36259), .B2(
        \REGISTERS[8][31] ), .ZN(n35618) );
  NAND4_X1 U221 ( .A1(n35615), .A2(n35616), .A3(n35617), .A4(n35618), .ZN(
        n35619) );
  AOI22_X1 U222 ( .A1(n36254), .A2(\REGISTERS[26][31] ), .B1(n36256), .B2(
        \REGISTERS[21][31] ), .ZN(n35620) );
  AOI22_X1 U223 ( .A1(n36251), .A2(\REGISTERS[1][31] ), .B1(n36252), .B2(
        \REGISTERS[7][31] ), .ZN(n35621) );
  AOI222_X1 U224 ( .A1(n36248), .A2(\REGISTERS[20][31] ), .B1(n36249), .B2(
        \REGISTERS[5][31] ), .C1(n36247), .C2(\REGISTERS[18][31] ), .ZN(n35622) );
  NAND3_X1 U225 ( .A1(n35620), .A2(n35621), .A3(n35622), .ZN(n35623) );
  AOI22_X1 U226 ( .A1(n36244), .A2(\REGISTERS[28][31] ), .B1(n36246), .B2(
        \REGISTERS[19][31] ), .ZN(n35624) );
  AOI22_X1 U227 ( .A1(n36243), .A2(\REGISTERS[6][31] ), .B1(n36257), .B2(
        \REGISTERS[23][31] ), .ZN(n35625) );
  AOI22_X1 U228 ( .A1(n36253), .A2(\REGISTERS[24][31] ), .B1(n36241), .B2(
        \REGISTERS[10][31] ), .ZN(n35626) );
  AOI22_X1 U229 ( .A1(n36239), .A2(\REGISTERS[12][31] ), .B1(n36266), .B2(
        \REGISTERS[27][31] ), .ZN(n35627) );
  NAND4_X1 U230 ( .A1(n35624), .A2(n35625), .A3(n35626), .A4(n35627), .ZN(
        n35628) );
  OR4_X1 U231 ( .A1(n35614), .A2(n35619), .A3(n35623), .A4(n35628), .ZN(
        OUTB[31]) );
  AOI22_X1 U232 ( .A1(n36781), .A2(\REGISTERS[9][31] ), .B1(n36782), .B2(
        \REGISTERS[10][31] ), .ZN(n35629) );
  AOI22_X1 U233 ( .A1(n36783), .A2(\REGISTERS[18][31] ), .B1(n36784), .B2(
        \REGISTERS[2][31] ), .ZN(n35630) );
  AOI22_X1 U234 ( .A1(n36786), .A2(\REGISTERS[3][31] ), .B1(n36785), .B2(
        \REGISTERS[31][31] ), .ZN(n35631) );
  AOI22_X1 U235 ( .A1(n36787), .A2(\REGISTERS[8][31] ), .B1(n36788), .B2(
        \REGISTERS[30][31] ), .ZN(n35632) );
  NAND4_X1 U236 ( .A1(n35629), .A2(n35630), .A3(n35631), .A4(n35632), .ZN(
        n35633) );
  AOI22_X1 U237 ( .A1(n36793), .A2(\REGISTERS[29][31] ), .B1(n36794), .B2(
        \REGISTERS[11][31] ), .ZN(n35634) );
  AOI22_X1 U238 ( .A1(n36795), .A2(\REGISTERS[16][31] ), .B1(n36796), .B2(
        \REGISTERS[1][31] ), .ZN(n35635) );
  AOI22_X1 U239 ( .A1(n36797), .A2(\REGISTERS[24][31] ), .B1(n36798), .B2(
        \REGISTERS[12][31] ), .ZN(n35636) );
  AOI22_X1 U240 ( .A1(n36800), .A2(\REGISTERS[20][31] ), .B1(n36799), .B2(
        \REGISTERS[15][31] ), .ZN(n35637) );
  NAND4_X1 U241 ( .A1(n35634), .A2(n35635), .A3(n35636), .A4(n35637), .ZN(
        n35638) );
  AOI22_X1 U242 ( .A1(n36759), .A2(\REGISTERS[5][31] ), .B1(n36758), .B2(
        \REGISTERS[22][31] ), .ZN(n35639) );
  AOI22_X1 U243 ( .A1(n36760), .A2(\REGISTERS[21][31] ), .B1(n36761), .B2(
        \REGISTERS[25][31] ), .ZN(n35640) );
  AOI222_X1 U244 ( .A1(n36763), .A2(\REGISTERS[17][31] ), .B1(n36762), .B2(
        \REGISTERS[23][31] ), .C1(n36764), .C2(\REGISTERS[19][31] ), .ZN(
        n35641) );
  NAND3_X1 U245 ( .A1(n35639), .A2(n35640), .A3(n35641), .ZN(n35642) );
  AOI22_X1 U246 ( .A1(n36769), .A2(\REGISTERS[13][31] ), .B1(n36770), .B2(
        \REGISTERS[14][31] ), .ZN(n35643) );
  AOI22_X1 U247 ( .A1(n36771), .A2(\REGISTERS[4][31] ), .B1(n36772), .B2(
        \REGISTERS[27][31] ), .ZN(n35644) );
  AOI22_X1 U248 ( .A1(n36773), .A2(\REGISTERS[28][31] ), .B1(n36774), .B2(
        \REGISTERS[6][31] ), .ZN(n35645) );
  AOI22_X1 U249 ( .A1(n36776), .A2(\REGISTERS[26][31] ), .B1(n36775), .B2(
        \REGISTERS[7][31] ), .ZN(n35646) );
  NAND4_X1 U250 ( .A1(n35643), .A2(n35644), .A3(n35645), .A4(n35646), .ZN(
        n35647) );
  OR4_X1 U251 ( .A1(n35633), .A2(n35638), .A3(n35642), .A4(n35647), .ZN(
        OUTA[31]) );
  AOI22_X1 U252 ( .A1(n36240), .A2(\REGISTERS[30][30] ), .B1(n36237), .B2(
        \REGISTERS[14][30] ), .ZN(n35648) );
  AOI22_X1 U253 ( .A1(n36238), .A2(\REGISTERS[3][30] ), .B1(n36242), .B2(
        \REGISTERS[4][30] ), .ZN(n35649) );
  AOI22_X1 U254 ( .A1(n36250), .A2(\REGISTERS[17][30] ), .B1(n36245), .B2(
        \REGISTERS[22][30] ), .ZN(n35650) );
  AOI22_X1 U255 ( .A1(n36260), .A2(\REGISTERS[15][30] ), .B1(n36258), .B2(
        \REGISTERS[9][30] ), .ZN(n35651) );
  NAND4_X1 U256 ( .A1(n35648), .A2(n35649), .A3(n35650), .A4(n35651), .ZN(
        n35652) );
  AOI22_X1 U257 ( .A1(n36262), .A2(\REGISTERS[16][30] ), .B1(n36263), .B2(
        \REGISTERS[25][30] ), .ZN(n35653) );
  AOI22_X1 U258 ( .A1(n36265), .A2(\REGISTERS[11][30] ), .B1(n36264), .B2(
        \REGISTERS[2][30] ), .ZN(n35654) );
  AOI22_X1 U259 ( .A1(n36267), .A2(\REGISTERS[31][30] ), .B1(n36261), .B2(
        \REGISTERS[13][30] ), .ZN(n35655) );
  AOI22_X1 U260 ( .A1(n36255), .A2(\REGISTERS[29][30] ), .B1(n36259), .B2(
        \REGISTERS[8][30] ), .ZN(n35656) );
  NAND4_X1 U261 ( .A1(n35653), .A2(n35654), .A3(n35655), .A4(n35656), .ZN(
        n35657) );
  AOI22_X1 U262 ( .A1(n36254), .A2(\REGISTERS[26][30] ), .B1(n36256), .B2(
        \REGISTERS[21][30] ), .ZN(n35658) );
  AOI22_X1 U263 ( .A1(n36251), .A2(\REGISTERS[1][30] ), .B1(n36252), .B2(
        \REGISTERS[7][30] ), .ZN(n35659) );
  AOI222_X1 U264 ( .A1(n36248), .A2(\REGISTERS[20][30] ), .B1(n36249), .B2(
        \REGISTERS[5][30] ), .C1(n36247), .C2(\REGISTERS[18][30] ), .ZN(n35660) );
  NAND3_X1 U265 ( .A1(n35658), .A2(n35659), .A3(n35660), .ZN(n35661) );
  AOI22_X1 U266 ( .A1(n36244), .A2(\REGISTERS[28][30] ), .B1(n36246), .B2(
        \REGISTERS[19][30] ), .ZN(n35662) );
  AOI22_X1 U267 ( .A1(n36243), .A2(\REGISTERS[6][30] ), .B1(n36257), .B2(
        \REGISTERS[23][30] ), .ZN(n35663) );
  AOI22_X1 U268 ( .A1(n36253), .A2(\REGISTERS[24][30] ), .B1(n36241), .B2(
        \REGISTERS[10][30] ), .ZN(n35664) );
  AOI22_X1 U269 ( .A1(n36239), .A2(\REGISTERS[12][30] ), .B1(n36266), .B2(
        \REGISTERS[27][30] ), .ZN(n35665) );
  NAND4_X1 U270 ( .A1(n35662), .A2(n35663), .A3(n35664), .A4(n35665), .ZN(
        n35666) );
  OR4_X1 U271 ( .A1(n35652), .A2(n35657), .A3(n35661), .A4(n35666), .ZN(
        OUTB[30]) );
  AOI22_X1 U272 ( .A1(n36240), .A2(\REGISTERS[30][29] ), .B1(n36237), .B2(
        \REGISTERS[14][29] ), .ZN(n35667) );
  AOI22_X1 U273 ( .A1(n36238), .A2(\REGISTERS[3][29] ), .B1(n36242), .B2(
        \REGISTERS[4][29] ), .ZN(n35668) );
  AOI22_X1 U274 ( .A1(n36250), .A2(\REGISTERS[17][29] ), .B1(n36245), .B2(
        \REGISTERS[22][29] ), .ZN(n35669) );
  AOI22_X1 U275 ( .A1(n36260), .A2(\REGISTERS[15][29] ), .B1(n36258), .B2(
        \REGISTERS[9][29] ), .ZN(n35670) );
  NAND4_X1 U276 ( .A1(n35667), .A2(n35668), .A3(n35669), .A4(n35670), .ZN(
        n35671) );
  AOI22_X1 U277 ( .A1(n36262), .A2(\REGISTERS[16][29] ), .B1(n36263), .B2(
        \REGISTERS[25][29] ), .ZN(n35672) );
  AOI22_X1 U278 ( .A1(n36265), .A2(\REGISTERS[11][29] ), .B1(n36264), .B2(
        \REGISTERS[2][29] ), .ZN(n35673) );
  AOI22_X1 U279 ( .A1(n36267), .A2(\REGISTERS[31][29] ), .B1(n36261), .B2(
        \REGISTERS[13][29] ), .ZN(n35674) );
  AOI22_X1 U280 ( .A1(n36255), .A2(\REGISTERS[29][29] ), .B1(n36259), .B2(
        \REGISTERS[8][29] ), .ZN(n35675) );
  NAND4_X1 U281 ( .A1(n35672), .A2(n35673), .A3(n35674), .A4(n35675), .ZN(
        n35676) );
  AOI22_X1 U282 ( .A1(n36254), .A2(\REGISTERS[26][29] ), .B1(n36256), .B2(
        \REGISTERS[21][29] ), .ZN(n35677) );
  AOI22_X1 U283 ( .A1(n36251), .A2(\REGISTERS[1][29] ), .B1(n36252), .B2(
        \REGISTERS[7][29] ), .ZN(n35678) );
  AOI222_X1 U284 ( .A1(n36248), .A2(\REGISTERS[20][29] ), .B1(n36249), .B2(
        \REGISTERS[5][29] ), .C1(n36247), .C2(\REGISTERS[18][29] ), .ZN(n35679) );
  NAND3_X1 U285 ( .A1(n35677), .A2(n35678), .A3(n35679), .ZN(n35680) );
  AOI22_X1 U286 ( .A1(n36244), .A2(\REGISTERS[28][29] ), .B1(n36246), .B2(
        \REGISTERS[19][29] ), .ZN(n35681) );
  AOI22_X1 U287 ( .A1(n36243), .A2(\REGISTERS[6][29] ), .B1(n36257), .B2(
        \REGISTERS[23][29] ), .ZN(n35682) );
  AOI22_X1 U288 ( .A1(n36253), .A2(\REGISTERS[24][29] ), .B1(n36241), .B2(
        \REGISTERS[10][29] ), .ZN(n35683) );
  AOI22_X1 U289 ( .A1(n36239), .A2(\REGISTERS[12][29] ), .B1(n36266), .B2(
        \REGISTERS[27][29] ), .ZN(n35684) );
  NAND4_X1 U290 ( .A1(n35681), .A2(n35682), .A3(n35683), .A4(n35684), .ZN(
        n35685) );
  OR4_X1 U291 ( .A1(n35671), .A2(n35676), .A3(n35680), .A4(n35685), .ZN(
        OUTB[29]) );
  AOI22_X1 U292 ( .A1(n36240), .A2(\REGISTERS[30][28] ), .B1(n36237), .B2(
        \REGISTERS[14][28] ), .ZN(n35686) );
  AOI22_X1 U293 ( .A1(n36238), .A2(\REGISTERS[3][28] ), .B1(n36242), .B2(
        \REGISTERS[4][28] ), .ZN(n35687) );
  AOI22_X1 U294 ( .A1(n36250), .A2(\REGISTERS[17][28] ), .B1(n36245), .B2(
        \REGISTERS[22][28] ), .ZN(n35688) );
  AOI22_X1 U295 ( .A1(n36260), .A2(\REGISTERS[15][28] ), .B1(n36258), .B2(
        \REGISTERS[9][28] ), .ZN(n35689) );
  NAND4_X1 U296 ( .A1(n35686), .A2(n35687), .A3(n35688), .A4(n35689), .ZN(
        n35690) );
  AOI22_X1 U297 ( .A1(n36262), .A2(\REGISTERS[16][28] ), .B1(n36263), .B2(
        \REGISTERS[25][28] ), .ZN(n35691) );
  AOI22_X1 U298 ( .A1(n36265), .A2(\REGISTERS[11][28] ), .B1(n36264), .B2(
        \REGISTERS[2][28] ), .ZN(n35692) );
  AOI22_X1 U299 ( .A1(n36267), .A2(\REGISTERS[31][28] ), .B1(n36261), .B2(
        \REGISTERS[13][28] ), .ZN(n35693) );
  AOI22_X1 U300 ( .A1(n36255), .A2(\REGISTERS[29][28] ), .B1(n36259), .B2(
        \REGISTERS[8][28] ), .ZN(n35694) );
  NAND4_X1 U301 ( .A1(n35691), .A2(n35692), .A3(n35693), .A4(n35694), .ZN(
        n35695) );
  AOI22_X1 U302 ( .A1(n36254), .A2(\REGISTERS[26][28] ), .B1(n36256), .B2(
        \REGISTERS[21][28] ), .ZN(n35696) );
  AOI22_X1 U303 ( .A1(n36251), .A2(\REGISTERS[1][28] ), .B1(n36252), .B2(
        \REGISTERS[7][28] ), .ZN(n35697) );
  AOI222_X1 U304 ( .A1(n36248), .A2(\REGISTERS[20][28] ), .B1(n36249), .B2(
        \REGISTERS[5][28] ), .C1(n36247), .C2(\REGISTERS[18][28] ), .ZN(n35698) );
  NAND3_X1 U305 ( .A1(n35696), .A2(n35697), .A3(n35698), .ZN(n35699) );
  AOI22_X1 U306 ( .A1(n36244), .A2(\REGISTERS[28][28] ), .B1(n36246), .B2(
        \REGISTERS[19][28] ), .ZN(n35700) );
  AOI22_X1 U307 ( .A1(n36243), .A2(\REGISTERS[6][28] ), .B1(n36257), .B2(
        \REGISTERS[23][28] ), .ZN(n35701) );
  AOI22_X1 U308 ( .A1(n36253), .A2(\REGISTERS[24][28] ), .B1(n36241), .B2(
        \REGISTERS[10][28] ), .ZN(n35702) );
  AOI22_X1 U309 ( .A1(n36239), .A2(\REGISTERS[12][28] ), .B1(n36266), .B2(
        \REGISTERS[27][28] ), .ZN(n35703) );
  NAND4_X1 U310 ( .A1(n35700), .A2(n35701), .A3(n35702), .A4(n35703), .ZN(
        n35704) );
  OR4_X1 U311 ( .A1(n35690), .A2(n35695), .A3(n35699), .A4(n35704), .ZN(
        OUTB[28]) );
  AOI22_X1 U312 ( .A1(n36240), .A2(\REGISTERS[30][27] ), .B1(n36237), .B2(
        \REGISTERS[14][27] ), .ZN(n35705) );
  AOI22_X1 U313 ( .A1(n36238), .A2(\REGISTERS[3][27] ), .B1(n36242), .B2(
        \REGISTERS[4][27] ), .ZN(n35706) );
  AOI22_X1 U314 ( .A1(n36250), .A2(\REGISTERS[17][27] ), .B1(n36245), .B2(
        \REGISTERS[22][27] ), .ZN(n35707) );
  AOI22_X1 U315 ( .A1(n36260), .A2(\REGISTERS[15][27] ), .B1(n36258), .B2(
        \REGISTERS[9][27] ), .ZN(n35708) );
  NAND4_X1 U316 ( .A1(n35705), .A2(n35706), .A3(n35707), .A4(n35708), .ZN(
        n35709) );
  AOI22_X1 U317 ( .A1(n36262), .A2(\REGISTERS[16][27] ), .B1(n36263), .B2(
        \REGISTERS[25][27] ), .ZN(n35710) );
  AOI22_X1 U318 ( .A1(n36265), .A2(\REGISTERS[11][27] ), .B1(n36264), .B2(
        \REGISTERS[2][27] ), .ZN(n35711) );
  AOI22_X1 U319 ( .A1(n36267), .A2(\REGISTERS[31][27] ), .B1(n36261), .B2(
        \REGISTERS[13][27] ), .ZN(n35712) );
  AOI22_X1 U320 ( .A1(n36255), .A2(\REGISTERS[29][27] ), .B1(n36259), .B2(
        \REGISTERS[8][27] ), .ZN(n35713) );
  NAND4_X1 U321 ( .A1(n35710), .A2(n35711), .A3(n35712), .A4(n35713), .ZN(
        n35714) );
  AOI22_X1 U322 ( .A1(n36254), .A2(\REGISTERS[26][27] ), .B1(n36256), .B2(
        \REGISTERS[21][27] ), .ZN(n35715) );
  AOI22_X1 U323 ( .A1(n36251), .A2(\REGISTERS[1][27] ), .B1(n36252), .B2(
        \REGISTERS[7][27] ), .ZN(n35716) );
  AOI222_X1 U324 ( .A1(n36248), .A2(\REGISTERS[20][27] ), .B1(n36249), .B2(
        \REGISTERS[5][27] ), .C1(n36247), .C2(\REGISTERS[18][27] ), .ZN(n35717) );
  NAND3_X1 U325 ( .A1(n35715), .A2(n35716), .A3(n35717), .ZN(n35718) );
  AOI22_X1 U326 ( .A1(n36244), .A2(\REGISTERS[28][27] ), .B1(n36246), .B2(
        \REGISTERS[19][27] ), .ZN(n35719) );
  AOI22_X1 U327 ( .A1(n36243), .A2(\REGISTERS[6][27] ), .B1(n36257), .B2(
        \REGISTERS[23][27] ), .ZN(n35720) );
  AOI22_X1 U328 ( .A1(n36253), .A2(\REGISTERS[24][27] ), .B1(n36241), .B2(
        \REGISTERS[10][27] ), .ZN(n35721) );
  AOI22_X1 U329 ( .A1(n36239), .A2(\REGISTERS[12][27] ), .B1(n36266), .B2(
        \REGISTERS[27][27] ), .ZN(n35722) );
  NAND4_X1 U330 ( .A1(n35719), .A2(n35720), .A3(n35721), .A4(n35722), .ZN(
        n35723) );
  OR4_X1 U331 ( .A1(n35709), .A2(n35714), .A3(n35718), .A4(n35723), .ZN(
        OUTB[27]) );
  AOI22_X1 U332 ( .A1(n36240), .A2(\REGISTERS[30][26] ), .B1(n36237), .B2(
        \REGISTERS[14][26] ), .ZN(n35724) );
  AOI22_X1 U333 ( .A1(n36238), .A2(\REGISTERS[3][26] ), .B1(n36242), .B2(
        \REGISTERS[4][26] ), .ZN(n35725) );
  AOI22_X1 U334 ( .A1(n36250), .A2(\REGISTERS[17][26] ), .B1(n36245), .B2(
        \REGISTERS[22][26] ), .ZN(n35726) );
  AOI22_X1 U335 ( .A1(n36260), .A2(\REGISTERS[15][26] ), .B1(n36258), .B2(
        \REGISTERS[9][26] ), .ZN(n35727) );
  NAND4_X1 U336 ( .A1(n35724), .A2(n35725), .A3(n35726), .A4(n35727), .ZN(
        n35728) );
  AOI22_X1 U337 ( .A1(n36262), .A2(\REGISTERS[16][26] ), .B1(n36263), .B2(
        \REGISTERS[25][26] ), .ZN(n35729) );
  AOI22_X1 U338 ( .A1(n36265), .A2(\REGISTERS[11][26] ), .B1(n36264), .B2(
        \REGISTERS[2][26] ), .ZN(n35730) );
  AOI22_X1 U339 ( .A1(n36267), .A2(\REGISTERS[31][26] ), .B1(n36261), .B2(
        \REGISTERS[13][26] ), .ZN(n35731) );
  AOI22_X1 U340 ( .A1(n36255), .A2(\REGISTERS[29][26] ), .B1(n36259), .B2(
        \REGISTERS[8][26] ), .ZN(n35732) );
  NAND4_X1 U341 ( .A1(n35729), .A2(n35730), .A3(n35731), .A4(n35732), .ZN(
        n35733) );
  AOI22_X1 U342 ( .A1(n36254), .A2(\REGISTERS[26][26] ), .B1(n36256), .B2(
        \REGISTERS[21][26] ), .ZN(n35734) );
  AOI22_X1 U343 ( .A1(n36251), .A2(\REGISTERS[1][26] ), .B1(n36252), .B2(
        \REGISTERS[7][26] ), .ZN(n35735) );
  AOI222_X1 U344 ( .A1(n36248), .A2(\REGISTERS[20][26] ), .B1(n36249), .B2(
        \REGISTERS[5][26] ), .C1(n36247), .C2(\REGISTERS[18][26] ), .ZN(n35736) );
  NAND3_X1 U345 ( .A1(n35734), .A2(n35735), .A3(n35736), .ZN(n35737) );
  AOI22_X1 U346 ( .A1(n36244), .A2(\REGISTERS[28][26] ), .B1(n36246), .B2(
        \REGISTERS[19][26] ), .ZN(n35738) );
  AOI22_X1 U347 ( .A1(n36243), .A2(\REGISTERS[6][26] ), .B1(n36257), .B2(
        \REGISTERS[23][26] ), .ZN(n35739) );
  AOI22_X1 U348 ( .A1(n36253), .A2(\REGISTERS[24][26] ), .B1(n36241), .B2(
        \REGISTERS[10][26] ), .ZN(n35740) );
  AOI22_X1 U349 ( .A1(n36239), .A2(\REGISTERS[12][26] ), .B1(n36266), .B2(
        \REGISTERS[27][26] ), .ZN(n35741) );
  NAND4_X1 U350 ( .A1(n35738), .A2(n35739), .A3(n35740), .A4(n35741), .ZN(
        n35742) );
  OR4_X1 U351 ( .A1(n35728), .A2(n35733), .A3(n35737), .A4(n35742), .ZN(
        OUTB[26]) );
  AOI22_X1 U352 ( .A1(n36240), .A2(\REGISTERS[30][25] ), .B1(n36237), .B2(
        \REGISTERS[14][25] ), .ZN(n35743) );
  AOI22_X1 U353 ( .A1(n36238), .A2(\REGISTERS[3][25] ), .B1(n36242), .B2(
        \REGISTERS[4][25] ), .ZN(n35744) );
  AOI22_X1 U354 ( .A1(n36250), .A2(\REGISTERS[17][25] ), .B1(n36245), .B2(
        \REGISTERS[22][25] ), .ZN(n35745) );
  AOI22_X1 U355 ( .A1(n36260), .A2(\REGISTERS[15][25] ), .B1(n36258), .B2(
        \REGISTERS[9][25] ), .ZN(n35746) );
  NAND4_X1 U356 ( .A1(n35743), .A2(n35744), .A3(n35745), .A4(n35746), .ZN(
        n35747) );
  AOI22_X1 U357 ( .A1(n36262), .A2(\REGISTERS[16][25] ), .B1(n36263), .B2(
        \REGISTERS[25][25] ), .ZN(n35748) );
  AOI22_X1 U358 ( .A1(n36265), .A2(\REGISTERS[11][25] ), .B1(n36264), .B2(
        \REGISTERS[2][25] ), .ZN(n35749) );
  AOI22_X1 U359 ( .A1(n36267), .A2(\REGISTERS[31][25] ), .B1(n36261), .B2(
        \REGISTERS[13][25] ), .ZN(n35750) );
  AOI22_X1 U360 ( .A1(n36255), .A2(\REGISTERS[29][25] ), .B1(n36259), .B2(
        \REGISTERS[8][25] ), .ZN(n35751) );
  NAND4_X1 U361 ( .A1(n35748), .A2(n35749), .A3(n35750), .A4(n35751), .ZN(
        n35752) );
  AOI22_X1 U362 ( .A1(n36254), .A2(\REGISTERS[26][25] ), .B1(n36256), .B2(
        \REGISTERS[21][25] ), .ZN(n35753) );
  AOI22_X1 U363 ( .A1(n36251), .A2(\REGISTERS[1][25] ), .B1(n36252), .B2(
        \REGISTERS[7][25] ), .ZN(n35754) );
  AOI222_X1 U364 ( .A1(n36248), .A2(\REGISTERS[20][25] ), .B1(n36249), .B2(
        \REGISTERS[5][25] ), .C1(n36247), .C2(\REGISTERS[18][25] ), .ZN(n35755) );
  NAND3_X1 U365 ( .A1(n35753), .A2(n35754), .A3(n35755), .ZN(n35756) );
  AOI22_X1 U366 ( .A1(n36244), .A2(\REGISTERS[28][25] ), .B1(n36246), .B2(
        \REGISTERS[19][25] ), .ZN(n35757) );
  AOI22_X1 U367 ( .A1(n36243), .A2(\REGISTERS[6][25] ), .B1(n36257), .B2(
        \REGISTERS[23][25] ), .ZN(n35758) );
  AOI22_X1 U368 ( .A1(n36253), .A2(\REGISTERS[24][25] ), .B1(n36241), .B2(
        \REGISTERS[10][25] ), .ZN(n35759) );
  AOI22_X1 U369 ( .A1(n36239), .A2(\REGISTERS[12][25] ), .B1(n36266), .B2(
        \REGISTERS[27][25] ), .ZN(n35760) );
  NAND4_X1 U370 ( .A1(n35757), .A2(n35758), .A3(n35759), .A4(n35760), .ZN(
        n35761) );
  OR4_X1 U371 ( .A1(n35747), .A2(n35752), .A3(n35756), .A4(n35761), .ZN(
        OUTB[25]) );
  AOI22_X1 U372 ( .A1(n36240), .A2(\REGISTERS[30][24] ), .B1(n36237), .B2(
        \REGISTERS[14][24] ), .ZN(n35762) );
  AOI22_X1 U373 ( .A1(n36238), .A2(\REGISTERS[3][24] ), .B1(n36242), .B2(
        \REGISTERS[4][24] ), .ZN(n35763) );
  AOI22_X1 U374 ( .A1(n36250), .A2(\REGISTERS[17][24] ), .B1(n36245), .B2(
        \REGISTERS[22][24] ), .ZN(n35764) );
  AOI22_X1 U375 ( .A1(n36260), .A2(\REGISTERS[15][24] ), .B1(n36258), .B2(
        \REGISTERS[9][24] ), .ZN(n35765) );
  NAND4_X1 U376 ( .A1(n35762), .A2(n35763), .A3(n35764), .A4(n35765), .ZN(
        n35766) );
  AOI22_X1 U377 ( .A1(n36262), .A2(\REGISTERS[16][24] ), .B1(n36263), .B2(
        \REGISTERS[25][24] ), .ZN(n35767) );
  AOI22_X1 U378 ( .A1(n36265), .A2(\REGISTERS[11][24] ), .B1(n36264), .B2(
        \REGISTERS[2][24] ), .ZN(n35768) );
  AOI22_X1 U379 ( .A1(n36267), .A2(\REGISTERS[31][24] ), .B1(n36261), .B2(
        \REGISTERS[13][24] ), .ZN(n35769) );
  AOI22_X1 U380 ( .A1(n36255), .A2(\REGISTERS[29][24] ), .B1(n36259), .B2(
        \REGISTERS[8][24] ), .ZN(n35770) );
  NAND4_X1 U381 ( .A1(n35767), .A2(n35768), .A3(n35769), .A4(n35770), .ZN(
        n35771) );
  AOI22_X1 U382 ( .A1(n36254), .A2(\REGISTERS[26][24] ), .B1(n36256), .B2(
        \REGISTERS[21][24] ), .ZN(n35772) );
  AOI22_X1 U383 ( .A1(n36251), .A2(\REGISTERS[1][24] ), .B1(n36252), .B2(
        \REGISTERS[7][24] ), .ZN(n35773) );
  AOI222_X1 U384 ( .A1(n36248), .A2(\REGISTERS[20][24] ), .B1(n36249), .B2(
        \REGISTERS[5][24] ), .C1(n36247), .C2(\REGISTERS[18][24] ), .ZN(n35774) );
  NAND3_X1 U385 ( .A1(n35772), .A2(n35773), .A3(n35774), .ZN(n35775) );
  AOI22_X1 U386 ( .A1(n36244), .A2(\REGISTERS[28][24] ), .B1(n36246), .B2(
        \REGISTERS[19][24] ), .ZN(n35776) );
  AOI22_X1 U387 ( .A1(n36243), .A2(\REGISTERS[6][24] ), .B1(n36257), .B2(
        \REGISTERS[23][24] ), .ZN(n35777) );
  AOI22_X1 U388 ( .A1(n36253), .A2(\REGISTERS[24][24] ), .B1(n36241), .B2(
        \REGISTERS[10][24] ), .ZN(n35778) );
  AOI22_X1 U389 ( .A1(n36239), .A2(\REGISTERS[12][24] ), .B1(n36266), .B2(
        \REGISTERS[27][24] ), .ZN(n35779) );
  NAND4_X1 U390 ( .A1(n35776), .A2(n35777), .A3(n35778), .A4(n35779), .ZN(
        n35780) );
  OR4_X1 U391 ( .A1(n35766), .A2(n35771), .A3(n35775), .A4(n35780), .ZN(
        OUTB[24]) );
  AOI22_X1 U392 ( .A1(n36240), .A2(\REGISTERS[30][23] ), .B1(n36237), .B2(
        \REGISTERS[14][23] ), .ZN(n35781) );
  AOI22_X1 U393 ( .A1(n36238), .A2(\REGISTERS[3][23] ), .B1(n36242), .B2(
        \REGISTERS[4][23] ), .ZN(n35782) );
  AOI22_X1 U394 ( .A1(n36250), .A2(\REGISTERS[17][23] ), .B1(n36245), .B2(
        \REGISTERS[22][23] ), .ZN(n35783) );
  AOI22_X1 U395 ( .A1(n36260), .A2(\REGISTERS[15][23] ), .B1(n36258), .B2(
        \REGISTERS[9][23] ), .ZN(n35784) );
  NAND4_X1 U396 ( .A1(n35781), .A2(n35782), .A3(n35783), .A4(n35784), .ZN(
        n35785) );
  AOI22_X1 U397 ( .A1(n36262), .A2(\REGISTERS[16][23] ), .B1(n36263), .B2(
        \REGISTERS[25][23] ), .ZN(n35786) );
  AOI22_X1 U398 ( .A1(n36265), .A2(\REGISTERS[11][23] ), .B1(n36264), .B2(
        \REGISTERS[2][23] ), .ZN(n35787) );
  AOI22_X1 U399 ( .A1(n36267), .A2(\REGISTERS[31][23] ), .B1(n36261), .B2(
        \REGISTERS[13][23] ), .ZN(n35788) );
  AOI22_X1 U400 ( .A1(n36255), .A2(\REGISTERS[29][23] ), .B1(n36259), .B2(
        \REGISTERS[8][23] ), .ZN(n35789) );
  NAND4_X1 U401 ( .A1(n35786), .A2(n35787), .A3(n35788), .A4(n35789), .ZN(
        n35790) );
  AOI22_X1 U402 ( .A1(n36254), .A2(\REGISTERS[26][23] ), .B1(n36256), .B2(
        \REGISTERS[21][23] ), .ZN(n35791) );
  AOI22_X1 U403 ( .A1(n36251), .A2(\REGISTERS[1][23] ), .B1(n36252), .B2(
        \REGISTERS[7][23] ), .ZN(n35792) );
  AOI222_X1 U404 ( .A1(n36248), .A2(\REGISTERS[20][23] ), .B1(n36249), .B2(
        \REGISTERS[5][23] ), .C1(n36247), .C2(\REGISTERS[18][23] ), .ZN(n35793) );
  NAND3_X1 U405 ( .A1(n35791), .A2(n35792), .A3(n35793), .ZN(n35794) );
  AOI22_X1 U406 ( .A1(n36244), .A2(\REGISTERS[28][23] ), .B1(n36246), .B2(
        \REGISTERS[19][23] ), .ZN(n35795) );
  AOI22_X1 U407 ( .A1(n36243), .A2(\REGISTERS[6][23] ), .B1(n36257), .B2(
        \REGISTERS[23][23] ), .ZN(n35796) );
  AOI22_X1 U408 ( .A1(n36253), .A2(\REGISTERS[24][23] ), .B1(n36241), .B2(
        \REGISTERS[10][23] ), .ZN(n35797) );
  AOI22_X1 U409 ( .A1(n36239), .A2(\REGISTERS[12][23] ), .B1(n36266), .B2(
        \REGISTERS[27][23] ), .ZN(n35798) );
  NAND4_X1 U410 ( .A1(n35795), .A2(n35796), .A3(n35797), .A4(n35798), .ZN(
        n35799) );
  OR4_X1 U411 ( .A1(n35785), .A2(n35790), .A3(n35794), .A4(n35799), .ZN(
        OUTB[23]) );
  AOI22_X1 U412 ( .A1(n36240), .A2(\REGISTERS[30][22] ), .B1(n36237), .B2(
        \REGISTERS[14][22] ), .ZN(n35800) );
  AOI22_X1 U413 ( .A1(n36238), .A2(\REGISTERS[3][22] ), .B1(n36242), .B2(
        \REGISTERS[4][22] ), .ZN(n35801) );
  AOI22_X1 U414 ( .A1(n36250), .A2(\REGISTERS[17][22] ), .B1(n36245), .B2(
        \REGISTERS[22][22] ), .ZN(n35802) );
  AOI22_X1 U415 ( .A1(n36260), .A2(\REGISTERS[15][22] ), .B1(n36258), .B2(
        \REGISTERS[9][22] ), .ZN(n35803) );
  NAND4_X1 U416 ( .A1(n35800), .A2(n35801), .A3(n35802), .A4(n35803), .ZN(
        n35804) );
  AOI22_X1 U417 ( .A1(n36262), .A2(\REGISTERS[16][22] ), .B1(n36263), .B2(
        \REGISTERS[25][22] ), .ZN(n35805) );
  AOI22_X1 U418 ( .A1(n36265), .A2(\REGISTERS[11][22] ), .B1(n36264), .B2(
        \REGISTERS[2][22] ), .ZN(n35806) );
  AOI22_X1 U419 ( .A1(n36267), .A2(\REGISTERS[31][22] ), .B1(n36261), .B2(
        \REGISTERS[13][22] ), .ZN(n35807) );
  AOI22_X1 U420 ( .A1(n36255), .A2(\REGISTERS[29][22] ), .B1(n36259), .B2(
        \REGISTERS[8][22] ), .ZN(n35808) );
  NAND4_X1 U421 ( .A1(n35805), .A2(n35806), .A3(n35807), .A4(n35808), .ZN(
        n35809) );
  AOI22_X1 U422 ( .A1(n36254), .A2(\REGISTERS[26][22] ), .B1(n36256), .B2(
        \REGISTERS[21][22] ), .ZN(n35810) );
  AOI22_X1 U423 ( .A1(n36251), .A2(\REGISTERS[1][22] ), .B1(n36252), .B2(
        \REGISTERS[7][22] ), .ZN(n35811) );
  AOI222_X1 U424 ( .A1(n36248), .A2(\REGISTERS[20][22] ), .B1(n36249), .B2(
        \REGISTERS[5][22] ), .C1(n36247), .C2(\REGISTERS[18][22] ), .ZN(n35812) );
  NAND3_X1 U425 ( .A1(n35810), .A2(n35811), .A3(n35812), .ZN(n35813) );
  AOI22_X1 U426 ( .A1(n36244), .A2(\REGISTERS[28][22] ), .B1(n36246), .B2(
        \REGISTERS[19][22] ), .ZN(n35814) );
  AOI22_X1 U427 ( .A1(n36243), .A2(\REGISTERS[6][22] ), .B1(n36257), .B2(
        \REGISTERS[23][22] ), .ZN(n35815) );
  AOI22_X1 U428 ( .A1(n36253), .A2(\REGISTERS[24][22] ), .B1(n36241), .B2(
        \REGISTERS[10][22] ), .ZN(n35816) );
  AOI22_X1 U429 ( .A1(n36239), .A2(\REGISTERS[12][22] ), .B1(n36266), .B2(
        \REGISTERS[27][22] ), .ZN(n35817) );
  NAND4_X1 U430 ( .A1(n35814), .A2(n35815), .A3(n35816), .A4(n35817), .ZN(
        n35818) );
  OR4_X1 U431 ( .A1(n35804), .A2(n35809), .A3(n35813), .A4(n35818), .ZN(
        OUTB[22]) );
  AOI22_X1 U432 ( .A1(n36240), .A2(\REGISTERS[30][21] ), .B1(n36237), .B2(
        \REGISTERS[14][21] ), .ZN(n35819) );
  AOI22_X1 U433 ( .A1(n36238), .A2(\REGISTERS[3][21] ), .B1(n36242), .B2(
        \REGISTERS[4][21] ), .ZN(n35820) );
  AOI22_X1 U434 ( .A1(n36250), .A2(\REGISTERS[17][21] ), .B1(n36245), .B2(
        \REGISTERS[22][21] ), .ZN(n35821) );
  AOI22_X1 U435 ( .A1(n36260), .A2(\REGISTERS[15][21] ), .B1(n36258), .B2(
        \REGISTERS[9][21] ), .ZN(n35822) );
  NAND4_X1 U436 ( .A1(n35819), .A2(n35820), .A3(n35821), .A4(n35822), .ZN(
        n35823) );
  AOI22_X1 U437 ( .A1(n36262), .A2(\REGISTERS[16][21] ), .B1(n36263), .B2(
        \REGISTERS[25][21] ), .ZN(n35824) );
  AOI22_X1 U438 ( .A1(n36265), .A2(\REGISTERS[11][21] ), .B1(n36264), .B2(
        \REGISTERS[2][21] ), .ZN(n35825) );
  AOI22_X1 U439 ( .A1(n36267), .A2(\REGISTERS[31][21] ), .B1(n36261), .B2(
        \REGISTERS[13][21] ), .ZN(n35826) );
  AOI22_X1 U440 ( .A1(n36255), .A2(\REGISTERS[29][21] ), .B1(n36259), .B2(
        \REGISTERS[8][21] ), .ZN(n35827) );
  NAND4_X1 U441 ( .A1(n35824), .A2(n35825), .A3(n35826), .A4(n35827), .ZN(
        n35828) );
  AOI22_X1 U442 ( .A1(n36254), .A2(\REGISTERS[26][21] ), .B1(n36256), .B2(
        \REGISTERS[21][21] ), .ZN(n35829) );
  AOI22_X1 U443 ( .A1(n36251), .A2(\REGISTERS[1][21] ), .B1(n36252), .B2(
        \REGISTERS[7][21] ), .ZN(n35830) );
  AOI222_X1 U444 ( .A1(n36248), .A2(\REGISTERS[20][21] ), .B1(n36249), .B2(
        \REGISTERS[5][21] ), .C1(n36247), .C2(\REGISTERS[18][21] ), .ZN(n35831) );
  NAND3_X1 U445 ( .A1(n35829), .A2(n35830), .A3(n35831), .ZN(n35832) );
  AOI22_X1 U446 ( .A1(n36244), .A2(\REGISTERS[28][21] ), .B1(n36246), .B2(
        \REGISTERS[19][21] ), .ZN(n35833) );
  AOI22_X1 U447 ( .A1(n36243), .A2(\REGISTERS[6][21] ), .B1(n36257), .B2(
        \REGISTERS[23][21] ), .ZN(n35834) );
  AOI22_X1 U448 ( .A1(n36253), .A2(\REGISTERS[24][21] ), .B1(n36241), .B2(
        \REGISTERS[10][21] ), .ZN(n35835) );
  AOI22_X1 U449 ( .A1(n36239), .A2(\REGISTERS[12][21] ), .B1(n36266), .B2(
        \REGISTERS[27][21] ), .ZN(n35836) );
  NAND4_X1 U450 ( .A1(n35833), .A2(n35834), .A3(n35835), .A4(n35836), .ZN(
        n35837) );
  OR4_X1 U451 ( .A1(n35823), .A2(n35828), .A3(n35832), .A4(n35837), .ZN(
        OUTB[21]) );
  AOI22_X1 U452 ( .A1(n36240), .A2(\REGISTERS[30][20] ), .B1(n36237), .B2(
        \REGISTERS[14][20] ), .ZN(n35838) );
  AOI22_X1 U453 ( .A1(n36238), .A2(\REGISTERS[3][20] ), .B1(n36242), .B2(
        \REGISTERS[4][20] ), .ZN(n35839) );
  AOI22_X1 U454 ( .A1(n36250), .A2(\REGISTERS[17][20] ), .B1(n36245), .B2(
        \REGISTERS[22][20] ), .ZN(n35840) );
  AOI22_X1 U455 ( .A1(n36260), .A2(\REGISTERS[15][20] ), .B1(n36258), .B2(
        \REGISTERS[9][20] ), .ZN(n35841) );
  NAND4_X1 U456 ( .A1(n35838), .A2(n35839), .A3(n35840), .A4(n35841), .ZN(
        n35842) );
  AOI22_X1 U457 ( .A1(n36262), .A2(\REGISTERS[16][20] ), .B1(n36263), .B2(
        \REGISTERS[25][20] ), .ZN(n35843) );
  AOI22_X1 U458 ( .A1(n36265), .A2(\REGISTERS[11][20] ), .B1(n36264), .B2(
        \REGISTERS[2][20] ), .ZN(n35844) );
  AOI22_X1 U459 ( .A1(n36267), .A2(\REGISTERS[31][20] ), .B1(n36261), .B2(
        \REGISTERS[13][20] ), .ZN(n35845) );
  AOI22_X1 U460 ( .A1(n36255), .A2(\REGISTERS[29][20] ), .B1(n36259), .B2(
        \REGISTERS[8][20] ), .ZN(n35846) );
  NAND4_X1 U461 ( .A1(n35843), .A2(n35844), .A3(n35845), .A4(n35846), .ZN(
        n35847) );
  AOI22_X1 U462 ( .A1(n36254), .A2(\REGISTERS[26][20] ), .B1(n36256), .B2(
        \REGISTERS[21][20] ), .ZN(n35848) );
  AOI22_X1 U463 ( .A1(n36251), .A2(\REGISTERS[1][20] ), .B1(n36252), .B2(
        \REGISTERS[7][20] ), .ZN(n35849) );
  AOI222_X1 U464 ( .A1(n36248), .A2(\REGISTERS[20][20] ), .B1(n36249), .B2(
        \REGISTERS[5][20] ), .C1(n36247), .C2(\REGISTERS[18][20] ), .ZN(n35850) );
  NAND3_X1 U465 ( .A1(n35848), .A2(n35849), .A3(n35850), .ZN(n35851) );
  AOI22_X1 U466 ( .A1(n36244), .A2(\REGISTERS[28][20] ), .B1(n36246), .B2(
        \REGISTERS[19][20] ), .ZN(n35852) );
  AOI22_X1 U467 ( .A1(n36243), .A2(\REGISTERS[6][20] ), .B1(n36257), .B2(
        \REGISTERS[23][20] ), .ZN(n35853) );
  AOI22_X1 U468 ( .A1(n36253), .A2(\REGISTERS[24][20] ), .B1(n36241), .B2(
        \REGISTERS[10][20] ), .ZN(n35854) );
  AOI22_X1 U469 ( .A1(n36239), .A2(\REGISTERS[12][20] ), .B1(n36266), .B2(
        \REGISTERS[27][20] ), .ZN(n35855) );
  NAND4_X1 U470 ( .A1(n35852), .A2(n35853), .A3(n35854), .A4(n35855), .ZN(
        n35856) );
  OR4_X1 U471 ( .A1(n35842), .A2(n35847), .A3(n35851), .A4(n35856), .ZN(
        OUTB[20]) );
  AOI22_X1 U472 ( .A1(n36240), .A2(\REGISTERS[30][19] ), .B1(n36237), .B2(
        \REGISTERS[14][19] ), .ZN(n35857) );
  AOI22_X1 U473 ( .A1(n36238), .A2(\REGISTERS[3][19] ), .B1(n36242), .B2(
        \REGISTERS[4][19] ), .ZN(n35858) );
  AOI22_X1 U474 ( .A1(n36250), .A2(\REGISTERS[17][19] ), .B1(n36245), .B2(
        \REGISTERS[22][19] ), .ZN(n35859) );
  AOI22_X1 U475 ( .A1(n36260), .A2(\REGISTERS[15][19] ), .B1(n36258), .B2(
        \REGISTERS[9][19] ), .ZN(n35860) );
  NAND4_X1 U476 ( .A1(n35857), .A2(n35858), .A3(n35859), .A4(n35860), .ZN(
        n35861) );
  AOI22_X1 U477 ( .A1(n36262), .A2(\REGISTERS[16][19] ), .B1(n36263), .B2(
        \REGISTERS[25][19] ), .ZN(n35862) );
  AOI22_X1 U478 ( .A1(n36265), .A2(\REGISTERS[11][19] ), .B1(n36264), .B2(
        \REGISTERS[2][19] ), .ZN(n35863) );
  AOI22_X1 U479 ( .A1(n36267), .A2(\REGISTERS[31][19] ), .B1(n36261), .B2(
        \REGISTERS[13][19] ), .ZN(n35864) );
  AOI22_X1 U480 ( .A1(n36255), .A2(\REGISTERS[29][19] ), .B1(n36259), .B2(
        \REGISTERS[8][19] ), .ZN(n35865) );
  NAND4_X1 U481 ( .A1(n35862), .A2(n35863), .A3(n35864), .A4(n35865), .ZN(
        n35866) );
  AOI22_X1 U482 ( .A1(n36254), .A2(\REGISTERS[26][19] ), .B1(n36256), .B2(
        \REGISTERS[21][19] ), .ZN(n35867) );
  AOI22_X1 U483 ( .A1(n36251), .A2(\REGISTERS[1][19] ), .B1(n36252), .B2(
        \REGISTERS[7][19] ), .ZN(n35868) );
  AOI222_X1 U484 ( .A1(n36248), .A2(\REGISTERS[20][19] ), .B1(n36249), .B2(
        \REGISTERS[5][19] ), .C1(n36247), .C2(\REGISTERS[18][19] ), .ZN(n35869) );
  NAND3_X1 U485 ( .A1(n35867), .A2(n35868), .A3(n35869), .ZN(n35870) );
  AOI22_X1 U486 ( .A1(n36244), .A2(\REGISTERS[28][19] ), .B1(n36246), .B2(
        \REGISTERS[19][19] ), .ZN(n35871) );
  AOI22_X1 U487 ( .A1(n36243), .A2(\REGISTERS[6][19] ), .B1(n36257), .B2(
        \REGISTERS[23][19] ), .ZN(n35872) );
  AOI22_X1 U488 ( .A1(n36253), .A2(\REGISTERS[24][19] ), .B1(n36241), .B2(
        \REGISTERS[10][19] ), .ZN(n35873) );
  AOI22_X1 U489 ( .A1(n36239), .A2(\REGISTERS[12][19] ), .B1(n36266), .B2(
        \REGISTERS[27][19] ), .ZN(n35874) );
  NAND4_X1 U490 ( .A1(n35871), .A2(n35872), .A3(n35873), .A4(n35874), .ZN(
        n35875) );
  OR4_X1 U491 ( .A1(n35861), .A2(n35866), .A3(n35870), .A4(n35875), .ZN(
        OUTB[19]) );
  AOI22_X1 U492 ( .A1(n36240), .A2(\REGISTERS[30][18] ), .B1(n36237), .B2(
        \REGISTERS[14][18] ), .ZN(n35876) );
  AOI22_X1 U493 ( .A1(n36238), .A2(\REGISTERS[3][18] ), .B1(n36242), .B2(
        \REGISTERS[4][18] ), .ZN(n35877) );
  AOI22_X1 U494 ( .A1(n36250), .A2(\REGISTERS[17][18] ), .B1(n36245), .B2(
        \REGISTERS[22][18] ), .ZN(n35878) );
  AOI22_X1 U495 ( .A1(n36260), .A2(\REGISTERS[15][18] ), .B1(n36258), .B2(
        \REGISTERS[9][18] ), .ZN(n35879) );
  NAND4_X1 U496 ( .A1(n35876), .A2(n35877), .A3(n35878), .A4(n35879), .ZN(
        n35880) );
  AOI22_X1 U497 ( .A1(n36262), .A2(\REGISTERS[16][18] ), .B1(n36263), .B2(
        \REGISTERS[25][18] ), .ZN(n35881) );
  AOI22_X1 U498 ( .A1(n36265), .A2(\REGISTERS[11][18] ), .B1(n36264), .B2(
        \REGISTERS[2][18] ), .ZN(n35882) );
  AOI22_X1 U499 ( .A1(n36267), .A2(\REGISTERS[31][18] ), .B1(n36261), .B2(
        \REGISTERS[13][18] ), .ZN(n35883) );
  AOI22_X1 U500 ( .A1(n36255), .A2(\REGISTERS[29][18] ), .B1(n36259), .B2(
        \REGISTERS[8][18] ), .ZN(n35884) );
  NAND4_X1 U501 ( .A1(n35881), .A2(n35882), .A3(n35883), .A4(n35884), .ZN(
        n35885) );
  AOI22_X1 U502 ( .A1(n36254), .A2(\REGISTERS[26][18] ), .B1(n36256), .B2(
        \REGISTERS[21][18] ), .ZN(n35886) );
  AOI22_X1 U503 ( .A1(n36251), .A2(\REGISTERS[1][18] ), .B1(n36252), .B2(
        \REGISTERS[7][18] ), .ZN(n35887) );
  AOI222_X1 U504 ( .A1(n36248), .A2(\REGISTERS[20][18] ), .B1(n36249), .B2(
        \REGISTERS[5][18] ), .C1(n36247), .C2(\REGISTERS[18][18] ), .ZN(n35888) );
  NAND3_X1 U505 ( .A1(n35886), .A2(n35887), .A3(n35888), .ZN(n35889) );
  AOI22_X1 U506 ( .A1(n36244), .A2(\REGISTERS[28][18] ), .B1(n36246), .B2(
        \REGISTERS[19][18] ), .ZN(n35890) );
  AOI22_X1 U507 ( .A1(n36243), .A2(\REGISTERS[6][18] ), .B1(n36257), .B2(
        \REGISTERS[23][18] ), .ZN(n35891) );
  AOI22_X1 U508 ( .A1(n36253), .A2(\REGISTERS[24][18] ), .B1(n36241), .B2(
        \REGISTERS[10][18] ), .ZN(n35892) );
  AOI22_X1 U509 ( .A1(n36239), .A2(\REGISTERS[12][18] ), .B1(n36266), .B2(
        \REGISTERS[27][18] ), .ZN(n35893) );
  NAND4_X1 U510 ( .A1(n35890), .A2(n35891), .A3(n35892), .A4(n35893), .ZN(
        n35894) );
  OR4_X1 U511 ( .A1(n35880), .A2(n35885), .A3(n35889), .A4(n35894), .ZN(
        OUTB[18]) );
  AOI22_X1 U512 ( .A1(n36240), .A2(\REGISTERS[30][17] ), .B1(n36237), .B2(
        \REGISTERS[14][17] ), .ZN(n35895) );
  AOI22_X1 U513 ( .A1(n36238), .A2(\REGISTERS[3][17] ), .B1(n36242), .B2(
        \REGISTERS[4][17] ), .ZN(n35896) );
  AOI22_X1 U514 ( .A1(n36250), .A2(\REGISTERS[17][17] ), .B1(n36245), .B2(
        \REGISTERS[22][17] ), .ZN(n35897) );
  AOI22_X1 U515 ( .A1(n36260), .A2(\REGISTERS[15][17] ), .B1(n36258), .B2(
        \REGISTERS[9][17] ), .ZN(n35898) );
  NAND4_X1 U516 ( .A1(n35895), .A2(n35896), .A3(n35897), .A4(n35898), .ZN(
        n35899) );
  AOI22_X1 U517 ( .A1(n36262), .A2(\REGISTERS[16][17] ), .B1(n36263), .B2(
        \REGISTERS[25][17] ), .ZN(n35900) );
  AOI22_X1 U518 ( .A1(n36265), .A2(\REGISTERS[11][17] ), .B1(n36264), .B2(
        \REGISTERS[2][17] ), .ZN(n35901) );
  AOI22_X1 U519 ( .A1(n36267), .A2(\REGISTERS[31][17] ), .B1(n36261), .B2(
        \REGISTERS[13][17] ), .ZN(n35902) );
  AOI22_X1 U520 ( .A1(n36255), .A2(\REGISTERS[29][17] ), .B1(n36259), .B2(
        \REGISTERS[8][17] ), .ZN(n35903) );
  NAND4_X1 U521 ( .A1(n35900), .A2(n35901), .A3(n35902), .A4(n35903), .ZN(
        n35904) );
  AOI22_X1 U522 ( .A1(n36254), .A2(\REGISTERS[26][17] ), .B1(n36256), .B2(
        \REGISTERS[21][17] ), .ZN(n35905) );
  AOI22_X1 U523 ( .A1(n36251), .A2(\REGISTERS[1][17] ), .B1(n36252), .B2(
        \REGISTERS[7][17] ), .ZN(n35906) );
  AOI222_X1 U524 ( .A1(n36248), .A2(\REGISTERS[20][17] ), .B1(n36249), .B2(
        \REGISTERS[5][17] ), .C1(n36247), .C2(\REGISTERS[18][17] ), .ZN(n35907) );
  NAND3_X1 U525 ( .A1(n35905), .A2(n35906), .A3(n35907), .ZN(n35908) );
  AOI22_X1 U526 ( .A1(n36244), .A2(\REGISTERS[28][17] ), .B1(n36246), .B2(
        \REGISTERS[19][17] ), .ZN(n35909) );
  AOI22_X1 U527 ( .A1(n36243), .A2(\REGISTERS[6][17] ), .B1(n36257), .B2(
        \REGISTERS[23][17] ), .ZN(n35910) );
  AOI22_X1 U528 ( .A1(n36253), .A2(\REGISTERS[24][17] ), .B1(n36241), .B2(
        \REGISTERS[10][17] ), .ZN(n35911) );
  AOI22_X1 U529 ( .A1(n36239), .A2(\REGISTERS[12][17] ), .B1(n36266), .B2(
        \REGISTERS[27][17] ), .ZN(n35912) );
  NAND4_X1 U530 ( .A1(n35909), .A2(n35910), .A3(n35911), .A4(n35912), .ZN(
        n35913) );
  OR4_X1 U531 ( .A1(n35899), .A2(n35904), .A3(n35908), .A4(n35913), .ZN(
        OUTB[17]) );
  AOI22_X1 U532 ( .A1(n36240), .A2(\REGISTERS[30][16] ), .B1(n36237), .B2(
        \REGISTERS[14][16] ), .ZN(n35914) );
  AOI22_X1 U533 ( .A1(n36238), .A2(\REGISTERS[3][16] ), .B1(n36242), .B2(
        \REGISTERS[4][16] ), .ZN(n35915) );
  AOI22_X1 U534 ( .A1(n36250), .A2(\REGISTERS[17][16] ), .B1(n36245), .B2(
        \REGISTERS[22][16] ), .ZN(n35916) );
  AOI22_X1 U535 ( .A1(n36260), .A2(\REGISTERS[15][16] ), .B1(n36258), .B2(
        \REGISTERS[9][16] ), .ZN(n35917) );
  NAND4_X1 U536 ( .A1(n35914), .A2(n35915), .A3(n35916), .A4(n35917), .ZN(
        n35918) );
  AOI22_X1 U537 ( .A1(n36262), .A2(\REGISTERS[16][16] ), .B1(n36263), .B2(
        \REGISTERS[25][16] ), .ZN(n35919) );
  AOI22_X1 U538 ( .A1(n36265), .A2(\REGISTERS[11][16] ), .B1(n36264), .B2(
        \REGISTERS[2][16] ), .ZN(n35920) );
  AOI22_X1 U539 ( .A1(n36267), .A2(\REGISTERS[31][16] ), .B1(n36261), .B2(
        \REGISTERS[13][16] ), .ZN(n35921) );
  AOI22_X1 U540 ( .A1(n36255), .A2(\REGISTERS[29][16] ), .B1(n36259), .B2(
        \REGISTERS[8][16] ), .ZN(n35922) );
  NAND4_X1 U541 ( .A1(n35919), .A2(n35920), .A3(n35921), .A4(n35922), .ZN(
        n35923) );
  AOI22_X1 U542 ( .A1(n36254), .A2(\REGISTERS[26][16] ), .B1(n36256), .B2(
        \REGISTERS[21][16] ), .ZN(n35924) );
  AOI22_X1 U543 ( .A1(n36251), .A2(\REGISTERS[1][16] ), .B1(n36252), .B2(
        \REGISTERS[7][16] ), .ZN(n35925) );
  AOI222_X1 U544 ( .A1(n36248), .A2(\REGISTERS[20][16] ), .B1(n36249), .B2(
        \REGISTERS[5][16] ), .C1(n36247), .C2(\REGISTERS[18][16] ), .ZN(n35926) );
  NAND3_X1 U545 ( .A1(n35924), .A2(n35925), .A3(n35926), .ZN(n35927) );
  AOI22_X1 U546 ( .A1(n36244), .A2(\REGISTERS[28][16] ), .B1(n36246), .B2(
        \REGISTERS[19][16] ), .ZN(n35928) );
  AOI22_X1 U547 ( .A1(n36243), .A2(\REGISTERS[6][16] ), .B1(n36257), .B2(
        \REGISTERS[23][16] ), .ZN(n35929) );
  AOI22_X1 U548 ( .A1(n36253), .A2(\REGISTERS[24][16] ), .B1(n36241), .B2(
        \REGISTERS[10][16] ), .ZN(n35930) );
  AOI22_X1 U549 ( .A1(n36239), .A2(\REGISTERS[12][16] ), .B1(n36266), .B2(
        \REGISTERS[27][16] ), .ZN(n35931) );
  NAND4_X1 U550 ( .A1(n35928), .A2(n35929), .A3(n35930), .A4(n35931), .ZN(
        n35932) );
  OR4_X1 U551 ( .A1(n35918), .A2(n35923), .A3(n35927), .A4(n35932), .ZN(
        OUTB[16]) );
  AOI22_X1 U552 ( .A1(n36240), .A2(\REGISTERS[30][15] ), .B1(n36237), .B2(
        \REGISTERS[14][15] ), .ZN(n35933) );
  AOI22_X1 U553 ( .A1(n36238), .A2(\REGISTERS[3][15] ), .B1(n36242), .B2(
        \REGISTERS[4][15] ), .ZN(n35934) );
  AOI22_X1 U554 ( .A1(n36250), .A2(\REGISTERS[17][15] ), .B1(n36245), .B2(
        \REGISTERS[22][15] ), .ZN(n35935) );
  AOI22_X1 U555 ( .A1(n36260), .A2(\REGISTERS[15][15] ), .B1(n36258), .B2(
        \REGISTERS[9][15] ), .ZN(n35936) );
  NAND4_X1 U556 ( .A1(n35933), .A2(n35934), .A3(n35935), .A4(n35936), .ZN(
        n35937) );
  AOI22_X1 U557 ( .A1(n36262), .A2(\REGISTERS[16][15] ), .B1(n36263), .B2(
        \REGISTERS[25][15] ), .ZN(n35938) );
  AOI22_X1 U558 ( .A1(n36265), .A2(\REGISTERS[11][15] ), .B1(n36264), .B2(
        \REGISTERS[2][15] ), .ZN(n35939) );
  AOI22_X1 U559 ( .A1(n36267), .A2(\REGISTERS[31][15] ), .B1(n36261), .B2(
        \REGISTERS[13][15] ), .ZN(n35940) );
  AOI22_X1 U560 ( .A1(n36255), .A2(\REGISTERS[29][15] ), .B1(n36259), .B2(
        \REGISTERS[8][15] ), .ZN(n35941) );
  NAND4_X1 U561 ( .A1(n35938), .A2(n35939), .A3(n35940), .A4(n35941), .ZN(
        n35942) );
  AOI22_X1 U562 ( .A1(n36254), .A2(\REGISTERS[26][15] ), .B1(n36256), .B2(
        \REGISTERS[21][15] ), .ZN(n35943) );
  AOI22_X1 U563 ( .A1(n36251), .A2(\REGISTERS[1][15] ), .B1(n36252), .B2(
        \REGISTERS[7][15] ), .ZN(n35944) );
  AOI222_X1 U564 ( .A1(n36248), .A2(\REGISTERS[20][15] ), .B1(n36249), .B2(
        \REGISTERS[5][15] ), .C1(n36247), .C2(\REGISTERS[18][15] ), .ZN(n35945) );
  NAND3_X1 U565 ( .A1(n35943), .A2(n35944), .A3(n35945), .ZN(n35946) );
  AOI22_X1 U566 ( .A1(n36244), .A2(\REGISTERS[28][15] ), .B1(n36246), .B2(
        \REGISTERS[19][15] ), .ZN(n35947) );
  AOI22_X1 U567 ( .A1(n36243), .A2(\REGISTERS[6][15] ), .B1(n36257), .B2(
        \REGISTERS[23][15] ), .ZN(n35948) );
  AOI22_X1 U568 ( .A1(n36253), .A2(\REGISTERS[24][15] ), .B1(n36241), .B2(
        \REGISTERS[10][15] ), .ZN(n35949) );
  AOI22_X1 U569 ( .A1(n36239), .A2(\REGISTERS[12][15] ), .B1(n36266), .B2(
        \REGISTERS[27][15] ), .ZN(n35950) );
  NAND4_X1 U570 ( .A1(n35947), .A2(n35948), .A3(n35949), .A4(n35950), .ZN(
        n35951) );
  OR4_X1 U571 ( .A1(n35937), .A2(n35942), .A3(n35946), .A4(n35951), .ZN(
        OUTB[15]) );
  AOI22_X1 U572 ( .A1(n36240), .A2(\REGISTERS[30][14] ), .B1(n36237), .B2(
        \REGISTERS[14][14] ), .ZN(n35952) );
  AOI22_X1 U573 ( .A1(n36238), .A2(\REGISTERS[3][14] ), .B1(n36242), .B2(
        \REGISTERS[4][14] ), .ZN(n35953) );
  AOI22_X1 U574 ( .A1(n36250), .A2(\REGISTERS[17][14] ), .B1(n36245), .B2(
        \REGISTERS[22][14] ), .ZN(n35954) );
  AOI22_X1 U575 ( .A1(n36260), .A2(\REGISTERS[15][14] ), .B1(n36258), .B2(
        \REGISTERS[9][14] ), .ZN(n35955) );
  NAND4_X1 U576 ( .A1(n35952), .A2(n35953), .A3(n35954), .A4(n35955), .ZN(
        n35956) );
  AOI22_X1 U577 ( .A1(n36262), .A2(\REGISTERS[16][14] ), .B1(n36263), .B2(
        \REGISTERS[25][14] ), .ZN(n35957) );
  AOI22_X1 U578 ( .A1(n36265), .A2(\REGISTERS[11][14] ), .B1(n36264), .B2(
        \REGISTERS[2][14] ), .ZN(n35958) );
  AOI22_X1 U579 ( .A1(n36267), .A2(\REGISTERS[31][14] ), .B1(n36261), .B2(
        \REGISTERS[13][14] ), .ZN(n35959) );
  AOI22_X1 U580 ( .A1(n36255), .A2(\REGISTERS[29][14] ), .B1(n36259), .B2(
        \REGISTERS[8][14] ), .ZN(n35960) );
  NAND4_X1 U581 ( .A1(n35957), .A2(n35958), .A3(n35959), .A4(n35960), .ZN(
        n35961) );
  AOI22_X1 U582 ( .A1(n36254), .A2(\REGISTERS[26][14] ), .B1(n36256), .B2(
        \REGISTERS[21][14] ), .ZN(n35962) );
  AOI22_X1 U583 ( .A1(n36251), .A2(\REGISTERS[1][14] ), .B1(n36252), .B2(
        \REGISTERS[7][14] ), .ZN(n35963) );
  AOI222_X1 U584 ( .A1(n36248), .A2(\REGISTERS[20][14] ), .B1(n36249), .B2(
        \REGISTERS[5][14] ), .C1(n36247), .C2(\REGISTERS[18][14] ), .ZN(n35964) );
  NAND3_X1 U585 ( .A1(n35962), .A2(n35963), .A3(n35964), .ZN(n35965) );
  AOI22_X1 U586 ( .A1(n36244), .A2(\REGISTERS[28][14] ), .B1(n36246), .B2(
        \REGISTERS[19][14] ), .ZN(n35966) );
  AOI22_X1 U587 ( .A1(n36243), .A2(\REGISTERS[6][14] ), .B1(n36257), .B2(
        \REGISTERS[23][14] ), .ZN(n35967) );
  AOI22_X1 U588 ( .A1(n36253), .A2(\REGISTERS[24][14] ), .B1(n36241), .B2(
        \REGISTERS[10][14] ), .ZN(n35968) );
  AOI22_X1 U589 ( .A1(n36239), .A2(\REGISTERS[12][14] ), .B1(n36266), .B2(
        \REGISTERS[27][14] ), .ZN(n35969) );
  NAND4_X1 U590 ( .A1(n35966), .A2(n35967), .A3(n35968), .A4(n35969), .ZN(
        n35970) );
  OR4_X1 U591 ( .A1(n35956), .A2(n35961), .A3(n35965), .A4(n35970), .ZN(
        OUTB[14]) );
  AOI22_X1 U592 ( .A1(n36240), .A2(\REGISTERS[30][13] ), .B1(n36237), .B2(
        \REGISTERS[14][13] ), .ZN(n35971) );
  AOI22_X1 U593 ( .A1(n36238), .A2(\REGISTERS[3][13] ), .B1(n36242), .B2(
        \REGISTERS[4][13] ), .ZN(n35972) );
  AOI22_X1 U594 ( .A1(n36250), .A2(\REGISTERS[17][13] ), .B1(n36245), .B2(
        \REGISTERS[22][13] ), .ZN(n35973) );
  AOI22_X1 U595 ( .A1(n36260), .A2(\REGISTERS[15][13] ), .B1(n36258), .B2(
        \REGISTERS[9][13] ), .ZN(n35974) );
  NAND4_X1 U596 ( .A1(n35971), .A2(n35972), .A3(n35973), .A4(n35974), .ZN(
        n35975) );
  AOI22_X1 U597 ( .A1(n36262), .A2(\REGISTERS[16][13] ), .B1(n36263), .B2(
        \REGISTERS[25][13] ), .ZN(n35976) );
  AOI22_X1 U598 ( .A1(n36265), .A2(\REGISTERS[11][13] ), .B1(n36264), .B2(
        \REGISTERS[2][13] ), .ZN(n35977) );
  AOI22_X1 U599 ( .A1(n36267), .A2(\REGISTERS[31][13] ), .B1(n36261), .B2(
        \REGISTERS[13][13] ), .ZN(n35978) );
  AOI22_X1 U600 ( .A1(n36255), .A2(\REGISTERS[29][13] ), .B1(n36259), .B2(
        \REGISTERS[8][13] ), .ZN(n35979) );
  NAND4_X1 U601 ( .A1(n35976), .A2(n35977), .A3(n35978), .A4(n35979), .ZN(
        n35980) );
  AOI22_X1 U602 ( .A1(n36254), .A2(\REGISTERS[26][13] ), .B1(n36256), .B2(
        \REGISTERS[21][13] ), .ZN(n35981) );
  AOI22_X1 U603 ( .A1(n36251), .A2(\REGISTERS[1][13] ), .B1(n36252), .B2(
        \REGISTERS[7][13] ), .ZN(n35982) );
  AOI222_X1 U604 ( .A1(n36248), .A2(\REGISTERS[20][13] ), .B1(n36249), .B2(
        \REGISTERS[5][13] ), .C1(n36247), .C2(\REGISTERS[18][13] ), .ZN(n35983) );
  NAND3_X1 U605 ( .A1(n35981), .A2(n35982), .A3(n35983), .ZN(n35984) );
  AOI22_X1 U606 ( .A1(n36244), .A2(\REGISTERS[28][13] ), .B1(n36246), .B2(
        \REGISTERS[19][13] ), .ZN(n35985) );
  AOI22_X1 U607 ( .A1(n36243), .A2(\REGISTERS[6][13] ), .B1(n36257), .B2(
        \REGISTERS[23][13] ), .ZN(n35986) );
  AOI22_X1 U608 ( .A1(n36253), .A2(\REGISTERS[24][13] ), .B1(n36241), .B2(
        \REGISTERS[10][13] ), .ZN(n35987) );
  AOI22_X1 U609 ( .A1(n36239), .A2(\REGISTERS[12][13] ), .B1(n36266), .B2(
        \REGISTERS[27][13] ), .ZN(n35988) );
  NAND4_X1 U610 ( .A1(n35985), .A2(n35986), .A3(n35987), .A4(n35988), .ZN(
        n35989) );
  OR4_X1 U611 ( .A1(n35975), .A2(n35980), .A3(n35984), .A4(n35989), .ZN(
        OUTB[13]) );
  AOI22_X1 U612 ( .A1(n36240), .A2(\REGISTERS[30][12] ), .B1(n36237), .B2(
        \REGISTERS[14][12] ), .ZN(n35990) );
  AOI22_X1 U613 ( .A1(n36238), .A2(\REGISTERS[3][12] ), .B1(n36242), .B2(
        \REGISTERS[4][12] ), .ZN(n35991) );
  AOI22_X1 U614 ( .A1(n36250), .A2(\REGISTERS[17][12] ), .B1(n36245), .B2(
        \REGISTERS[22][12] ), .ZN(n35992) );
  AOI22_X1 U615 ( .A1(n36260), .A2(\REGISTERS[15][12] ), .B1(n36258), .B2(
        \REGISTERS[9][12] ), .ZN(n35993) );
  NAND4_X1 U616 ( .A1(n35990), .A2(n35991), .A3(n35992), .A4(n35993), .ZN(
        n35994) );
  AOI22_X1 U617 ( .A1(n36262), .A2(\REGISTERS[16][12] ), .B1(n36263), .B2(
        \REGISTERS[25][12] ), .ZN(n35995) );
  AOI22_X1 U618 ( .A1(n36265), .A2(\REGISTERS[11][12] ), .B1(n36264), .B2(
        \REGISTERS[2][12] ), .ZN(n35996) );
  AOI22_X1 U619 ( .A1(n36267), .A2(\REGISTERS[31][12] ), .B1(n36261), .B2(
        \REGISTERS[13][12] ), .ZN(n35997) );
  AOI22_X1 U620 ( .A1(n36255), .A2(\REGISTERS[29][12] ), .B1(n36259), .B2(
        \REGISTERS[8][12] ), .ZN(n35998) );
  NAND4_X1 U621 ( .A1(n35995), .A2(n35996), .A3(n35997), .A4(n35998), .ZN(
        n35999) );
  AOI22_X1 U622 ( .A1(n36254), .A2(\REGISTERS[26][12] ), .B1(n36256), .B2(
        \REGISTERS[21][12] ), .ZN(n36000) );
  AOI22_X1 U623 ( .A1(n36251), .A2(\REGISTERS[1][12] ), .B1(n36252), .B2(
        \REGISTERS[7][12] ), .ZN(n36001) );
  AOI222_X1 U624 ( .A1(n36248), .A2(\REGISTERS[20][12] ), .B1(n36249), .B2(
        \REGISTERS[5][12] ), .C1(n36247), .C2(\REGISTERS[18][12] ), .ZN(n36002) );
  NAND3_X1 U625 ( .A1(n36000), .A2(n36001), .A3(n36002), .ZN(n36003) );
  AOI22_X1 U626 ( .A1(n36244), .A2(\REGISTERS[28][12] ), .B1(n36246), .B2(
        \REGISTERS[19][12] ), .ZN(n36004) );
  AOI22_X1 U627 ( .A1(n36243), .A2(\REGISTERS[6][12] ), .B1(n36257), .B2(
        \REGISTERS[23][12] ), .ZN(n36005) );
  AOI22_X1 U628 ( .A1(n36253), .A2(\REGISTERS[24][12] ), .B1(n36241), .B2(
        \REGISTERS[10][12] ), .ZN(n36006) );
  AOI22_X1 U629 ( .A1(n36239), .A2(\REGISTERS[12][12] ), .B1(n36266), .B2(
        \REGISTERS[27][12] ), .ZN(n36007) );
  NAND4_X1 U630 ( .A1(n36004), .A2(n36005), .A3(n36006), .A4(n36007), .ZN(
        n36008) );
  OR4_X1 U631 ( .A1(n35994), .A2(n35999), .A3(n36003), .A4(n36008), .ZN(
        OUTB[12]) );
  AOI22_X1 U632 ( .A1(n36240), .A2(\REGISTERS[30][11] ), .B1(n36237), .B2(
        \REGISTERS[14][11] ), .ZN(n36009) );
  AOI22_X1 U633 ( .A1(n36238), .A2(\REGISTERS[3][11] ), .B1(n36242), .B2(
        \REGISTERS[4][11] ), .ZN(n36010) );
  AOI22_X1 U634 ( .A1(n36250), .A2(\REGISTERS[17][11] ), .B1(n36245), .B2(
        \REGISTERS[22][11] ), .ZN(n36011) );
  AOI22_X1 U635 ( .A1(n36260), .A2(\REGISTERS[15][11] ), .B1(n36258), .B2(
        \REGISTERS[9][11] ), .ZN(n36012) );
  NAND4_X1 U636 ( .A1(n36009), .A2(n36010), .A3(n36011), .A4(n36012), .ZN(
        n36013) );
  AOI22_X1 U637 ( .A1(n36262), .A2(\REGISTERS[16][11] ), .B1(n36263), .B2(
        \REGISTERS[25][11] ), .ZN(n36014) );
  AOI22_X1 U638 ( .A1(n36265), .A2(\REGISTERS[11][11] ), .B1(n36264), .B2(
        \REGISTERS[2][11] ), .ZN(n36015) );
  AOI22_X1 U639 ( .A1(n36267), .A2(\REGISTERS[31][11] ), .B1(n36261), .B2(
        \REGISTERS[13][11] ), .ZN(n36016) );
  AOI22_X1 U640 ( .A1(n36255), .A2(\REGISTERS[29][11] ), .B1(n36259), .B2(
        \REGISTERS[8][11] ), .ZN(n36017) );
  NAND4_X1 U641 ( .A1(n36014), .A2(n36015), .A3(n36016), .A4(n36017), .ZN(
        n36018) );
  AOI22_X1 U642 ( .A1(n36254), .A2(\REGISTERS[26][11] ), .B1(n36256), .B2(
        \REGISTERS[21][11] ), .ZN(n36019) );
  AOI22_X1 U643 ( .A1(n36251), .A2(\REGISTERS[1][11] ), .B1(n36252), .B2(
        \REGISTERS[7][11] ), .ZN(n36020) );
  AOI222_X1 U644 ( .A1(n36248), .A2(\REGISTERS[20][11] ), .B1(n36249), .B2(
        \REGISTERS[5][11] ), .C1(n36247), .C2(\REGISTERS[18][11] ), .ZN(n36021) );
  NAND3_X1 U645 ( .A1(n36019), .A2(n36020), .A3(n36021), .ZN(n36022) );
  AOI22_X1 U646 ( .A1(n36244), .A2(\REGISTERS[28][11] ), .B1(n36246), .B2(
        \REGISTERS[19][11] ), .ZN(n36023) );
  AOI22_X1 U647 ( .A1(n36243), .A2(\REGISTERS[6][11] ), .B1(n36257), .B2(
        \REGISTERS[23][11] ), .ZN(n36024) );
  AOI22_X1 U648 ( .A1(n36253), .A2(\REGISTERS[24][11] ), .B1(n36241), .B2(
        \REGISTERS[10][11] ), .ZN(n36025) );
  AOI22_X1 U649 ( .A1(n36239), .A2(\REGISTERS[12][11] ), .B1(n36266), .B2(
        \REGISTERS[27][11] ), .ZN(n36026) );
  NAND4_X1 U650 ( .A1(n36023), .A2(n36024), .A3(n36025), .A4(n36026), .ZN(
        n36027) );
  OR4_X1 U651 ( .A1(n36013), .A2(n36018), .A3(n36022), .A4(n36027), .ZN(
        OUTB[11]) );
  AOI22_X1 U652 ( .A1(n36240), .A2(\REGISTERS[30][10] ), .B1(n36237), .B2(
        \REGISTERS[14][10] ), .ZN(n36028) );
  AOI22_X1 U653 ( .A1(n36238), .A2(\REGISTERS[3][10] ), .B1(n36242), .B2(
        \REGISTERS[4][10] ), .ZN(n36029) );
  AOI22_X1 U654 ( .A1(n36250), .A2(\REGISTERS[17][10] ), .B1(n36245), .B2(
        \REGISTERS[22][10] ), .ZN(n36030) );
  AOI22_X1 U655 ( .A1(n36260), .A2(\REGISTERS[15][10] ), .B1(n36258), .B2(
        \REGISTERS[9][10] ), .ZN(n36031) );
  NAND4_X1 U656 ( .A1(n36028), .A2(n36029), .A3(n36030), .A4(n36031), .ZN(
        n36032) );
  AOI22_X1 U657 ( .A1(n36262), .A2(\REGISTERS[16][10] ), .B1(n36263), .B2(
        \REGISTERS[25][10] ), .ZN(n36033) );
  AOI22_X1 U658 ( .A1(n36265), .A2(\REGISTERS[11][10] ), .B1(n36264), .B2(
        \REGISTERS[2][10] ), .ZN(n36034) );
  AOI22_X1 U659 ( .A1(n36267), .A2(\REGISTERS[31][10] ), .B1(n36261), .B2(
        \REGISTERS[13][10] ), .ZN(n36035) );
  AOI22_X1 U660 ( .A1(n36255), .A2(\REGISTERS[29][10] ), .B1(n36259), .B2(
        \REGISTERS[8][10] ), .ZN(n36036) );
  NAND4_X1 U661 ( .A1(n36033), .A2(n36034), .A3(n36035), .A4(n36036), .ZN(
        n36037) );
  AOI22_X1 U662 ( .A1(n36254), .A2(\REGISTERS[26][10] ), .B1(n36256), .B2(
        \REGISTERS[21][10] ), .ZN(n36038) );
  AOI22_X1 U663 ( .A1(n36251), .A2(\REGISTERS[1][10] ), .B1(n36252), .B2(
        \REGISTERS[7][10] ), .ZN(n36039) );
  AOI222_X1 U664 ( .A1(n36248), .A2(\REGISTERS[20][10] ), .B1(n36249), .B2(
        \REGISTERS[5][10] ), .C1(n36247), .C2(\REGISTERS[18][10] ), .ZN(n36040) );
  NAND3_X1 U665 ( .A1(n36038), .A2(n36039), .A3(n36040), .ZN(n36041) );
  AOI22_X1 U666 ( .A1(n36244), .A2(\REGISTERS[28][10] ), .B1(n36246), .B2(
        \REGISTERS[19][10] ), .ZN(n36042) );
  AOI22_X1 U667 ( .A1(n36243), .A2(\REGISTERS[6][10] ), .B1(n36257), .B2(
        \REGISTERS[23][10] ), .ZN(n36043) );
  AOI22_X1 U668 ( .A1(n36253), .A2(\REGISTERS[24][10] ), .B1(n36241), .B2(
        \REGISTERS[10][10] ), .ZN(n36044) );
  AOI22_X1 U669 ( .A1(n36239), .A2(\REGISTERS[12][10] ), .B1(n36266), .B2(
        \REGISTERS[27][10] ), .ZN(n36045) );
  NAND4_X1 U670 ( .A1(n36042), .A2(n36043), .A3(n36044), .A4(n36045), .ZN(
        n36046) );
  OR4_X1 U671 ( .A1(n36032), .A2(n36037), .A3(n36041), .A4(n36046), .ZN(
        OUTB[10]) );
  AOI22_X1 U672 ( .A1(n36240), .A2(\REGISTERS[30][9] ), .B1(n36237), .B2(
        \REGISTERS[14][9] ), .ZN(n36047) );
  AOI22_X1 U673 ( .A1(n36238), .A2(\REGISTERS[3][9] ), .B1(n36242), .B2(
        \REGISTERS[4][9] ), .ZN(n36048) );
  AOI22_X1 U674 ( .A1(n36250), .A2(\REGISTERS[17][9] ), .B1(n36245), .B2(
        \REGISTERS[22][9] ), .ZN(n36049) );
  AOI22_X1 U675 ( .A1(n36260), .A2(\REGISTERS[15][9] ), .B1(n36258), .B2(
        \REGISTERS[9][9] ), .ZN(n36050) );
  NAND4_X1 U676 ( .A1(n36047), .A2(n36048), .A3(n36049), .A4(n36050), .ZN(
        n36051) );
  AOI22_X1 U677 ( .A1(n36262), .A2(\REGISTERS[16][9] ), .B1(n36263), .B2(
        \REGISTERS[25][9] ), .ZN(n36052) );
  AOI22_X1 U678 ( .A1(n36265), .A2(\REGISTERS[11][9] ), .B1(n36264), .B2(
        \REGISTERS[2][9] ), .ZN(n36053) );
  AOI22_X1 U679 ( .A1(n36267), .A2(\REGISTERS[31][9] ), .B1(n36261), .B2(
        \REGISTERS[13][9] ), .ZN(n36054) );
  AOI22_X1 U680 ( .A1(n36255), .A2(\REGISTERS[29][9] ), .B1(n36259), .B2(
        \REGISTERS[8][9] ), .ZN(n36055) );
  NAND4_X1 U681 ( .A1(n36052), .A2(n36053), .A3(n36054), .A4(n36055), .ZN(
        n36056) );
  AOI22_X1 U682 ( .A1(n36254), .A2(\REGISTERS[26][9] ), .B1(n36256), .B2(
        \REGISTERS[21][9] ), .ZN(n36057) );
  AOI22_X1 U683 ( .A1(n36251), .A2(\REGISTERS[1][9] ), .B1(n36252), .B2(
        \REGISTERS[7][9] ), .ZN(n36058) );
  AOI222_X1 U684 ( .A1(n36248), .A2(\REGISTERS[20][9] ), .B1(n36249), .B2(
        \REGISTERS[5][9] ), .C1(n36247), .C2(\REGISTERS[18][9] ), .ZN(n36059)
         );
  NAND3_X1 U685 ( .A1(n36057), .A2(n36058), .A3(n36059), .ZN(n36060) );
  AOI22_X1 U686 ( .A1(n36244), .A2(\REGISTERS[28][9] ), .B1(n36246), .B2(
        \REGISTERS[19][9] ), .ZN(n36061) );
  AOI22_X1 U687 ( .A1(n36243), .A2(\REGISTERS[6][9] ), .B1(n36257), .B2(
        \REGISTERS[23][9] ), .ZN(n36062) );
  AOI22_X1 U688 ( .A1(n36253), .A2(\REGISTERS[24][9] ), .B1(n36241), .B2(
        \REGISTERS[10][9] ), .ZN(n36063) );
  AOI22_X1 U689 ( .A1(n36239), .A2(\REGISTERS[12][9] ), .B1(n36266), .B2(
        \REGISTERS[27][9] ), .ZN(n36064) );
  NAND4_X1 U690 ( .A1(n36061), .A2(n36062), .A3(n36063), .A4(n36064), .ZN(
        n36065) );
  OR4_X1 U691 ( .A1(n36051), .A2(n36056), .A3(n36060), .A4(n36065), .ZN(
        OUTB[9]) );
  AOI22_X1 U692 ( .A1(n36240), .A2(\REGISTERS[30][8] ), .B1(n36237), .B2(
        \REGISTERS[14][8] ), .ZN(n36066) );
  AOI22_X1 U693 ( .A1(n36238), .A2(\REGISTERS[3][8] ), .B1(n36242), .B2(
        \REGISTERS[4][8] ), .ZN(n36067) );
  AOI22_X1 U694 ( .A1(n36250), .A2(\REGISTERS[17][8] ), .B1(n36245), .B2(
        \REGISTERS[22][8] ), .ZN(n36068) );
  AOI22_X1 U695 ( .A1(n36260), .A2(\REGISTERS[15][8] ), .B1(n36258), .B2(
        \REGISTERS[9][8] ), .ZN(n36069) );
  NAND4_X1 U696 ( .A1(n36066), .A2(n36067), .A3(n36068), .A4(n36069), .ZN(
        n36070) );
  AOI22_X1 U697 ( .A1(n36262), .A2(\REGISTERS[16][8] ), .B1(n36263), .B2(
        \REGISTERS[25][8] ), .ZN(n36071) );
  AOI22_X1 U698 ( .A1(n36265), .A2(\REGISTERS[11][8] ), .B1(n36264), .B2(
        \REGISTERS[2][8] ), .ZN(n36072) );
  AOI22_X1 U699 ( .A1(n36267), .A2(\REGISTERS[31][8] ), .B1(n36261), .B2(
        \REGISTERS[13][8] ), .ZN(n36073) );
  AOI22_X1 U700 ( .A1(n36255), .A2(\REGISTERS[29][8] ), .B1(n36259), .B2(
        \REGISTERS[8][8] ), .ZN(n36074) );
  NAND4_X1 U701 ( .A1(n36071), .A2(n36072), .A3(n36073), .A4(n36074), .ZN(
        n36075) );
  AOI22_X1 U702 ( .A1(n36254), .A2(\REGISTERS[26][8] ), .B1(n36256), .B2(
        \REGISTERS[21][8] ), .ZN(n36076) );
  AOI22_X1 U703 ( .A1(n36251), .A2(\REGISTERS[1][8] ), .B1(n36252), .B2(
        \REGISTERS[7][8] ), .ZN(n36077) );
  AOI222_X1 U704 ( .A1(n36248), .A2(\REGISTERS[20][8] ), .B1(n36249), .B2(
        \REGISTERS[5][8] ), .C1(n36247), .C2(\REGISTERS[18][8] ), .ZN(n36078)
         );
  NAND3_X1 U705 ( .A1(n36076), .A2(n36077), .A3(n36078), .ZN(n36079) );
  AOI22_X1 U706 ( .A1(n36244), .A2(\REGISTERS[28][8] ), .B1(n36246), .B2(
        \REGISTERS[19][8] ), .ZN(n36080) );
  AOI22_X1 U707 ( .A1(n36243), .A2(\REGISTERS[6][8] ), .B1(n36257), .B2(
        \REGISTERS[23][8] ), .ZN(n36081) );
  AOI22_X1 U708 ( .A1(n36253), .A2(\REGISTERS[24][8] ), .B1(n36241), .B2(
        \REGISTERS[10][8] ), .ZN(n36082) );
  AOI22_X1 U709 ( .A1(n36239), .A2(\REGISTERS[12][8] ), .B1(n36266), .B2(
        \REGISTERS[27][8] ), .ZN(n36083) );
  NAND4_X1 U710 ( .A1(n36080), .A2(n36081), .A3(n36082), .A4(n36083), .ZN(
        n36084) );
  OR4_X1 U711 ( .A1(n36070), .A2(n36075), .A3(n36079), .A4(n36084), .ZN(
        OUTB[8]) );
  AOI22_X1 U712 ( .A1(n36240), .A2(\REGISTERS[30][7] ), .B1(n36237), .B2(
        \REGISTERS[14][7] ), .ZN(n36085) );
  AOI22_X1 U713 ( .A1(n36238), .A2(\REGISTERS[3][7] ), .B1(n36242), .B2(
        \REGISTERS[4][7] ), .ZN(n36086) );
  AOI22_X1 U714 ( .A1(n36250), .A2(\REGISTERS[17][7] ), .B1(n36245), .B2(
        \REGISTERS[22][7] ), .ZN(n36087) );
  AOI22_X1 U715 ( .A1(n36260), .A2(\REGISTERS[15][7] ), .B1(n36258), .B2(
        \REGISTERS[9][7] ), .ZN(n36088) );
  NAND4_X1 U716 ( .A1(n36085), .A2(n36086), .A3(n36087), .A4(n36088), .ZN(
        n36089) );
  AOI22_X1 U717 ( .A1(n36262), .A2(\REGISTERS[16][7] ), .B1(n36263), .B2(
        \REGISTERS[25][7] ), .ZN(n36090) );
  AOI22_X1 U718 ( .A1(n36265), .A2(\REGISTERS[11][7] ), .B1(n36264), .B2(
        \REGISTERS[2][7] ), .ZN(n36091) );
  AOI22_X1 U719 ( .A1(n36267), .A2(\REGISTERS[31][7] ), .B1(n36261), .B2(
        \REGISTERS[13][7] ), .ZN(n36092) );
  AOI22_X1 U720 ( .A1(n36255), .A2(\REGISTERS[29][7] ), .B1(n36259), .B2(
        \REGISTERS[8][7] ), .ZN(n36093) );
  NAND4_X1 U721 ( .A1(n36090), .A2(n36091), .A3(n36092), .A4(n36093), .ZN(
        n36094) );
  AOI22_X1 U722 ( .A1(n36254), .A2(\REGISTERS[26][7] ), .B1(n36256), .B2(
        \REGISTERS[21][7] ), .ZN(n36095) );
  AOI22_X1 U723 ( .A1(n36251), .A2(\REGISTERS[1][7] ), .B1(n36252), .B2(
        \REGISTERS[7][7] ), .ZN(n36096) );
  AOI222_X1 U724 ( .A1(n36248), .A2(\REGISTERS[20][7] ), .B1(n36249), .B2(
        \REGISTERS[5][7] ), .C1(n36247), .C2(\REGISTERS[18][7] ), .ZN(n36097)
         );
  NAND3_X1 U725 ( .A1(n36095), .A2(n36096), .A3(n36097), .ZN(n36098) );
  AOI22_X1 U726 ( .A1(n36244), .A2(\REGISTERS[28][7] ), .B1(n36246), .B2(
        \REGISTERS[19][7] ), .ZN(n36099) );
  AOI22_X1 U727 ( .A1(n36243), .A2(\REGISTERS[6][7] ), .B1(n36257), .B2(
        \REGISTERS[23][7] ), .ZN(n36100) );
  AOI22_X1 U728 ( .A1(n36253), .A2(\REGISTERS[24][7] ), .B1(n36241), .B2(
        \REGISTERS[10][7] ), .ZN(n36101) );
  AOI22_X1 U729 ( .A1(n36239), .A2(\REGISTERS[12][7] ), .B1(n36266), .B2(
        \REGISTERS[27][7] ), .ZN(n36102) );
  NAND4_X1 U730 ( .A1(n36099), .A2(n36100), .A3(n36101), .A4(n36102), .ZN(
        n36103) );
  OR4_X1 U731 ( .A1(n36089), .A2(n36094), .A3(n36098), .A4(n36103), .ZN(
        OUTB[7]) );
  AOI22_X1 U732 ( .A1(n36240), .A2(\REGISTERS[30][6] ), .B1(n36237), .B2(
        \REGISTERS[14][6] ), .ZN(n36104) );
  AOI22_X1 U733 ( .A1(n36238), .A2(\REGISTERS[3][6] ), .B1(n36242), .B2(
        \REGISTERS[4][6] ), .ZN(n36105) );
  AOI22_X1 U734 ( .A1(n36250), .A2(\REGISTERS[17][6] ), .B1(n36245), .B2(
        \REGISTERS[22][6] ), .ZN(n36106) );
  AOI22_X1 U735 ( .A1(n36260), .A2(\REGISTERS[15][6] ), .B1(n36258), .B2(
        \REGISTERS[9][6] ), .ZN(n36107) );
  NAND4_X1 U736 ( .A1(n36104), .A2(n36105), .A3(n36106), .A4(n36107), .ZN(
        n36108) );
  AOI22_X1 U737 ( .A1(n36262), .A2(\REGISTERS[16][6] ), .B1(n36263), .B2(
        \REGISTERS[25][6] ), .ZN(n36109) );
  AOI22_X1 U738 ( .A1(n36265), .A2(\REGISTERS[11][6] ), .B1(n36264), .B2(
        \REGISTERS[2][6] ), .ZN(n36110) );
  AOI22_X1 U739 ( .A1(n36267), .A2(\REGISTERS[31][6] ), .B1(n36261), .B2(
        \REGISTERS[13][6] ), .ZN(n36111) );
  AOI22_X1 U740 ( .A1(n36255), .A2(\REGISTERS[29][6] ), .B1(n36259), .B2(
        \REGISTERS[8][6] ), .ZN(n36112) );
  NAND4_X1 U741 ( .A1(n36109), .A2(n36110), .A3(n36111), .A4(n36112), .ZN(
        n36113) );
  AOI22_X1 U742 ( .A1(n36254), .A2(\REGISTERS[26][6] ), .B1(n36256), .B2(
        \REGISTERS[21][6] ), .ZN(n36114) );
  AOI22_X1 U743 ( .A1(n36251), .A2(\REGISTERS[1][6] ), .B1(n36252), .B2(
        \REGISTERS[7][6] ), .ZN(n36115) );
  AOI222_X1 U744 ( .A1(n36248), .A2(\REGISTERS[20][6] ), .B1(n36249), .B2(
        \REGISTERS[5][6] ), .C1(n36247), .C2(\REGISTERS[18][6] ), .ZN(n36116)
         );
  NAND3_X1 U745 ( .A1(n36114), .A2(n36115), .A3(n36116), .ZN(n36117) );
  AOI22_X1 U746 ( .A1(n36244), .A2(\REGISTERS[28][6] ), .B1(n36246), .B2(
        \REGISTERS[19][6] ), .ZN(n36118) );
  AOI22_X1 U747 ( .A1(n36243), .A2(\REGISTERS[6][6] ), .B1(n36257), .B2(
        \REGISTERS[23][6] ), .ZN(n36119) );
  AOI22_X1 U748 ( .A1(n36253), .A2(\REGISTERS[24][6] ), .B1(n36241), .B2(
        \REGISTERS[10][6] ), .ZN(n36120) );
  AOI22_X1 U749 ( .A1(n36239), .A2(\REGISTERS[12][6] ), .B1(n36266), .B2(
        \REGISTERS[27][6] ), .ZN(n36121) );
  NAND4_X1 U750 ( .A1(n36118), .A2(n36119), .A3(n36120), .A4(n36121), .ZN(
        n36122) );
  OR4_X1 U751 ( .A1(n36108), .A2(n36113), .A3(n36117), .A4(n36122), .ZN(
        OUTB[6]) );
  AOI22_X1 U752 ( .A1(n36240), .A2(\REGISTERS[30][5] ), .B1(n36237), .B2(
        \REGISTERS[14][5] ), .ZN(n36123) );
  AOI22_X1 U753 ( .A1(n36238), .A2(\REGISTERS[3][5] ), .B1(n36242), .B2(
        \REGISTERS[4][5] ), .ZN(n36124) );
  AOI22_X1 U754 ( .A1(n36250), .A2(\REGISTERS[17][5] ), .B1(n36245), .B2(
        \REGISTERS[22][5] ), .ZN(n36125) );
  AOI22_X1 U755 ( .A1(n36260), .A2(\REGISTERS[15][5] ), .B1(n36258), .B2(
        \REGISTERS[9][5] ), .ZN(n36126) );
  NAND4_X1 U756 ( .A1(n36123), .A2(n36124), .A3(n36125), .A4(n36126), .ZN(
        n36127) );
  AOI22_X1 U757 ( .A1(n36262), .A2(\REGISTERS[16][5] ), .B1(n36263), .B2(
        \REGISTERS[25][5] ), .ZN(n36128) );
  AOI22_X1 U758 ( .A1(n36265), .A2(\REGISTERS[11][5] ), .B1(n36264), .B2(
        \REGISTERS[2][5] ), .ZN(n36129) );
  AOI22_X1 U759 ( .A1(n36267), .A2(\REGISTERS[31][5] ), .B1(n36261), .B2(
        \REGISTERS[13][5] ), .ZN(n36130) );
  AOI22_X1 U760 ( .A1(n36255), .A2(\REGISTERS[29][5] ), .B1(n36259), .B2(
        \REGISTERS[8][5] ), .ZN(n36131) );
  NAND4_X1 U761 ( .A1(n36128), .A2(n36129), .A3(n36130), .A4(n36131), .ZN(
        n36132) );
  AOI22_X1 U762 ( .A1(n36254), .A2(\REGISTERS[26][5] ), .B1(n36256), .B2(
        \REGISTERS[21][5] ), .ZN(n36133) );
  AOI22_X1 U763 ( .A1(n36251), .A2(\REGISTERS[1][5] ), .B1(n36252), .B2(
        \REGISTERS[7][5] ), .ZN(n36134) );
  AOI222_X1 U764 ( .A1(n36248), .A2(\REGISTERS[20][5] ), .B1(n36249), .B2(
        \REGISTERS[5][5] ), .C1(n36247), .C2(\REGISTERS[18][5] ), .ZN(n36135)
         );
  NAND3_X1 U765 ( .A1(n36133), .A2(n36134), .A3(n36135), .ZN(n36136) );
  AOI22_X1 U766 ( .A1(n36244), .A2(\REGISTERS[28][5] ), .B1(n36246), .B2(
        \REGISTERS[19][5] ), .ZN(n36137) );
  AOI22_X1 U767 ( .A1(n36243), .A2(\REGISTERS[6][5] ), .B1(n36257), .B2(
        \REGISTERS[23][5] ), .ZN(n36138) );
  AOI22_X1 U768 ( .A1(n36253), .A2(\REGISTERS[24][5] ), .B1(n36241), .B2(
        \REGISTERS[10][5] ), .ZN(n36139) );
  AOI22_X1 U769 ( .A1(n36239), .A2(\REGISTERS[12][5] ), .B1(n36266), .B2(
        \REGISTERS[27][5] ), .ZN(n36140) );
  NAND4_X1 U770 ( .A1(n36137), .A2(n36138), .A3(n36139), .A4(n36140), .ZN(
        n36141) );
  OR4_X1 U771 ( .A1(n36127), .A2(n36132), .A3(n36136), .A4(n36141), .ZN(
        OUTB[5]) );
  AOI22_X1 U772 ( .A1(n36240), .A2(\REGISTERS[30][4] ), .B1(n36237), .B2(
        \REGISTERS[14][4] ), .ZN(n36142) );
  AOI22_X1 U773 ( .A1(n36238), .A2(\REGISTERS[3][4] ), .B1(n36242), .B2(
        \REGISTERS[4][4] ), .ZN(n36143) );
  AOI22_X1 U774 ( .A1(n36250), .A2(\REGISTERS[17][4] ), .B1(n36245), .B2(
        \REGISTERS[22][4] ), .ZN(n36144) );
  AOI22_X1 U775 ( .A1(n36260), .A2(\REGISTERS[15][4] ), .B1(n36258), .B2(
        \REGISTERS[9][4] ), .ZN(n36145) );
  NAND4_X1 U776 ( .A1(n36142), .A2(n36143), .A3(n36144), .A4(n36145), .ZN(
        n36146) );
  AOI22_X1 U777 ( .A1(n36262), .A2(\REGISTERS[16][4] ), .B1(n36263), .B2(
        \REGISTERS[25][4] ), .ZN(n36147) );
  AOI22_X1 U778 ( .A1(n36265), .A2(\REGISTERS[11][4] ), .B1(n36264), .B2(
        \REGISTERS[2][4] ), .ZN(n36148) );
  AOI22_X1 U779 ( .A1(n36267), .A2(\REGISTERS[31][4] ), .B1(n36261), .B2(
        \REGISTERS[13][4] ), .ZN(n36149) );
  AOI22_X1 U780 ( .A1(n36255), .A2(\REGISTERS[29][4] ), .B1(n36259), .B2(
        \REGISTERS[8][4] ), .ZN(n36150) );
  NAND4_X1 U781 ( .A1(n36147), .A2(n36148), .A3(n36149), .A4(n36150), .ZN(
        n36151) );
  AOI22_X1 U782 ( .A1(n36254), .A2(\REGISTERS[26][4] ), .B1(n36256), .B2(
        \REGISTERS[21][4] ), .ZN(n36152) );
  AOI22_X1 U783 ( .A1(n36251), .A2(\REGISTERS[1][4] ), .B1(n36252), .B2(
        \REGISTERS[7][4] ), .ZN(n36153) );
  AOI222_X1 U784 ( .A1(n36248), .A2(\REGISTERS[20][4] ), .B1(n36249), .B2(
        \REGISTERS[5][4] ), .C1(n36247), .C2(\REGISTERS[18][4] ), .ZN(n36154)
         );
  NAND3_X1 U785 ( .A1(n36152), .A2(n36153), .A3(n36154), .ZN(n36155) );
  AOI22_X1 U786 ( .A1(n36244), .A2(\REGISTERS[28][4] ), .B1(n36246), .B2(
        \REGISTERS[19][4] ), .ZN(n36156) );
  AOI22_X1 U787 ( .A1(n36243), .A2(\REGISTERS[6][4] ), .B1(n36257), .B2(
        \REGISTERS[23][4] ), .ZN(n36157) );
  AOI22_X1 U788 ( .A1(n36253), .A2(\REGISTERS[24][4] ), .B1(n36241), .B2(
        \REGISTERS[10][4] ), .ZN(n36158) );
  AOI22_X1 U789 ( .A1(n36239), .A2(\REGISTERS[12][4] ), .B1(n36266), .B2(
        \REGISTERS[27][4] ), .ZN(n36159) );
  NAND4_X1 U790 ( .A1(n36156), .A2(n36157), .A3(n36158), .A4(n36159), .ZN(
        n36160) );
  OR4_X1 U791 ( .A1(n36146), .A2(n36151), .A3(n36155), .A4(n36160), .ZN(
        OUTB[4]) );
  AOI22_X1 U792 ( .A1(n36240), .A2(\REGISTERS[30][3] ), .B1(n36237), .B2(
        \REGISTERS[14][3] ), .ZN(n36161) );
  AOI22_X1 U793 ( .A1(n36238), .A2(\REGISTERS[3][3] ), .B1(n36242), .B2(
        \REGISTERS[4][3] ), .ZN(n36162) );
  AOI22_X1 U794 ( .A1(n36250), .A2(\REGISTERS[17][3] ), .B1(n36245), .B2(
        \REGISTERS[22][3] ), .ZN(n36163) );
  AOI22_X1 U795 ( .A1(n36260), .A2(\REGISTERS[15][3] ), .B1(n36258), .B2(
        \REGISTERS[9][3] ), .ZN(n36164) );
  NAND4_X1 U796 ( .A1(n36161), .A2(n36162), .A3(n36163), .A4(n36164), .ZN(
        n36165) );
  AOI22_X1 U797 ( .A1(n36262), .A2(\REGISTERS[16][3] ), .B1(n36263), .B2(
        \REGISTERS[25][3] ), .ZN(n36166) );
  AOI22_X1 U798 ( .A1(n36265), .A2(\REGISTERS[11][3] ), .B1(n36264), .B2(
        \REGISTERS[2][3] ), .ZN(n36167) );
  AOI22_X1 U799 ( .A1(n36855), .A2(\REGISTERS[31][3] ), .B1(n36261), .B2(
        \REGISTERS[13][3] ), .ZN(n36168) );
  AOI22_X1 U800 ( .A1(n36255), .A2(\REGISTERS[29][3] ), .B1(n36259), .B2(
        \REGISTERS[8][3] ), .ZN(n36169) );
  NAND4_X1 U801 ( .A1(n36166), .A2(n36167), .A3(n36168), .A4(n36169), .ZN(
        n36170) );
  AOI22_X1 U802 ( .A1(n36254), .A2(\REGISTERS[26][3] ), .B1(n36256), .B2(
        \REGISTERS[21][3] ), .ZN(n36171) );
  AOI22_X1 U803 ( .A1(n36251), .A2(\REGISTERS[1][3] ), .B1(n36252), .B2(
        \REGISTERS[7][3] ), .ZN(n36172) );
  AOI222_X1 U804 ( .A1(n36248), .A2(\REGISTERS[20][3] ), .B1(n36249), .B2(
        \REGISTERS[5][3] ), .C1(n36247), .C2(\REGISTERS[18][3] ), .ZN(n36173)
         );
  NAND3_X1 U805 ( .A1(n36171), .A2(n36172), .A3(n36173), .ZN(n36174) );
  AOI22_X1 U806 ( .A1(n36244), .A2(\REGISTERS[28][3] ), .B1(n36246), .B2(
        \REGISTERS[19][3] ), .ZN(n36175) );
  AOI22_X1 U807 ( .A1(n36243), .A2(\REGISTERS[6][3] ), .B1(n36257), .B2(
        \REGISTERS[23][3] ), .ZN(n36176) );
  AOI22_X1 U808 ( .A1(n36253), .A2(\REGISTERS[24][3] ), .B1(n36241), .B2(
        \REGISTERS[10][3] ), .ZN(n36177) );
  AOI22_X1 U809 ( .A1(n36239), .A2(\REGISTERS[12][3] ), .B1(n36266), .B2(
        \REGISTERS[27][3] ), .ZN(n36178) );
  NAND4_X1 U810 ( .A1(n36175), .A2(n36176), .A3(n36177), .A4(n36178), .ZN(
        n36179) );
  OR4_X1 U811 ( .A1(n36165), .A2(n36170), .A3(n36174), .A4(n36179), .ZN(
        OUTB[3]) );
  AOI22_X1 U812 ( .A1(n36240), .A2(\REGISTERS[30][2] ), .B1(n36237), .B2(
        \REGISTERS[14][2] ), .ZN(n36180) );
  AOI22_X1 U813 ( .A1(n36238), .A2(\REGISTERS[3][2] ), .B1(n36242), .B2(
        \REGISTERS[4][2] ), .ZN(n36181) );
  AOI22_X1 U814 ( .A1(n36250), .A2(\REGISTERS[17][2] ), .B1(n36245), .B2(
        \REGISTERS[22][2] ), .ZN(n36182) );
  AOI22_X1 U815 ( .A1(n36260), .A2(\REGISTERS[15][2] ), .B1(n36258), .B2(
        \REGISTERS[9][2] ), .ZN(n36183) );
  NAND4_X1 U816 ( .A1(n36180), .A2(n36181), .A3(n36182), .A4(n36183), .ZN(
        n36184) );
  AOI22_X1 U817 ( .A1(n36262), .A2(\REGISTERS[16][2] ), .B1(n36263), .B2(
        \REGISTERS[25][2] ), .ZN(n36185) );
  AOI22_X1 U818 ( .A1(n36265), .A2(\REGISTERS[11][2] ), .B1(n36264), .B2(
        \REGISTERS[2][2] ), .ZN(n36186) );
  AOI22_X1 U819 ( .A1(n36267), .A2(\REGISTERS[31][2] ), .B1(n36261), .B2(
        \REGISTERS[13][2] ), .ZN(n36187) );
  AOI22_X1 U820 ( .A1(n36255), .A2(\REGISTERS[29][2] ), .B1(n36259), .B2(
        \REGISTERS[8][2] ), .ZN(n36188) );
  NAND4_X1 U821 ( .A1(n36185), .A2(n36186), .A3(n36187), .A4(n36188), .ZN(
        n36189) );
  AOI22_X1 U822 ( .A1(n36254), .A2(\REGISTERS[26][2] ), .B1(n36256), .B2(
        \REGISTERS[21][2] ), .ZN(n36190) );
  AOI22_X1 U823 ( .A1(n36251), .A2(\REGISTERS[1][2] ), .B1(n36252), .B2(
        \REGISTERS[7][2] ), .ZN(n36191) );
  AOI222_X1 U824 ( .A1(n36248), .A2(\REGISTERS[20][2] ), .B1(n36249), .B2(
        \REGISTERS[5][2] ), .C1(n36247), .C2(\REGISTERS[18][2] ), .ZN(n36192)
         );
  NAND3_X1 U825 ( .A1(n36190), .A2(n36191), .A3(n36192), .ZN(n36193) );
  AOI22_X1 U826 ( .A1(n36244), .A2(\REGISTERS[28][2] ), .B1(n36246), .B2(
        \REGISTERS[19][2] ), .ZN(n36194) );
  AOI22_X1 U827 ( .A1(n36243), .A2(\REGISTERS[6][2] ), .B1(n36257), .B2(
        \REGISTERS[23][2] ), .ZN(n36195) );
  AOI22_X1 U828 ( .A1(n36253), .A2(\REGISTERS[24][2] ), .B1(n36241), .B2(
        \REGISTERS[10][2] ), .ZN(n36196) );
  AOI22_X1 U829 ( .A1(n36239), .A2(\REGISTERS[12][2] ), .B1(n36266), .B2(
        \REGISTERS[27][2] ), .ZN(n36197) );
  NAND4_X1 U830 ( .A1(n36194), .A2(n36195), .A3(n36196), .A4(n36197), .ZN(
        n36198) );
  OR4_X1 U831 ( .A1(n36184), .A2(n36189), .A3(n36193), .A4(n36198), .ZN(
        OUTB[2]) );
  AOI22_X1 U832 ( .A1(n36240), .A2(\REGISTERS[30][1] ), .B1(n36237), .B2(
        \REGISTERS[14][1] ), .ZN(n36199) );
  AOI22_X1 U833 ( .A1(n36238), .A2(\REGISTERS[3][1] ), .B1(n36242), .B2(
        \REGISTERS[4][1] ), .ZN(n36200) );
  AOI22_X1 U834 ( .A1(n36250), .A2(\REGISTERS[17][1] ), .B1(n36245), .B2(
        \REGISTERS[22][1] ), .ZN(n36201) );
  AOI22_X1 U835 ( .A1(n36260), .A2(\REGISTERS[15][1] ), .B1(n36258), .B2(
        \REGISTERS[9][1] ), .ZN(n36202) );
  NAND4_X1 U836 ( .A1(n36199), .A2(n36200), .A3(n36201), .A4(n36202), .ZN(
        n36203) );
  AOI22_X1 U837 ( .A1(n36262), .A2(\REGISTERS[16][1] ), .B1(n36263), .B2(
        \REGISTERS[25][1] ), .ZN(n36204) );
  AOI22_X1 U838 ( .A1(n36265), .A2(\REGISTERS[11][1] ), .B1(n36264), .B2(
        \REGISTERS[2][1] ), .ZN(n36205) );
  AOI22_X1 U839 ( .A1(n36267), .A2(\REGISTERS[31][1] ), .B1(n36261), .B2(
        \REGISTERS[13][1] ), .ZN(n36206) );
  AOI22_X1 U840 ( .A1(n36255), .A2(\REGISTERS[29][1] ), .B1(n36259), .B2(
        \REGISTERS[8][1] ), .ZN(n36207) );
  NAND4_X1 U841 ( .A1(n36204), .A2(n36205), .A3(n36206), .A4(n36207), .ZN(
        n36208) );
  AOI22_X1 U842 ( .A1(n36254), .A2(\REGISTERS[26][1] ), .B1(n36256), .B2(
        \REGISTERS[21][1] ), .ZN(n36209) );
  AOI22_X1 U843 ( .A1(n36251), .A2(\REGISTERS[1][1] ), .B1(n36252), .B2(
        \REGISTERS[7][1] ), .ZN(n36210) );
  AOI222_X1 U844 ( .A1(n36248), .A2(\REGISTERS[20][1] ), .B1(n36249), .B2(
        \REGISTERS[5][1] ), .C1(n36247), .C2(\REGISTERS[18][1] ), .ZN(n36211)
         );
  NAND3_X1 U845 ( .A1(n36209), .A2(n36210), .A3(n36211), .ZN(n36212) );
  AOI22_X1 U846 ( .A1(n36244), .A2(\REGISTERS[28][1] ), .B1(n36246), .B2(
        \REGISTERS[19][1] ), .ZN(n36213) );
  AOI22_X1 U847 ( .A1(n36243), .A2(\REGISTERS[6][1] ), .B1(n36257), .B2(
        \REGISTERS[23][1] ), .ZN(n36214) );
  AOI22_X1 U848 ( .A1(n36253), .A2(\REGISTERS[24][1] ), .B1(n36241), .B2(
        \REGISTERS[10][1] ), .ZN(n36215) );
  AOI22_X1 U849 ( .A1(n36239), .A2(\REGISTERS[12][1] ), .B1(n36266), .B2(
        \REGISTERS[27][1] ), .ZN(n36216) );
  NAND4_X1 U850 ( .A1(n36213), .A2(n36214), .A3(n36215), .A4(n36216), .ZN(
        n36217) );
  OR4_X1 U851 ( .A1(n36203), .A2(n36208), .A3(n36212), .A4(n36217), .ZN(
        OUTB[1]) );
  AOI22_X1 U852 ( .A1(n36240), .A2(\REGISTERS[30][0] ), .B1(n36237), .B2(
        \REGISTERS[14][0] ), .ZN(n36218) );
  AOI22_X1 U853 ( .A1(n36238), .A2(\REGISTERS[3][0] ), .B1(n36242), .B2(
        \REGISTERS[4][0] ), .ZN(n36219) );
  AOI22_X1 U854 ( .A1(n36250), .A2(\REGISTERS[17][0] ), .B1(n36245), .B2(
        \REGISTERS[22][0] ), .ZN(n36220) );
  AOI22_X1 U855 ( .A1(n36260), .A2(\REGISTERS[15][0] ), .B1(n36258), .B2(
        \REGISTERS[9][0] ), .ZN(n36221) );
  NAND4_X1 U856 ( .A1(n36218), .A2(n36219), .A3(n36220), .A4(n36221), .ZN(
        n36222) );
  AOI22_X1 U857 ( .A1(n36262), .A2(\REGISTERS[16][0] ), .B1(n36263), .B2(
        \REGISTERS[25][0] ), .ZN(n36223) );
  AOI22_X1 U858 ( .A1(n36265), .A2(\REGISTERS[11][0] ), .B1(n36264), .B2(
        \REGISTERS[2][0] ), .ZN(n36224) );
  AOI22_X1 U859 ( .A1(n36267), .A2(\REGISTERS[31][0] ), .B1(n36261), .B2(
        \REGISTERS[13][0] ), .ZN(n36225) );
  AOI22_X1 U860 ( .A1(n36255), .A2(\REGISTERS[29][0] ), .B1(n36259), .B2(
        \REGISTERS[8][0] ), .ZN(n36226) );
  NAND4_X1 U861 ( .A1(n36223), .A2(n36224), .A3(n36225), .A4(n36226), .ZN(
        n36227) );
  AOI22_X1 U862 ( .A1(n36254), .A2(\REGISTERS[26][0] ), .B1(n36256), .B2(
        \REGISTERS[21][0] ), .ZN(n36228) );
  AOI22_X1 U863 ( .A1(n36251), .A2(\REGISTERS[1][0] ), .B1(n36252), .B2(
        \REGISTERS[7][0] ), .ZN(n36229) );
  AOI222_X1 U864 ( .A1(n36248), .A2(\REGISTERS[20][0] ), .B1(n36249), .B2(
        \REGISTERS[5][0] ), .C1(n36247), .C2(\REGISTERS[18][0] ), .ZN(n36230)
         );
  NAND3_X1 U865 ( .A1(n36228), .A2(n36229), .A3(n36230), .ZN(n36231) );
  AOI22_X1 U866 ( .A1(n36244), .A2(\REGISTERS[28][0] ), .B1(n36246), .B2(
        \REGISTERS[19][0] ), .ZN(n36232) );
  AOI22_X1 U867 ( .A1(n36243), .A2(\REGISTERS[6][0] ), .B1(n36257), .B2(
        \REGISTERS[23][0] ), .ZN(n36233) );
  AOI22_X1 U868 ( .A1(n36253), .A2(\REGISTERS[24][0] ), .B1(n36241), .B2(
        \REGISTERS[10][0] ), .ZN(n36234) );
  AOI22_X1 U869 ( .A1(n36239), .A2(\REGISTERS[12][0] ), .B1(n36266), .B2(
        \REGISTERS[27][0] ), .ZN(n36235) );
  NAND4_X1 U870 ( .A1(n36232), .A2(n36233), .A3(n36234), .A4(n36235), .ZN(
        n36236) );
  OR4_X1 U871 ( .A1(n36222), .A2(n36227), .A3(n36231), .A4(n36236), .ZN(
        OUTB[0]) );
  BUF_X2 U872 ( .A(n36844), .Z(n36237) );
  BUF_X2 U873 ( .A(n36845), .Z(n36238) );
  BUF_X2 U874 ( .A(n36841), .Z(n36239) );
  BUF_X2 U875 ( .A(n36843), .Z(n36240) );
  BUF_X2 U876 ( .A(n36840), .Z(n36241) );
  BUF_X2 U877 ( .A(n36846), .Z(n36242) );
  BUF_X2 U878 ( .A(n36837), .Z(n36243) );
  BUF_X2 U879 ( .A(n36835), .Z(n36244) );
  BUF_X2 U880 ( .A(n36848), .Z(n36245) );
  BUF_X2 U881 ( .A(n36836), .Z(n36246) );
  BUF_X2 U882 ( .A(n36834), .Z(n36247) );
  BUF_X2 U883 ( .A(n36832), .Z(n36248) );
  BUF_X2 U884 ( .A(n36833), .Z(n36249) );
  BUF_X2 U885 ( .A(n36847), .Z(n36250) );
  BUF_X2 U886 ( .A(n36830), .Z(n36251) );
  BUF_X2 U887 ( .A(n36831), .Z(n36252) );
  BUF_X2 U888 ( .A(n36839), .Z(n36253) );
  BUF_X2 U889 ( .A(n36828), .Z(n36254) );
  BUF_X2 U890 ( .A(n36857), .Z(n36255) );
  BUF_X2 U891 ( .A(n36829), .Z(n36256) );
  BUF_X2 U892 ( .A(n36838), .Z(n36257) );
  BUF_X2 U893 ( .A(n36850), .Z(n36258) );
  BUF_X2 U894 ( .A(n36858), .Z(n36259) );
  BUF_X2 U895 ( .A(n36849), .Z(n36260) );
  BUF_X2 U896 ( .A(n36856), .Z(n36261) );
  BUF_X2 U897 ( .A(n36851), .Z(n36262) );
  BUF_X2 U898 ( .A(n36852), .Z(n36263) );
  BUF_X2 U899 ( .A(n36854), .Z(n36264) );
  BUF_X2 U900 ( .A(n36853), .Z(n36265) );
  BUF_X2 U901 ( .A(n36842), .Z(n36266) );
  BUF_X2 U902 ( .A(n36855), .Z(n36267) );
  NOR3_X2 U903 ( .A1(ADD_RDA[2]), .A2(n36357), .A3(n36356), .ZN(n36784) );
  BUF_X1 U904 ( .A(n36784), .Z(n36286) );
  BUF_X1 U905 ( .A(n36771), .Z(n36277) );
  BUF_X1 U906 ( .A(n36760), .Z(n36270) );
  BUF_X1 U907 ( .A(n36800), .Z(n36298) );
  BUF_X1 U908 ( .A(n36787), .Z(n36289) );
  BUF_X1 U909 ( .A(n36788), .Z(n36290) );
  BUF_X1 U910 ( .A(n36786), .Z(n36288) );
  BUF_X1 U911 ( .A(n36782), .Z(n36284) );
  BUF_X1 U912 ( .A(n36776), .Z(n36282) );
  BUF_X1 U913 ( .A(n36763), .Z(n36273) );
  BUF_X1 U914 ( .A(n36761), .Z(n36271) );
  BUF_X1 U915 ( .A(n36759), .Z(n36269) );
  BUF_X1 U916 ( .A(n36798), .Z(n36296) );
  BUF_X1 U917 ( .A(n36796), .Z(n36294) );
  BUF_X1 U918 ( .A(n36794), .Z(n36292) );
  BUF_X1 U919 ( .A(n36772), .Z(n36278) );
  BUF_X1 U920 ( .A(n36783), .Z(n36285) );
  BUF_X1 U921 ( .A(n36764), .Z(n36274) );
  BUF_X1 U922 ( .A(n36762), .Z(n36272) );
  BUF_X1 U923 ( .A(n36775), .Z(n36281) );
  BUF_X1 U924 ( .A(n36799), .Z(n36297) );
  BUF_X1 U925 ( .A(n36797), .Z(n36295) );
  BUF_X1 U926 ( .A(n36795), .Z(n36293) );
  BUF_X1 U927 ( .A(n36793), .Z(n36291) );
  BUF_X1 U928 ( .A(n36781), .Z(n36283) );
  BUF_X1 U929 ( .A(n36773), .Z(n36279) );
  BUF_X1 U930 ( .A(n36774), .Z(n36280) );
  BUF_X1 U931 ( .A(n36769), .Z(n36275) );
  BUF_X1 U932 ( .A(n36770), .Z(n36276) );
  BUF_X1 U933 ( .A(n36758), .Z(n36268) );
  BUF_X1 U934 ( .A(n36785), .Z(n36287) );
  INV_X1 U935 ( .A(ADD_RDA[2]), .ZN(n36352) );
  INV_X1 U936 ( .A(ADD_RDA[4]), .ZN(n36350) );
  INV_X1 U937 ( .A(ADD_RDA[1]), .ZN(n36357) );
  INV_X1 U938 ( .A(ADD_RDB[3]), .ZN(n36810) );
  OR4_X1 U939 ( .A1(n36717), .A2(n36716), .A3(n36715), .A4(n36714), .ZN(
        OUTA[6]) );
  OR4_X1 U940 ( .A1(n36697), .A2(n36696), .A3(n36695), .A4(n36694), .ZN(
        OUTA[5]) );
  OR4_X1 U941 ( .A1(n36657), .A2(n36656), .A3(n36655), .A4(n36654), .ZN(
        OUTA[3]) );
  OR4_X1 U942 ( .A1(n36677), .A2(n36676), .A3(n36675), .A4(n36674), .ZN(
        OUTA[4]) );
  OR4_X1 U943 ( .A1(n36637), .A2(n36636), .A3(n36635), .A4(n36634), .ZN(
        OUTA[30]) );
  OR4_X1 U944 ( .A1(n36511), .A2(n36510), .A3(n36509), .A4(n36508), .ZN(
        OUTA[1]) );
  OR4_X1 U945 ( .A1(n36427), .A2(n36426), .A3(n36425), .A4(n36424), .ZN(
        OUTA[12]) );
  OR4_X1 U946 ( .A1(n36447), .A2(n36446), .A3(n36445), .A4(n36444), .ZN(
        OUTA[13]) );
  OR4_X1 U947 ( .A1(n36387), .A2(n36386), .A3(n36385), .A4(n36384), .ZN(
        OUTA[10]) );
  OR4_X1 U948 ( .A1(n36407), .A2(n36406), .A3(n36405), .A4(n36404), .ZN(
        OUTA[11]) );
  OR4_X1 U949 ( .A1(n36467), .A2(n36466), .A3(n36465), .A4(n36464), .ZN(
        OUTA[14]) );
  OR4_X1 U950 ( .A1(n36487), .A2(n36486), .A3(n36485), .A4(n36484), .ZN(
        OUTA[15]) );
  OR4_X1 U951 ( .A1(n36737), .A2(n36736), .A3(n36735), .A4(n36734), .ZN(
        OUTA[7]) );
  OR4_X1 U952 ( .A1(n36577), .A2(n36576), .A3(n36575), .A4(n36574), .ZN(
        OUTA[28]) );
  OR4_X1 U953 ( .A1(n36537), .A2(n36536), .A3(n36535), .A4(n36534), .ZN(
        OUTA[26]) );
  OR4_X1 U954 ( .A1(n36557), .A2(n36556), .A3(n36555), .A4(n36554), .ZN(
        OUTA[27]) );
  OR4_X1 U955 ( .A1(n36617), .A2(n36616), .A3(n36615), .A4(n36614), .ZN(
        OUTA[2]) );
  OR4_X1 U956 ( .A1(n36597), .A2(n36596), .A3(n36595), .A4(n36594), .ZN(
        OUTA[29]) );
  OR4_X1 U957 ( .A1(n36757), .A2(n36756), .A3(n36755), .A4(n36754), .ZN(
        OUTA[8]) );
  OR4_X1 U958 ( .A1(n36808), .A2(n36807), .A3(n36806), .A4(n36805), .ZN(
        OUTA[9]) );
  NOR2_X1 U959 ( .A1(n36349), .A2(n36358), .ZN(n36764) );
  BUF_X1 U960 ( .A(N288), .Z(n36316) );
  BUF_X1 U961 ( .A(N300), .Z(n36304) );
  BUF_X1 U962 ( .A(N287), .Z(n36317) );
  BUF_X1 U963 ( .A(N283), .Z(n36321) );
  BUF_X1 U964 ( .A(N284), .Z(n36320) );
  BUF_X1 U965 ( .A(N285), .Z(n36319) );
  BUF_X1 U966 ( .A(N301), .Z(n36303) );
  BUF_X1 U967 ( .A(N286), .Z(n36318) );
  BUF_X1 U968 ( .A(N293), .Z(n36311) );
  BUF_X1 U969 ( .A(N294), .Z(n36310) );
  BUF_X1 U970 ( .A(N295), .Z(n36309) );
  BUF_X1 U971 ( .A(N296), .Z(n36308) );
  BUF_X1 U972 ( .A(N289), .Z(n36315) );
  BUF_X1 U973 ( .A(N299), .Z(n36305) );
  BUF_X1 U974 ( .A(N290), .Z(n36314) );
  BUF_X1 U975 ( .A(N291), .Z(n36313) );
  BUF_X1 U976 ( .A(N298), .Z(n36306) );
  BUF_X1 U977 ( .A(N297), .Z(n36307) );
  BUF_X1 U978 ( .A(N292), .Z(n36312) );
  BUF_X1 U979 ( .A(N276), .Z(n36328) );
  BUF_X1 U980 ( .A(N277), .Z(n36327) );
  BUF_X1 U981 ( .A(N305), .Z(n36299) );
  BUF_X1 U982 ( .A(N243), .Z(n36329) );
  BUF_X1 U983 ( .A(N278), .Z(n36326) );
  BUF_X1 U984 ( .A(N302), .Z(n36302) );
  BUF_X1 U985 ( .A(N303), .Z(n36301) );
  BUF_X1 U986 ( .A(N304), .Z(n36300) );
  BUF_X1 U987 ( .A(N282), .Z(n36322) );
  BUF_X1 U988 ( .A(N281), .Z(n36323) );
  BUF_X1 U989 ( .A(N280), .Z(n36324) );
  INV_X1 U990 ( .A(ADD_WR[0]), .ZN(n36332) );
  BUF_X1 U991 ( .A(N279), .Z(n36325) );
  AND2_X1 U992 ( .A1(RESET), .A2(DATAIN[6]), .ZN(N250) );
  AND2_X1 U993 ( .A1(RESET), .A2(DATAIN[5]), .ZN(N249) );
  AND2_X1 U994 ( .A1(RESET), .A2(DATAIN[3]), .ZN(N247) );
  AND2_X1 U995 ( .A1(RESET), .A2(DATAIN[17]), .ZN(N261) );
  AND2_X1 U996 ( .A1(RESET), .A2(DATAIN[18]), .ZN(N262) );
  AND2_X1 U997 ( .A1(RESET), .A2(DATAIN[19]), .ZN(N263) );
  AND2_X1 U998 ( .A1(RESET), .A2(DATAIN[16]), .ZN(N260) );
  AND2_X1 U999 ( .A1(RESET), .A2(DATAIN[15]), .ZN(N259) );
  AND2_X1 U1000 ( .A1(RESET), .A2(DATAIN[14]), .ZN(N258) );
  AND2_X1 U1001 ( .A1(RESET), .A2(DATAIN[13]), .ZN(N257) );
  AND2_X1 U1002 ( .A1(RESET), .A2(DATAIN[24]), .ZN(N268) );
  AND2_X1 U1003 ( .A1(RESET), .A2(DATAIN[20]), .ZN(N264) );
  AND2_X1 U1004 ( .A1(RESET), .A2(DATAIN[12]), .ZN(N256) );
  AND2_X1 U1005 ( .A1(RESET), .A2(DATAIN[11]), .ZN(N255) );
  AND2_X1 U1006 ( .A1(RESET), .A2(DATAIN[10]), .ZN(N254) );
  AND2_X1 U1007 ( .A1(RESET), .A2(DATAIN[9]), .ZN(N253) );
  AND2_X1 U1008 ( .A1(RESET), .A2(DATAIN[8]), .ZN(N252) );
  AND2_X1 U1009 ( .A1(RESET), .A2(DATAIN[7]), .ZN(N251) );
  AND2_X1 U1010 ( .A1(RESET), .A2(DATAIN[27]), .ZN(N271) );
  AND2_X1 U1011 ( .A1(RESET), .A2(DATAIN[26]), .ZN(N270) );
  AND2_X1 U1012 ( .A1(RESET), .A2(DATAIN[4]), .ZN(N248) );
  AND2_X1 U1013 ( .A1(RESET), .A2(DATAIN[30]), .ZN(N274) );
  AND2_X1 U1014 ( .A1(RESET), .A2(DATAIN[2]), .ZN(N246) );
  AND2_X1 U1015 ( .A1(RESET), .A2(DATAIN[1]), .ZN(N245) );
  AND2_X1 U1016 ( .A1(RESET), .A2(DATAIN[0]), .ZN(N244) );
  AND2_X1 U1017 ( .A1(RESET), .A2(DATAIN[31]), .ZN(N275) );
  AND2_X1 U1018 ( .A1(RESET), .A2(DATAIN[25]), .ZN(N269) );
  AND2_X1 U1019 ( .A1(RESET), .A2(DATAIN[29]), .ZN(N273) );
  AND2_X1 U1020 ( .A1(RESET), .A2(DATAIN[28]), .ZN(N272) );
  AND2_X1 U1021 ( .A1(RESET), .A2(DATAIN[22]), .ZN(N266) );
  AND2_X1 U1022 ( .A1(RESET), .A2(DATAIN[21]), .ZN(N265) );
  AND2_X1 U1023 ( .A1(RESET), .A2(DATAIN[23]), .ZN(N267) );
  NOR2_X1 U1024 ( .A1(n36823), .A2(n36826), .ZN(n36855) );
  NAND3_X1 U1025 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(ADD_WR[2]), .ZN(n36340)
         );
  NAND3_X1 U1026 ( .A1(WE), .A2(ADD_WR[3]), .A3(ADD_WR[4]), .ZN(n36334) );
  OAI21_X1 U1027 ( .B1(n36340), .B2(n36334), .A(RESET), .ZN(N243) );
  NAND3_X1 U1028 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n36332), .ZN(n36341) );
  OAI21_X1 U1029 ( .B1(n36334), .B2(n36341), .A(RESET), .ZN(N276) );
  INV_X1 U1030 ( .A(ADD_WR[1]), .ZN(n36330) );
  NAND3_X1 U1031 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n36330), .ZN(n36342) );
  OAI21_X1 U1032 ( .B1(n36334), .B2(n36342), .A(RESET), .ZN(N277) );
  NAND3_X1 U1033 ( .A1(ADD_WR[2]), .A2(n36332), .A3(n36330), .ZN(n36343) );
  OAI21_X1 U1034 ( .B1(n36334), .B2(n36343), .A(RESET), .ZN(N278) );
  NOR2_X1 U1035 ( .A1(ADD_WR[2]), .A2(n36330), .ZN(n36331) );
  NAND2_X1 U1036 ( .A1(ADD_WR[0]), .A2(n36331), .ZN(n36344) );
  OAI21_X1 U1037 ( .B1(n36334), .B2(n36344), .A(RESET), .ZN(N279) );
  NAND2_X1 U1038 ( .A1(n36331), .A2(n36332), .ZN(n36345) );
  OAI21_X1 U1039 ( .B1(n36334), .B2(n36345), .A(RESET), .ZN(N280) );
  NOR2_X1 U1040 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .ZN(n36333) );
  NAND2_X1 U1041 ( .A1(ADD_WR[0]), .A2(n36333), .ZN(n36347) );
  OAI21_X1 U1042 ( .B1(n36334), .B2(n36347), .A(RESET), .ZN(N281) );
  NAND2_X1 U1043 ( .A1(n36333), .A2(n36332), .ZN(n36337) );
  OAI21_X1 U1044 ( .B1(n36334), .B2(n36337), .A(RESET), .ZN(N282) );
  INV_X1 U1045 ( .A(ADD_WR[3]), .ZN(n36339) );
  NAND3_X1 U1046 ( .A1(WE), .A2(ADD_WR[4]), .A3(n36339), .ZN(n36335) );
  OAI21_X1 U1047 ( .B1(n36340), .B2(n36335), .A(RESET), .ZN(N283) );
  OAI21_X1 U1048 ( .B1(n36341), .B2(n36335), .A(RESET), .ZN(N284) );
  OAI21_X1 U1049 ( .B1(n36342), .B2(n36335), .A(RESET), .ZN(N285) );
  OAI21_X1 U1050 ( .B1(n36343), .B2(n36335), .A(RESET), .ZN(N286) );
  OAI21_X1 U1051 ( .B1(n36344), .B2(n36335), .A(RESET), .ZN(N287) );
  OAI21_X1 U1052 ( .B1(n36345), .B2(n36335), .A(RESET), .ZN(N288) );
  OAI21_X1 U1053 ( .B1(n36347), .B2(n36335), .A(RESET), .ZN(N289) );
  OAI21_X1 U1054 ( .B1(n36337), .B2(n36335), .A(RESET), .ZN(N290) );
  INV_X1 U1055 ( .A(ADD_WR[4]), .ZN(n36338) );
  NAND3_X1 U1056 ( .A1(ADD_WR[3]), .A2(WE), .A3(n36338), .ZN(n36336) );
  OAI21_X1 U1057 ( .B1(n36340), .B2(n36336), .A(RESET), .ZN(N291) );
  OAI21_X1 U1058 ( .B1(n36341), .B2(n36336), .A(RESET), .ZN(N292) );
  OAI21_X1 U1059 ( .B1(n36342), .B2(n36336), .A(RESET), .ZN(N293) );
  OAI21_X1 U1060 ( .B1(n36343), .B2(n36336), .A(RESET), .ZN(N294) );
  OAI21_X1 U1061 ( .B1(n36344), .B2(n36336), .A(RESET), .ZN(N295) );
  OAI21_X1 U1062 ( .B1(n36345), .B2(n36336), .A(RESET), .ZN(N296) );
  OAI21_X1 U1063 ( .B1(n36347), .B2(n36336), .A(RESET), .ZN(N297) );
  OAI21_X1 U1064 ( .B1(n36337), .B2(n36336), .A(RESET), .ZN(N298) );
  NAND3_X1 U1065 ( .A1(WE), .A2(n36339), .A3(n36338), .ZN(n36346) );
  OAI21_X1 U1066 ( .B1(n36340), .B2(n36346), .A(RESET), .ZN(N299) );
  OAI21_X1 U1067 ( .B1(n36341), .B2(n36346), .A(RESET), .ZN(N300) );
  OAI21_X1 U1068 ( .B1(n36342), .B2(n36346), .A(RESET), .ZN(N301) );
  OAI21_X1 U1069 ( .B1(n36343), .B2(n36346), .A(RESET), .ZN(N302) );
  OAI21_X1 U1070 ( .B1(n36344), .B2(n36346), .A(RESET), .ZN(N303) );
  OAI21_X1 U1071 ( .B1(n36345), .B2(n36346), .A(RESET), .ZN(N304) );
  OAI21_X1 U1072 ( .B1(n36347), .B2(n36346), .A(RESET), .ZN(N305) );
  NAND3_X1 U1073 ( .A1(RESET), .A2(ADD_RDA[2]), .A3(n36357), .ZN(n36365) );
  INV_X1 U1074 ( .A(ADD_RDA[3]), .ZN(n36348) );
  NAND3_X1 U1075 ( .A1(ADD_RDA[0]), .A2(n36350), .A3(n36348), .ZN(n36360) );
  NOR2_X1 U1076 ( .A1(n36365), .A2(n36360), .ZN(n36759) );
  NOR2_X1 U1077 ( .A1(ADD_RDA[3]), .A2(ADD_RDA[0]), .ZN(n36351) );
  NAND2_X1 U1078 ( .A1(ADD_RDA[4]), .A2(n36351), .ZN(n36364) );
  NAND3_X1 U1079 ( .A1(RESET), .A2(ADD_RDA[1]), .A3(ADD_RDA[2]), .ZN(n36367)
         );
  NOR2_X1 U1080 ( .A1(n36364), .A2(n36367), .ZN(n36758) );
  NAND3_X1 U1081 ( .A1(ADD_RDA[4]), .A2(ADD_RDA[3]), .A3(ADD_RDA[0]), .ZN(
        n36359) );
  NAND3_X1 U1082 ( .A1(RESET), .A2(n36357), .A3(n36352), .ZN(n36363) );
  NOR2_X1 U1083 ( .A1(n36359), .A2(n36363), .ZN(n36761) );
  NAND3_X1 U1084 ( .A1(ADD_RDA[4]), .A2(ADD_RDA[0]), .A3(n36348), .ZN(n36349)
         );
  NOR2_X1 U1085 ( .A1(n36349), .A2(n36365), .ZN(n36760) );
  NOR2_X1 U1086 ( .A1(n36349), .A2(n36363), .ZN(n36763) );
  NOR2_X1 U1087 ( .A1(n36349), .A2(n36367), .ZN(n36762) );
  NAND3_X1 U1088 ( .A1(ADD_RDA[1]), .A2(RESET), .A3(n36352), .ZN(n36358) );
  INV_X1 U1089 ( .A(ADD_RDA[0]), .ZN(n36354) );
  NAND3_X1 U1090 ( .A1(ADD_RDA[3]), .A2(n36350), .A3(n36354), .ZN(n36361) );
  NOR2_X1 U1091 ( .A1(n36367), .A2(n36361), .ZN(n36770) );
  NAND3_X1 U1092 ( .A1(ADD_RDA[3]), .A2(ADD_RDA[0]), .A3(n36350), .ZN(n36366)
         );
  NOR2_X1 U1093 ( .A1(n36365), .A2(n36366), .ZN(n36769) );
  NOR2_X1 U1094 ( .A1(n36358), .A2(n36359), .ZN(n36772) );
  NAND3_X1 U1095 ( .A1(RESET), .A2(n36351), .A3(n36350), .ZN(n36356) );
  NOR3_X1 U1096 ( .A1(ADD_RDA[1]), .A2(n36352), .A3(n36356), .ZN(n36771) );
  AOI22_X1 U1097 ( .A1(\REGISTERS[27][0] ), .A2(n36278), .B1(\REGISTERS[4][0] ), .B2(n36277), .ZN(n36355) );
  NAND2_X1 U1098 ( .A1(ADD_RDA[1]), .A2(ADD_RDA[2]), .ZN(n36353) );
  NOR2_X1 U1099 ( .A1(n36353), .A2(n36356), .ZN(n36774) );
  NAND3_X1 U1100 ( .A1(ADD_RDA[3]), .A2(ADD_RDA[4]), .A3(n36354), .ZN(n36362)
         );
  NOR2_X1 U1101 ( .A1(n36365), .A2(n36362), .ZN(n36773) );
  NOR2_X1 U1102 ( .A1(n36358), .A2(n36362), .ZN(n36776) );
  NOR2_X1 U1103 ( .A1(n36360), .A2(n36367), .ZN(n36775) );
  NOR2_X1 U1104 ( .A1(n36358), .A2(n36361), .ZN(n36782) );
  NOR2_X1 U1105 ( .A1(n36363), .A2(n36366), .ZN(n36781) );
  NOR2_X1 U1106 ( .A1(n36358), .A2(n36364), .ZN(n36783) );
  NOR2_X1 U1107 ( .A1(n36358), .A2(n36360), .ZN(n36786) );
  NOR2_X1 U1108 ( .A1(n36367), .A2(n36359), .ZN(n36785) );
  NOR2_X1 U1109 ( .A1(n36367), .A2(n36362), .ZN(n36788) );
  NOR2_X1 U1110 ( .A1(n36363), .A2(n36361), .ZN(n36787) );
  NOR2_X1 U1111 ( .A1(n36358), .A2(n36366), .ZN(n36794) );
  NOR2_X1 U1112 ( .A1(n36365), .A2(n36359), .ZN(n36793) );
  NOR2_X1 U1113 ( .A1(n36360), .A2(n36363), .ZN(n36796) );
  NOR2_X1 U1114 ( .A1(n36364), .A2(n36363), .ZN(n36795) );
  NOR2_X1 U1115 ( .A1(n36365), .A2(n36361), .ZN(n36798) );
  NOR2_X1 U1116 ( .A1(n36363), .A2(n36362), .ZN(n36797) );
  NOR2_X1 U1117 ( .A1(n36365), .A2(n36364), .ZN(n36800) );
  NOR2_X1 U1118 ( .A1(n36367), .A2(n36366), .ZN(n36799) );
  AOI22_X1 U1119 ( .A1(n36269), .A2(\REGISTERS[5][10] ), .B1(n36268), .B2(
        \REGISTERS[22][10] ), .ZN(n36371) );
  AOI22_X1 U1120 ( .A1(n36271), .A2(\REGISTERS[25][10] ), .B1(n36270), .B2(
        \REGISTERS[21][10] ), .ZN(n36370) );
  AOI22_X1 U1121 ( .A1(n36273), .A2(\REGISTERS[17][10] ), .B1(n36272), .B2(
        \REGISTERS[23][10] ), .ZN(n36369) );
  NAND2_X1 U1122 ( .A1(n36274), .A2(\REGISTERS[19][10] ), .ZN(n36368) );
  NAND4_X1 U1123 ( .A1(n36371), .A2(n36370), .A3(n36369), .A4(n36368), .ZN(
        n36387) );
  AOI22_X1 U1124 ( .A1(n36276), .A2(\REGISTERS[14][10] ), .B1(n36275), .B2(
        \REGISTERS[13][10] ), .ZN(n36375) );
  AOI22_X1 U1125 ( .A1(n36278), .A2(\REGISTERS[27][10] ), .B1(n36277), .B2(
        \REGISTERS[4][10] ), .ZN(n36374) );
  AOI22_X1 U1126 ( .A1(n36280), .A2(\REGISTERS[6][10] ), .B1(n36279), .B2(
        \REGISTERS[28][10] ), .ZN(n36373) );
  AOI22_X1 U1127 ( .A1(n36282), .A2(\REGISTERS[26][10] ), .B1(n36281), .B2(
        \REGISTERS[7][10] ), .ZN(n36372) );
  NAND4_X1 U1128 ( .A1(n36375), .A2(n36374), .A3(n36373), .A4(n36372), .ZN(
        n36386) );
  AOI22_X1 U1129 ( .A1(n36284), .A2(\REGISTERS[10][10] ), .B1(n36283), .B2(
        \REGISTERS[9][10] ), .ZN(n36379) );
  AOI22_X1 U1130 ( .A1(n36286), .A2(\REGISTERS[2][10] ), .B1(n36285), .B2(
        \REGISTERS[18][10] ), .ZN(n36378) );
  AOI22_X1 U1131 ( .A1(n36288), .A2(\REGISTERS[3][10] ), .B1(n36287), .B2(
        \REGISTERS[31][10] ), .ZN(n36377) );
  AOI22_X1 U1132 ( .A1(n36290), .A2(\REGISTERS[30][10] ), .B1(n36289), .B2(
        \REGISTERS[8][10] ), .ZN(n36376) );
  NAND4_X1 U1133 ( .A1(n36379), .A2(n36378), .A3(n36377), .A4(n36376), .ZN(
        n36385) );
  AOI22_X1 U1134 ( .A1(n36292), .A2(\REGISTERS[11][10] ), .B1(n36291), .B2(
        \REGISTERS[29][10] ), .ZN(n36383) );
  AOI22_X1 U1135 ( .A1(n36294), .A2(\REGISTERS[1][10] ), .B1(n36293), .B2(
        \REGISTERS[16][10] ), .ZN(n36382) );
  AOI22_X1 U1136 ( .A1(n36296), .A2(\REGISTERS[12][10] ), .B1(n36295), .B2(
        \REGISTERS[24][10] ), .ZN(n36381) );
  AOI22_X1 U1137 ( .A1(n36298), .A2(\REGISTERS[20][10] ), .B1(n36297), .B2(
        \REGISTERS[15][10] ), .ZN(n36380) );
  NAND4_X1 U1138 ( .A1(n36383), .A2(n36382), .A3(n36381), .A4(n36380), .ZN(
        n36384) );
  AOI22_X1 U1139 ( .A1(n36269), .A2(\REGISTERS[5][11] ), .B1(n36268), .B2(
        \REGISTERS[22][11] ), .ZN(n36391) );
  AOI22_X1 U1140 ( .A1(n36271), .A2(\REGISTERS[25][11] ), .B1(n36270), .B2(
        \REGISTERS[21][11] ), .ZN(n36390) );
  AOI22_X1 U1141 ( .A1(n36273), .A2(\REGISTERS[17][11] ), .B1(n36272), .B2(
        \REGISTERS[23][11] ), .ZN(n36389) );
  NAND2_X1 U1142 ( .A1(n36274), .A2(\REGISTERS[19][11] ), .ZN(n36388) );
  NAND4_X1 U1143 ( .A1(n36391), .A2(n36390), .A3(n36389), .A4(n36388), .ZN(
        n36407) );
  AOI22_X1 U1144 ( .A1(n36276), .A2(\REGISTERS[14][11] ), .B1(n36275), .B2(
        \REGISTERS[13][11] ), .ZN(n36395) );
  AOI22_X1 U1145 ( .A1(n36278), .A2(\REGISTERS[27][11] ), .B1(n36277), .B2(
        \REGISTERS[4][11] ), .ZN(n36394) );
  AOI22_X1 U1146 ( .A1(n36280), .A2(\REGISTERS[6][11] ), .B1(n36279), .B2(
        \REGISTERS[28][11] ), .ZN(n36393) );
  AOI22_X1 U1147 ( .A1(n36282), .A2(\REGISTERS[26][11] ), .B1(n36281), .B2(
        \REGISTERS[7][11] ), .ZN(n36392) );
  NAND4_X1 U1148 ( .A1(n36395), .A2(n36394), .A3(n36393), .A4(n36392), .ZN(
        n36406) );
  AOI22_X1 U1149 ( .A1(n36284), .A2(\REGISTERS[10][11] ), .B1(n36283), .B2(
        \REGISTERS[9][11] ), .ZN(n36399) );
  AOI22_X1 U1150 ( .A1(n36286), .A2(\REGISTERS[2][11] ), .B1(n36285), .B2(
        \REGISTERS[18][11] ), .ZN(n36398) );
  AOI22_X1 U1151 ( .A1(n36288), .A2(\REGISTERS[3][11] ), .B1(n36287), .B2(
        \REGISTERS[31][11] ), .ZN(n36397) );
  AOI22_X1 U1152 ( .A1(n36290), .A2(\REGISTERS[30][11] ), .B1(n36289), .B2(
        \REGISTERS[8][11] ), .ZN(n36396) );
  NAND4_X1 U1153 ( .A1(n36399), .A2(n36398), .A3(n36397), .A4(n36396), .ZN(
        n36405) );
  AOI22_X1 U1154 ( .A1(n36292), .A2(\REGISTERS[11][11] ), .B1(n36291), .B2(
        \REGISTERS[29][11] ), .ZN(n36403) );
  AOI22_X1 U1155 ( .A1(n36294), .A2(\REGISTERS[1][11] ), .B1(n36293), .B2(
        \REGISTERS[16][11] ), .ZN(n36402) );
  AOI22_X1 U1156 ( .A1(n36296), .A2(\REGISTERS[12][11] ), .B1(n36295), .B2(
        \REGISTERS[24][11] ), .ZN(n36401) );
  AOI22_X1 U1157 ( .A1(n36298), .A2(\REGISTERS[20][11] ), .B1(n36297), .B2(
        \REGISTERS[15][11] ), .ZN(n36400) );
  NAND4_X1 U1158 ( .A1(n36403), .A2(n36402), .A3(n36401), .A4(n36400), .ZN(
        n36404) );
  AOI22_X1 U1159 ( .A1(n36269), .A2(\REGISTERS[5][12] ), .B1(n36268), .B2(
        \REGISTERS[22][12] ), .ZN(n36411) );
  AOI22_X1 U1160 ( .A1(n36271), .A2(\REGISTERS[25][12] ), .B1(n36270), .B2(
        \REGISTERS[21][12] ), .ZN(n36410) );
  AOI22_X1 U1161 ( .A1(n36273), .A2(\REGISTERS[17][12] ), .B1(n36272), .B2(
        \REGISTERS[23][12] ), .ZN(n36409) );
  NAND2_X1 U1162 ( .A1(n36274), .A2(\REGISTERS[19][12] ), .ZN(n36408) );
  NAND4_X1 U1163 ( .A1(n36411), .A2(n36410), .A3(n36409), .A4(n36408), .ZN(
        n36427) );
  AOI22_X1 U1164 ( .A1(n36276), .A2(\REGISTERS[14][12] ), .B1(n36275), .B2(
        \REGISTERS[13][12] ), .ZN(n36415) );
  AOI22_X1 U1165 ( .A1(n36278), .A2(\REGISTERS[27][12] ), .B1(n36277), .B2(
        \REGISTERS[4][12] ), .ZN(n36414) );
  AOI22_X1 U1166 ( .A1(n36280), .A2(\REGISTERS[6][12] ), .B1(n36279), .B2(
        \REGISTERS[28][12] ), .ZN(n36413) );
  AOI22_X1 U1167 ( .A1(n36282), .A2(\REGISTERS[26][12] ), .B1(n36281), .B2(
        \REGISTERS[7][12] ), .ZN(n36412) );
  NAND4_X1 U1168 ( .A1(n36415), .A2(n36414), .A3(n36413), .A4(n36412), .ZN(
        n36426) );
  AOI22_X1 U1169 ( .A1(n36284), .A2(\REGISTERS[10][12] ), .B1(n36283), .B2(
        \REGISTERS[9][12] ), .ZN(n36419) );
  AOI22_X1 U1170 ( .A1(n36286), .A2(\REGISTERS[2][12] ), .B1(n36285), .B2(
        \REGISTERS[18][12] ), .ZN(n36418) );
  AOI22_X1 U1171 ( .A1(n36288), .A2(\REGISTERS[3][12] ), .B1(n36287), .B2(
        \REGISTERS[31][12] ), .ZN(n36417) );
  AOI22_X1 U1172 ( .A1(n36290), .A2(\REGISTERS[30][12] ), .B1(n36289), .B2(
        \REGISTERS[8][12] ), .ZN(n36416) );
  NAND4_X1 U1173 ( .A1(n36419), .A2(n36418), .A3(n36417), .A4(n36416), .ZN(
        n36425) );
  AOI22_X1 U1174 ( .A1(n36292), .A2(\REGISTERS[11][12] ), .B1(n36291), .B2(
        \REGISTERS[29][12] ), .ZN(n36423) );
  AOI22_X1 U1175 ( .A1(n36294), .A2(\REGISTERS[1][12] ), .B1(n36293), .B2(
        \REGISTERS[16][12] ), .ZN(n36422) );
  AOI22_X1 U1176 ( .A1(n36296), .A2(\REGISTERS[12][12] ), .B1(n36295), .B2(
        \REGISTERS[24][12] ), .ZN(n36421) );
  AOI22_X1 U1177 ( .A1(n36298), .A2(\REGISTERS[20][12] ), .B1(n36297), .B2(
        \REGISTERS[15][12] ), .ZN(n36420) );
  NAND4_X1 U1178 ( .A1(n36423), .A2(n36422), .A3(n36421), .A4(n36420), .ZN(
        n36424) );
  AOI22_X1 U1179 ( .A1(n36269), .A2(\REGISTERS[5][13] ), .B1(n36268), .B2(
        \REGISTERS[22][13] ), .ZN(n36431) );
  AOI22_X1 U1180 ( .A1(n36271), .A2(\REGISTERS[25][13] ), .B1(n36270), .B2(
        \REGISTERS[21][13] ), .ZN(n36430) );
  AOI22_X1 U1181 ( .A1(n36273), .A2(\REGISTERS[17][13] ), .B1(n36272), .B2(
        \REGISTERS[23][13] ), .ZN(n36429) );
  NAND2_X1 U1182 ( .A1(n36274), .A2(\REGISTERS[19][13] ), .ZN(n36428) );
  NAND4_X1 U1183 ( .A1(n36431), .A2(n36430), .A3(n36429), .A4(n36428), .ZN(
        n36447) );
  AOI22_X1 U1184 ( .A1(n36276), .A2(\REGISTERS[14][13] ), .B1(n36275), .B2(
        \REGISTERS[13][13] ), .ZN(n36435) );
  AOI22_X1 U1185 ( .A1(n36278), .A2(\REGISTERS[27][13] ), .B1(n36277), .B2(
        \REGISTERS[4][13] ), .ZN(n36434) );
  AOI22_X1 U1186 ( .A1(n36280), .A2(\REGISTERS[6][13] ), .B1(n36279), .B2(
        \REGISTERS[28][13] ), .ZN(n36433) );
  AOI22_X1 U1187 ( .A1(n36282), .A2(\REGISTERS[26][13] ), .B1(n36281), .B2(
        \REGISTERS[7][13] ), .ZN(n36432) );
  NAND4_X1 U1188 ( .A1(n36435), .A2(n36434), .A3(n36433), .A4(n36432), .ZN(
        n36446) );
  AOI22_X1 U1189 ( .A1(n36284), .A2(\REGISTERS[10][13] ), .B1(n36283), .B2(
        \REGISTERS[9][13] ), .ZN(n36439) );
  AOI22_X1 U1190 ( .A1(n36286), .A2(\REGISTERS[2][13] ), .B1(n36285), .B2(
        \REGISTERS[18][13] ), .ZN(n36438) );
  AOI22_X1 U1191 ( .A1(n36288), .A2(\REGISTERS[3][13] ), .B1(n36287), .B2(
        \REGISTERS[31][13] ), .ZN(n36437) );
  AOI22_X1 U1192 ( .A1(n36290), .A2(\REGISTERS[30][13] ), .B1(n36289), .B2(
        \REGISTERS[8][13] ), .ZN(n36436) );
  NAND4_X1 U1193 ( .A1(n36439), .A2(n36438), .A3(n36437), .A4(n36436), .ZN(
        n36445) );
  AOI22_X1 U1194 ( .A1(n36292), .A2(\REGISTERS[11][13] ), .B1(n36291), .B2(
        \REGISTERS[29][13] ), .ZN(n36443) );
  AOI22_X1 U1195 ( .A1(n36294), .A2(\REGISTERS[1][13] ), .B1(n36293), .B2(
        \REGISTERS[16][13] ), .ZN(n36442) );
  AOI22_X1 U1196 ( .A1(n36296), .A2(\REGISTERS[12][13] ), .B1(n36295), .B2(
        \REGISTERS[24][13] ), .ZN(n36441) );
  AOI22_X1 U1197 ( .A1(n36298), .A2(\REGISTERS[20][13] ), .B1(n36297), .B2(
        \REGISTERS[15][13] ), .ZN(n36440) );
  NAND4_X1 U1198 ( .A1(n36443), .A2(n36442), .A3(n36441), .A4(n36440), .ZN(
        n36444) );
  AOI22_X1 U1199 ( .A1(n36269), .A2(\REGISTERS[5][14] ), .B1(n36268), .B2(
        \REGISTERS[22][14] ), .ZN(n36451) );
  AOI22_X1 U1200 ( .A1(n36271), .A2(\REGISTERS[25][14] ), .B1(n36270), .B2(
        \REGISTERS[21][14] ), .ZN(n36450) );
  AOI22_X1 U1201 ( .A1(n36273), .A2(\REGISTERS[17][14] ), .B1(n36272), .B2(
        \REGISTERS[23][14] ), .ZN(n36449) );
  NAND2_X1 U1202 ( .A1(n36274), .A2(\REGISTERS[19][14] ), .ZN(n36448) );
  NAND4_X1 U1203 ( .A1(n36451), .A2(n36450), .A3(n36449), .A4(n36448), .ZN(
        n36467) );
  AOI22_X1 U1204 ( .A1(n36276), .A2(\REGISTERS[14][14] ), .B1(n36275), .B2(
        \REGISTERS[13][14] ), .ZN(n36455) );
  AOI22_X1 U1205 ( .A1(n36278), .A2(\REGISTERS[27][14] ), .B1(n36277), .B2(
        \REGISTERS[4][14] ), .ZN(n36454) );
  AOI22_X1 U1206 ( .A1(n36280), .A2(\REGISTERS[6][14] ), .B1(n36279), .B2(
        \REGISTERS[28][14] ), .ZN(n36453) );
  AOI22_X1 U1207 ( .A1(n36282), .A2(\REGISTERS[26][14] ), .B1(n36281), .B2(
        \REGISTERS[7][14] ), .ZN(n36452) );
  NAND4_X1 U1208 ( .A1(n36455), .A2(n36454), .A3(n36453), .A4(n36452), .ZN(
        n36466) );
  AOI22_X1 U1209 ( .A1(n36284), .A2(\REGISTERS[10][14] ), .B1(n36283), .B2(
        \REGISTERS[9][14] ), .ZN(n36459) );
  AOI22_X1 U1210 ( .A1(n36286), .A2(\REGISTERS[2][14] ), .B1(n36285), .B2(
        \REGISTERS[18][14] ), .ZN(n36458) );
  AOI22_X1 U1211 ( .A1(n36288), .A2(\REGISTERS[3][14] ), .B1(n36287), .B2(
        \REGISTERS[31][14] ), .ZN(n36457) );
  AOI22_X1 U1212 ( .A1(n36290), .A2(\REGISTERS[30][14] ), .B1(n36289), .B2(
        \REGISTERS[8][14] ), .ZN(n36456) );
  NAND4_X1 U1213 ( .A1(n36459), .A2(n36458), .A3(n36457), .A4(n36456), .ZN(
        n36465) );
  AOI22_X1 U1214 ( .A1(n36292), .A2(\REGISTERS[11][14] ), .B1(n36291), .B2(
        \REGISTERS[29][14] ), .ZN(n36463) );
  AOI22_X1 U1215 ( .A1(n36294), .A2(\REGISTERS[1][14] ), .B1(n36293), .B2(
        \REGISTERS[16][14] ), .ZN(n36462) );
  AOI22_X1 U1216 ( .A1(n36296), .A2(\REGISTERS[12][14] ), .B1(n36295), .B2(
        \REGISTERS[24][14] ), .ZN(n36461) );
  AOI22_X1 U1217 ( .A1(n36298), .A2(\REGISTERS[20][14] ), .B1(n36297), .B2(
        \REGISTERS[15][14] ), .ZN(n36460) );
  NAND4_X1 U1218 ( .A1(n36463), .A2(n36462), .A3(n36461), .A4(n36460), .ZN(
        n36464) );
  AOI22_X1 U1219 ( .A1(n36269), .A2(\REGISTERS[5][15] ), .B1(n36268), .B2(
        \REGISTERS[22][15] ), .ZN(n36471) );
  AOI22_X1 U1220 ( .A1(n36271), .A2(\REGISTERS[25][15] ), .B1(n36270), .B2(
        \REGISTERS[21][15] ), .ZN(n36470) );
  AOI22_X1 U1221 ( .A1(n36273), .A2(\REGISTERS[17][15] ), .B1(n36272), .B2(
        \REGISTERS[23][15] ), .ZN(n36469) );
  NAND2_X1 U1222 ( .A1(n36274), .A2(\REGISTERS[19][15] ), .ZN(n36468) );
  NAND4_X1 U1223 ( .A1(n36471), .A2(n36470), .A3(n36469), .A4(n36468), .ZN(
        n36487) );
  AOI22_X1 U1224 ( .A1(n36276), .A2(\REGISTERS[14][15] ), .B1(n36275), .B2(
        \REGISTERS[13][15] ), .ZN(n36475) );
  AOI22_X1 U1225 ( .A1(n36278), .A2(\REGISTERS[27][15] ), .B1(n36277), .B2(
        \REGISTERS[4][15] ), .ZN(n36474) );
  AOI22_X1 U1226 ( .A1(n36280), .A2(\REGISTERS[6][15] ), .B1(n36279), .B2(
        \REGISTERS[28][15] ), .ZN(n36473) );
  AOI22_X1 U1227 ( .A1(n36282), .A2(\REGISTERS[26][15] ), .B1(n36281), .B2(
        \REGISTERS[7][15] ), .ZN(n36472) );
  NAND4_X1 U1228 ( .A1(n36475), .A2(n36474), .A3(n36473), .A4(n36472), .ZN(
        n36486) );
  AOI22_X1 U1229 ( .A1(n36284), .A2(\REGISTERS[10][15] ), .B1(n36283), .B2(
        \REGISTERS[9][15] ), .ZN(n36479) );
  AOI22_X1 U1230 ( .A1(n36286), .A2(\REGISTERS[2][15] ), .B1(n36285), .B2(
        \REGISTERS[18][15] ), .ZN(n36478) );
  AOI22_X1 U1231 ( .A1(n36288), .A2(\REGISTERS[3][15] ), .B1(n36287), .B2(
        \REGISTERS[31][15] ), .ZN(n36477) );
  AOI22_X1 U1232 ( .A1(n36290), .A2(\REGISTERS[30][15] ), .B1(n36289), .B2(
        \REGISTERS[8][15] ), .ZN(n36476) );
  NAND4_X1 U1233 ( .A1(n36479), .A2(n36478), .A3(n36477), .A4(n36476), .ZN(
        n36485) );
  AOI22_X1 U1234 ( .A1(n36292), .A2(\REGISTERS[11][15] ), .B1(n36291), .B2(
        \REGISTERS[29][15] ), .ZN(n36483) );
  AOI22_X1 U1235 ( .A1(n36294), .A2(\REGISTERS[1][15] ), .B1(n36293), .B2(
        \REGISTERS[16][15] ), .ZN(n36482) );
  AOI22_X1 U1236 ( .A1(n36296), .A2(\REGISTERS[12][15] ), .B1(n36295), .B2(
        \REGISTERS[24][15] ), .ZN(n36481) );
  AOI22_X1 U1237 ( .A1(n36298), .A2(\REGISTERS[20][15] ), .B1(n36297), .B2(
        \REGISTERS[15][15] ), .ZN(n36480) );
  NAND4_X1 U1238 ( .A1(n36483), .A2(n36482), .A3(n36481), .A4(n36480), .ZN(
        n36484) );
  AOI22_X1 U1239 ( .A1(n36278), .A2(\REGISTERS[27][16] ), .B1(n36277), .B2(
        \REGISTERS[4][16] ), .ZN(n36488) );
  AOI22_X1 U1240 ( .A1(n36278), .A2(\REGISTERS[27][17] ), .B1(n36277), .B2(
        \REGISTERS[4][17] ), .ZN(n36489) );
  AOI22_X1 U1241 ( .A1(n36278), .A2(\REGISTERS[27][18] ), .B1(n36277), .B2(
        \REGISTERS[4][18] ), .ZN(n36490) );
  AOI22_X1 U1242 ( .A1(n36278), .A2(\REGISTERS[27][19] ), .B1(n36277), .B2(
        \REGISTERS[4][19] ), .ZN(n36491) );
  AOI22_X1 U1243 ( .A1(n36269), .A2(\REGISTERS[5][1] ), .B1(n36268), .B2(
        \REGISTERS[22][1] ), .ZN(n36495) );
  AOI22_X1 U1244 ( .A1(n36271), .A2(\REGISTERS[25][1] ), .B1(n36270), .B2(
        \REGISTERS[21][1] ), .ZN(n36494) );
  AOI22_X1 U1245 ( .A1(n36273), .A2(\REGISTERS[17][1] ), .B1(n36272), .B2(
        \REGISTERS[23][1] ), .ZN(n36493) );
  NAND2_X1 U1246 ( .A1(n36274), .A2(\REGISTERS[19][1] ), .ZN(n36492) );
  NAND4_X1 U1247 ( .A1(n36495), .A2(n36494), .A3(n36493), .A4(n36492), .ZN(
        n36511) );
  AOI22_X1 U1248 ( .A1(n36276), .A2(\REGISTERS[14][1] ), .B1(n36275), .B2(
        \REGISTERS[13][1] ), .ZN(n36499) );
  AOI22_X1 U1249 ( .A1(n36278), .A2(\REGISTERS[27][1] ), .B1(n36277), .B2(
        \REGISTERS[4][1] ), .ZN(n36498) );
  AOI22_X1 U1250 ( .A1(n36280), .A2(\REGISTERS[6][1] ), .B1(n36279), .B2(
        \REGISTERS[28][1] ), .ZN(n36497) );
  AOI22_X1 U1251 ( .A1(n36282), .A2(\REGISTERS[26][1] ), .B1(n36281), .B2(
        \REGISTERS[7][1] ), .ZN(n36496) );
  NAND4_X1 U1252 ( .A1(n36499), .A2(n36498), .A3(n36497), .A4(n36496), .ZN(
        n36510) );
  AOI22_X1 U1253 ( .A1(n36284), .A2(\REGISTERS[10][1] ), .B1(n36283), .B2(
        \REGISTERS[9][1] ), .ZN(n36503) );
  AOI22_X1 U1254 ( .A1(n36286), .A2(\REGISTERS[2][1] ), .B1(n36285), .B2(
        \REGISTERS[18][1] ), .ZN(n36502) );
  AOI22_X1 U1255 ( .A1(n36288), .A2(\REGISTERS[3][1] ), .B1(n36287), .B2(
        \REGISTERS[31][1] ), .ZN(n36501) );
  AOI22_X1 U1256 ( .A1(n36290), .A2(\REGISTERS[30][1] ), .B1(n36289), .B2(
        \REGISTERS[8][1] ), .ZN(n36500) );
  NAND4_X1 U1257 ( .A1(n36503), .A2(n36502), .A3(n36501), .A4(n36500), .ZN(
        n36509) );
  AOI22_X1 U1258 ( .A1(n36292), .A2(\REGISTERS[11][1] ), .B1(n36291), .B2(
        \REGISTERS[29][1] ), .ZN(n36507) );
  AOI22_X1 U1259 ( .A1(n36294), .A2(\REGISTERS[1][1] ), .B1(n36293), .B2(
        \REGISTERS[16][1] ), .ZN(n36506) );
  AOI22_X1 U1260 ( .A1(n36296), .A2(\REGISTERS[12][1] ), .B1(n36295), .B2(
        \REGISTERS[24][1] ), .ZN(n36505) );
  AOI22_X1 U1261 ( .A1(n36298), .A2(\REGISTERS[20][1] ), .B1(n36297), .B2(
        \REGISTERS[15][1] ), .ZN(n36504) );
  NAND4_X1 U1262 ( .A1(n36507), .A2(n36506), .A3(n36505), .A4(n36504), .ZN(
        n36508) );
  AOI22_X1 U1263 ( .A1(n36278), .A2(\REGISTERS[27][20] ), .B1(n36277), .B2(
        \REGISTERS[4][20] ), .ZN(n36512) );
  AOI22_X1 U1264 ( .A1(n36278), .A2(\REGISTERS[27][21] ), .B1(n36277), .B2(
        \REGISTERS[4][21] ), .ZN(n36513) );
  AOI22_X1 U1265 ( .A1(n36278), .A2(\REGISTERS[27][22] ), .B1(n36277), .B2(
        \REGISTERS[4][22] ), .ZN(n36514) );
  AOI22_X1 U1266 ( .A1(n36278), .A2(\REGISTERS[27][23] ), .B1(n36277), .B2(
        \REGISTERS[4][23] ), .ZN(n36515) );
  AOI22_X1 U1267 ( .A1(n36278), .A2(\REGISTERS[27][24] ), .B1(n36277), .B2(
        \REGISTERS[4][24] ), .ZN(n36516) );
  AOI22_X1 U1268 ( .A1(n36278), .A2(\REGISTERS[27][25] ), .B1(n36277), .B2(
        \REGISTERS[4][25] ), .ZN(n36517) );
  AOI22_X1 U1269 ( .A1(n36269), .A2(\REGISTERS[5][26] ), .B1(n36758), .B2(
        \REGISTERS[22][26] ), .ZN(n36521) );
  AOI22_X1 U1270 ( .A1(n36271), .A2(\REGISTERS[25][26] ), .B1(n36760), .B2(
        \REGISTERS[21][26] ), .ZN(n36520) );
  AOI22_X1 U1271 ( .A1(n36273), .A2(\REGISTERS[17][26] ), .B1(n36762), .B2(
        \REGISTERS[23][26] ), .ZN(n36519) );
  NAND2_X1 U1272 ( .A1(n36274), .A2(\REGISTERS[19][26] ), .ZN(n36518) );
  NAND4_X1 U1273 ( .A1(n36521), .A2(n36520), .A3(n36519), .A4(n36518), .ZN(
        n36537) );
  AOI22_X1 U1274 ( .A1(n36276), .A2(\REGISTERS[14][26] ), .B1(n36275), .B2(
        \REGISTERS[13][26] ), .ZN(n36525) );
  AOI22_X1 U1275 ( .A1(n36772), .A2(\REGISTERS[27][26] ), .B1(n36277), .B2(
        \REGISTERS[4][26] ), .ZN(n36524) );
  AOI22_X1 U1276 ( .A1(n36280), .A2(\REGISTERS[6][26] ), .B1(n36279), .B2(
        \REGISTERS[28][26] ), .ZN(n36523) );
  AOI22_X1 U1277 ( .A1(n36282), .A2(\REGISTERS[26][26] ), .B1(n36775), .B2(
        \REGISTERS[7][26] ), .ZN(n36522) );
  NAND4_X1 U1278 ( .A1(n36525), .A2(n36524), .A3(n36523), .A4(n36522), .ZN(
        n36536) );
  AOI22_X1 U1279 ( .A1(n36284), .A2(\REGISTERS[10][26] ), .B1(n36283), .B2(
        \REGISTERS[9][26] ), .ZN(n36529) );
  AOI22_X1 U1280 ( .A1(n36286), .A2(\REGISTERS[2][26] ), .B1(n36783), .B2(
        \REGISTERS[18][26] ), .ZN(n36528) );
  AOI22_X1 U1281 ( .A1(n36288), .A2(\REGISTERS[3][26] ), .B1(n36785), .B2(
        \REGISTERS[31][26] ), .ZN(n36527) );
  AOI22_X1 U1282 ( .A1(n36290), .A2(\REGISTERS[30][26] ), .B1(n36289), .B2(
        \REGISTERS[8][26] ), .ZN(n36526) );
  NAND4_X1 U1283 ( .A1(n36529), .A2(n36528), .A3(n36527), .A4(n36526), .ZN(
        n36535) );
  AOI22_X1 U1284 ( .A1(n36292), .A2(\REGISTERS[11][26] ), .B1(n36291), .B2(
        \REGISTERS[29][26] ), .ZN(n36533) );
  AOI22_X1 U1285 ( .A1(n36294), .A2(\REGISTERS[1][26] ), .B1(n36293), .B2(
        \REGISTERS[16][26] ), .ZN(n36532) );
  AOI22_X1 U1286 ( .A1(n36296), .A2(\REGISTERS[12][26] ), .B1(n36295), .B2(
        \REGISTERS[24][26] ), .ZN(n36531) );
  AOI22_X1 U1287 ( .A1(n36298), .A2(\REGISTERS[20][26] ), .B1(n36297), .B2(
        \REGISTERS[15][26] ), .ZN(n36530) );
  NAND4_X1 U1288 ( .A1(n36533), .A2(n36532), .A3(n36531), .A4(n36530), .ZN(
        n36534) );
  AOI22_X1 U1289 ( .A1(n36759), .A2(\REGISTERS[5][27] ), .B1(n36758), .B2(
        \REGISTERS[22][27] ), .ZN(n36541) );
  AOI22_X1 U1290 ( .A1(n36761), .A2(\REGISTERS[25][27] ), .B1(n36760), .B2(
        \REGISTERS[21][27] ), .ZN(n36540) );
  AOI22_X1 U1291 ( .A1(n36763), .A2(\REGISTERS[17][27] ), .B1(n36762), .B2(
        \REGISTERS[23][27] ), .ZN(n36539) );
  NAND2_X1 U1292 ( .A1(n36764), .A2(\REGISTERS[19][27] ), .ZN(n36538) );
  NAND4_X1 U1293 ( .A1(n36541), .A2(n36540), .A3(n36539), .A4(n36538), .ZN(
        n36557) );
  AOI22_X1 U1294 ( .A1(n36770), .A2(\REGISTERS[14][27] ), .B1(n36769), .B2(
        \REGISTERS[13][27] ), .ZN(n36545) );
  AOI22_X1 U1295 ( .A1(n36278), .A2(\REGISTERS[27][27] ), .B1(n36277), .B2(
        \REGISTERS[4][27] ), .ZN(n36544) );
  AOI22_X1 U1296 ( .A1(n36774), .A2(\REGISTERS[6][27] ), .B1(n36773), .B2(
        \REGISTERS[28][27] ), .ZN(n36543) );
  AOI22_X1 U1297 ( .A1(n36776), .A2(\REGISTERS[26][27] ), .B1(n36775), .B2(
        \REGISTERS[7][27] ), .ZN(n36542) );
  NAND4_X1 U1298 ( .A1(n36545), .A2(n36544), .A3(n36543), .A4(n36542), .ZN(
        n36556) );
  AOI22_X1 U1299 ( .A1(n36782), .A2(\REGISTERS[10][27] ), .B1(n36781), .B2(
        \REGISTERS[9][27] ), .ZN(n36549) );
  AOI22_X1 U1300 ( .A1(n36286), .A2(\REGISTERS[2][27] ), .B1(n36783), .B2(
        \REGISTERS[18][27] ), .ZN(n36548) );
  AOI22_X1 U1301 ( .A1(n36786), .A2(\REGISTERS[3][27] ), .B1(n36785), .B2(
        \REGISTERS[31][27] ), .ZN(n36547) );
  AOI22_X1 U1302 ( .A1(n36788), .A2(\REGISTERS[30][27] ), .B1(n36787), .B2(
        \REGISTERS[8][27] ), .ZN(n36546) );
  NAND4_X1 U1303 ( .A1(n36549), .A2(n36548), .A3(n36547), .A4(n36546), .ZN(
        n36555) );
  AOI22_X1 U1304 ( .A1(n36292), .A2(\REGISTERS[11][27] ), .B1(n36793), .B2(
        \REGISTERS[29][27] ), .ZN(n36553) );
  AOI22_X1 U1305 ( .A1(n36294), .A2(\REGISTERS[1][27] ), .B1(n36795), .B2(
        \REGISTERS[16][27] ), .ZN(n36552) );
  AOI22_X1 U1306 ( .A1(n36296), .A2(\REGISTERS[12][27] ), .B1(n36797), .B2(
        \REGISTERS[24][27] ), .ZN(n36551) );
  AOI22_X1 U1307 ( .A1(n36800), .A2(\REGISTERS[20][27] ), .B1(n36799), .B2(
        \REGISTERS[15][27] ), .ZN(n36550) );
  NAND4_X1 U1308 ( .A1(n36553), .A2(n36552), .A3(n36551), .A4(n36550), .ZN(
        n36554) );
  AOI22_X1 U1309 ( .A1(n36759), .A2(\REGISTERS[5][28] ), .B1(n36758), .B2(
        \REGISTERS[22][28] ), .ZN(n36561) );
  AOI22_X1 U1310 ( .A1(n36761), .A2(\REGISTERS[25][28] ), .B1(n36270), .B2(
        \REGISTERS[21][28] ), .ZN(n36560) );
  AOI22_X1 U1311 ( .A1(n36763), .A2(\REGISTERS[17][28] ), .B1(n36762), .B2(
        \REGISTERS[23][28] ), .ZN(n36559) );
  NAND2_X1 U1312 ( .A1(n36764), .A2(\REGISTERS[19][28] ), .ZN(n36558) );
  NAND4_X1 U1313 ( .A1(n36561), .A2(n36560), .A3(n36559), .A4(n36558), .ZN(
        n36577) );
  AOI22_X1 U1314 ( .A1(n36276), .A2(\REGISTERS[14][28] ), .B1(n36769), .B2(
        \REGISTERS[13][28] ), .ZN(n36565) );
  AOI22_X1 U1315 ( .A1(n36772), .A2(\REGISTERS[27][28] ), .B1(n36277), .B2(
        \REGISTERS[4][28] ), .ZN(n36564) );
  AOI22_X1 U1316 ( .A1(n36280), .A2(\REGISTERS[6][28] ), .B1(n36773), .B2(
        \REGISTERS[28][28] ), .ZN(n36563) );
  AOI22_X1 U1317 ( .A1(n36282), .A2(\REGISTERS[26][28] ), .B1(n36281), .B2(
        \REGISTERS[7][28] ), .ZN(n36562) );
  NAND4_X1 U1318 ( .A1(n36565), .A2(n36564), .A3(n36563), .A4(n36562), .ZN(
        n36576) );
  AOI22_X1 U1319 ( .A1(n36284), .A2(\REGISTERS[10][28] ), .B1(n36781), .B2(
        \REGISTERS[9][28] ), .ZN(n36569) );
  AOI22_X1 U1320 ( .A1(n36286), .A2(\REGISTERS[2][28] ), .B1(n36783), .B2(
        \REGISTERS[18][28] ), .ZN(n36568) );
  AOI22_X1 U1321 ( .A1(n36288), .A2(\REGISTERS[3][28] ), .B1(n36785), .B2(
        \REGISTERS[31][28] ), .ZN(n36567) );
  AOI22_X1 U1322 ( .A1(n36290), .A2(\REGISTERS[30][28] ), .B1(n36787), .B2(
        \REGISTERS[8][28] ), .ZN(n36566) );
  NAND4_X1 U1323 ( .A1(n36569), .A2(n36568), .A3(n36567), .A4(n36566), .ZN(
        n36575) );
  AOI22_X1 U1324 ( .A1(n36794), .A2(\REGISTERS[11][28] ), .B1(n36793), .B2(
        \REGISTERS[29][28] ), .ZN(n36573) );
  AOI22_X1 U1325 ( .A1(n36796), .A2(\REGISTERS[1][28] ), .B1(n36795), .B2(
        \REGISTERS[16][28] ), .ZN(n36572) );
  AOI22_X1 U1326 ( .A1(n36798), .A2(\REGISTERS[12][28] ), .B1(n36797), .B2(
        \REGISTERS[24][28] ), .ZN(n36571) );
  AOI22_X1 U1327 ( .A1(n36298), .A2(\REGISTERS[20][28] ), .B1(n36799), .B2(
        \REGISTERS[15][28] ), .ZN(n36570) );
  NAND4_X1 U1328 ( .A1(n36573), .A2(n36572), .A3(n36571), .A4(n36570), .ZN(
        n36574) );
  AOI22_X1 U1329 ( .A1(n36759), .A2(\REGISTERS[5][29] ), .B1(n36758), .B2(
        \REGISTERS[22][29] ), .ZN(n36581) );
  AOI22_X1 U1330 ( .A1(n36761), .A2(\REGISTERS[25][29] ), .B1(n36760), .B2(
        \REGISTERS[21][29] ), .ZN(n36580) );
  AOI22_X1 U1331 ( .A1(n36763), .A2(\REGISTERS[17][29] ), .B1(n36762), .B2(
        \REGISTERS[23][29] ), .ZN(n36579) );
  NAND2_X1 U1332 ( .A1(n36764), .A2(\REGISTERS[19][29] ), .ZN(n36578) );
  NAND4_X1 U1333 ( .A1(n36581), .A2(n36580), .A3(n36579), .A4(n36578), .ZN(
        n36597) );
  AOI22_X1 U1334 ( .A1(n36770), .A2(\REGISTERS[14][29] ), .B1(n36769), .B2(
        \REGISTERS[13][29] ), .ZN(n36585) );
  AOI22_X1 U1335 ( .A1(n36772), .A2(\REGISTERS[27][29] ), .B1(n36277), .B2(
        \REGISTERS[4][29] ), .ZN(n36584) );
  AOI22_X1 U1336 ( .A1(n36774), .A2(\REGISTERS[6][29] ), .B1(n36773), .B2(
        \REGISTERS[28][29] ), .ZN(n36583) );
  AOI22_X1 U1337 ( .A1(n36776), .A2(\REGISTERS[26][29] ), .B1(n36775), .B2(
        \REGISTERS[7][29] ), .ZN(n36582) );
  NAND4_X1 U1338 ( .A1(n36585), .A2(n36584), .A3(n36583), .A4(n36582), .ZN(
        n36596) );
  AOI22_X1 U1339 ( .A1(n36782), .A2(\REGISTERS[10][29] ), .B1(n36781), .B2(
        \REGISTERS[9][29] ), .ZN(n36589) );
  AOI22_X1 U1340 ( .A1(n36286), .A2(\REGISTERS[2][29] ), .B1(n36783), .B2(
        \REGISTERS[18][29] ), .ZN(n36588) );
  AOI22_X1 U1341 ( .A1(n36786), .A2(\REGISTERS[3][29] ), .B1(n36785), .B2(
        \REGISTERS[31][29] ), .ZN(n36587) );
  AOI22_X1 U1342 ( .A1(n36788), .A2(\REGISTERS[30][29] ), .B1(n36787), .B2(
        \REGISTERS[8][29] ), .ZN(n36586) );
  NAND4_X1 U1343 ( .A1(n36589), .A2(n36588), .A3(n36587), .A4(n36586), .ZN(
        n36595) );
  AOI22_X1 U1344 ( .A1(n36794), .A2(\REGISTERS[11][29] ), .B1(n36793), .B2(
        \REGISTERS[29][29] ), .ZN(n36593) );
  AOI22_X1 U1345 ( .A1(n36796), .A2(\REGISTERS[1][29] ), .B1(n36795), .B2(
        \REGISTERS[16][29] ), .ZN(n36592) );
  AOI22_X1 U1346 ( .A1(n36798), .A2(\REGISTERS[12][29] ), .B1(n36797), .B2(
        \REGISTERS[24][29] ), .ZN(n36591) );
  AOI22_X1 U1347 ( .A1(n36800), .A2(\REGISTERS[20][29] ), .B1(n36799), .B2(
        \REGISTERS[15][29] ), .ZN(n36590) );
  NAND4_X1 U1348 ( .A1(n36593), .A2(n36592), .A3(n36591), .A4(n36590), .ZN(
        n36594) );
  AOI22_X1 U1349 ( .A1(n36759), .A2(\REGISTERS[5][2] ), .B1(n36758), .B2(
        \REGISTERS[22][2] ), .ZN(n36601) );
  AOI22_X1 U1350 ( .A1(n36761), .A2(\REGISTERS[25][2] ), .B1(n36760), .B2(
        \REGISTERS[21][2] ), .ZN(n36600) );
  AOI22_X1 U1351 ( .A1(n36763), .A2(\REGISTERS[17][2] ), .B1(n36762), .B2(
        \REGISTERS[23][2] ), .ZN(n36599) );
  NAND2_X1 U1352 ( .A1(n36764), .A2(\REGISTERS[19][2] ), .ZN(n36598) );
  NAND4_X1 U1353 ( .A1(n36601), .A2(n36600), .A3(n36599), .A4(n36598), .ZN(
        n36617) );
  AOI22_X1 U1354 ( .A1(n36770), .A2(\REGISTERS[14][2] ), .B1(n36769), .B2(
        \REGISTERS[13][2] ), .ZN(n36605) );
  AOI22_X1 U1355 ( .A1(n36772), .A2(\REGISTERS[27][2] ), .B1(n36277), .B2(
        \REGISTERS[4][2] ), .ZN(n36604) );
  AOI22_X1 U1356 ( .A1(n36774), .A2(\REGISTERS[6][2] ), .B1(n36773), .B2(
        \REGISTERS[28][2] ), .ZN(n36603) );
  AOI22_X1 U1357 ( .A1(n36776), .A2(\REGISTERS[26][2] ), .B1(n36775), .B2(
        \REGISTERS[7][2] ), .ZN(n36602) );
  NAND4_X1 U1358 ( .A1(n36605), .A2(n36604), .A3(n36603), .A4(n36602), .ZN(
        n36616) );
  AOI22_X1 U1359 ( .A1(n36782), .A2(\REGISTERS[10][2] ), .B1(n36781), .B2(
        \REGISTERS[9][2] ), .ZN(n36609) );
  AOI22_X1 U1360 ( .A1(n36286), .A2(\REGISTERS[2][2] ), .B1(n36783), .B2(
        \REGISTERS[18][2] ), .ZN(n36608) );
  AOI22_X1 U1361 ( .A1(n36786), .A2(\REGISTERS[3][2] ), .B1(n36785), .B2(
        \REGISTERS[31][2] ), .ZN(n36607) );
  AOI22_X1 U1362 ( .A1(n36788), .A2(\REGISTERS[30][2] ), .B1(n36787), .B2(
        \REGISTERS[8][2] ), .ZN(n36606) );
  NAND4_X1 U1363 ( .A1(n36609), .A2(n36608), .A3(n36607), .A4(n36606), .ZN(
        n36615) );
  AOI22_X1 U1364 ( .A1(n36794), .A2(\REGISTERS[11][2] ), .B1(n36793), .B2(
        \REGISTERS[29][2] ), .ZN(n36613) );
  AOI22_X1 U1365 ( .A1(n36796), .A2(\REGISTERS[1][2] ), .B1(n36795), .B2(
        \REGISTERS[16][2] ), .ZN(n36612) );
  AOI22_X1 U1366 ( .A1(n36798), .A2(\REGISTERS[12][2] ), .B1(n36797), .B2(
        \REGISTERS[24][2] ), .ZN(n36611) );
  AOI22_X1 U1367 ( .A1(n36800), .A2(\REGISTERS[20][2] ), .B1(n36799), .B2(
        \REGISTERS[15][2] ), .ZN(n36610) );
  NAND4_X1 U1368 ( .A1(n36613), .A2(n36612), .A3(n36611), .A4(n36610), .ZN(
        n36614) );
  AOI22_X1 U1369 ( .A1(n36269), .A2(\REGISTERS[5][30] ), .B1(n36758), .B2(
        \REGISTERS[22][30] ), .ZN(n36621) );
  AOI22_X1 U1370 ( .A1(n36271), .A2(\REGISTERS[25][30] ), .B1(n36760), .B2(
        \REGISTERS[21][30] ), .ZN(n36620) );
  AOI22_X1 U1371 ( .A1(n36273), .A2(\REGISTERS[17][30] ), .B1(n36272), .B2(
        \REGISTERS[23][30] ), .ZN(n36619) );
  NAND2_X1 U1372 ( .A1(n36764), .A2(\REGISTERS[19][30] ), .ZN(n36618) );
  NAND4_X1 U1373 ( .A1(n36621), .A2(n36620), .A3(n36619), .A4(n36618), .ZN(
        n36637) );
  AOI22_X1 U1374 ( .A1(n36770), .A2(\REGISTERS[14][30] ), .B1(n36769), .B2(
        \REGISTERS[13][30] ), .ZN(n36625) );
  AOI22_X1 U1375 ( .A1(n36278), .A2(\REGISTERS[27][30] ), .B1(n36771), .B2(
        \REGISTERS[4][30] ), .ZN(n36624) );
  AOI22_X1 U1376 ( .A1(n36774), .A2(\REGISTERS[6][30] ), .B1(n36773), .B2(
        \REGISTERS[28][30] ), .ZN(n36623) );
  AOI22_X1 U1377 ( .A1(n36776), .A2(\REGISTERS[26][30] ), .B1(n36775), .B2(
        \REGISTERS[7][30] ), .ZN(n36622) );
  NAND4_X1 U1378 ( .A1(n36625), .A2(n36624), .A3(n36623), .A4(n36622), .ZN(
        n36636) );
  AOI22_X1 U1379 ( .A1(n36782), .A2(\REGISTERS[10][30] ), .B1(n36781), .B2(
        \REGISTERS[9][30] ), .ZN(n36629) );
  AOI22_X1 U1380 ( .A1(n36784), .A2(\REGISTERS[2][30] ), .B1(n36783), .B2(
        \REGISTERS[18][30] ), .ZN(n36628) );
  AOI22_X1 U1381 ( .A1(n36786), .A2(\REGISTERS[3][30] ), .B1(n36785), .B2(
        \REGISTERS[31][30] ), .ZN(n36627) );
  AOI22_X1 U1382 ( .A1(n36788), .A2(\REGISTERS[30][30] ), .B1(n36787), .B2(
        \REGISTERS[8][30] ), .ZN(n36626) );
  NAND4_X1 U1383 ( .A1(n36629), .A2(n36628), .A3(n36627), .A4(n36626), .ZN(
        n36635) );
  AOI22_X1 U1384 ( .A1(n36794), .A2(\REGISTERS[11][30] ), .B1(n36793), .B2(
        \REGISTERS[29][30] ), .ZN(n36633) );
  AOI22_X1 U1385 ( .A1(n36796), .A2(\REGISTERS[1][30] ), .B1(n36795), .B2(
        \REGISTERS[16][30] ), .ZN(n36632) );
  AOI22_X1 U1386 ( .A1(n36798), .A2(\REGISTERS[12][30] ), .B1(n36797), .B2(
        \REGISTERS[24][30] ), .ZN(n36631) );
  AOI22_X1 U1387 ( .A1(n36800), .A2(\REGISTERS[20][30] ), .B1(n36799), .B2(
        \REGISTERS[15][30] ), .ZN(n36630) );
  NAND4_X1 U1388 ( .A1(n36633), .A2(n36632), .A3(n36631), .A4(n36630), .ZN(
        n36634) );
  AOI22_X1 U1389 ( .A1(n36759), .A2(\REGISTERS[5][3] ), .B1(n36758), .B2(
        \REGISTERS[22][3] ), .ZN(n36641) );
  AOI22_X1 U1390 ( .A1(n36761), .A2(\REGISTERS[25][3] ), .B1(n36760), .B2(
        \REGISTERS[21][3] ), .ZN(n36640) );
  AOI22_X1 U1391 ( .A1(n36763), .A2(\REGISTERS[17][3] ), .B1(n36762), .B2(
        \REGISTERS[23][3] ), .ZN(n36639) );
  NAND2_X1 U1392 ( .A1(n36764), .A2(\REGISTERS[19][3] ), .ZN(n36638) );
  NAND4_X1 U1393 ( .A1(n36641), .A2(n36640), .A3(n36639), .A4(n36638), .ZN(
        n36657) );
  AOI22_X1 U1394 ( .A1(n36770), .A2(\REGISTERS[14][3] ), .B1(n36769), .B2(
        \REGISTERS[13][3] ), .ZN(n36645) );
  AOI22_X1 U1395 ( .A1(n36772), .A2(\REGISTERS[27][3] ), .B1(n36771), .B2(
        \REGISTERS[4][3] ), .ZN(n36644) );
  AOI22_X1 U1396 ( .A1(n36774), .A2(\REGISTERS[6][3] ), .B1(n36773), .B2(
        \REGISTERS[28][3] ), .ZN(n36643) );
  AOI22_X1 U1397 ( .A1(n36776), .A2(\REGISTERS[26][3] ), .B1(n36775), .B2(
        \REGISTERS[7][3] ), .ZN(n36642) );
  NAND4_X1 U1398 ( .A1(n36645), .A2(n36644), .A3(n36643), .A4(n36642), .ZN(
        n36656) );
  AOI22_X1 U1399 ( .A1(n36782), .A2(\REGISTERS[10][3] ), .B1(n36781), .B2(
        \REGISTERS[9][3] ), .ZN(n36649) );
  AOI22_X1 U1400 ( .A1(n36784), .A2(\REGISTERS[2][3] ), .B1(n36783), .B2(
        \REGISTERS[18][3] ), .ZN(n36648) );
  AOI22_X1 U1401 ( .A1(n36786), .A2(\REGISTERS[3][3] ), .B1(n36785), .B2(
        \REGISTERS[31][3] ), .ZN(n36647) );
  AOI22_X1 U1402 ( .A1(n36788), .A2(\REGISTERS[30][3] ), .B1(n36787), .B2(
        \REGISTERS[8][3] ), .ZN(n36646) );
  NAND4_X1 U1403 ( .A1(n36649), .A2(n36648), .A3(n36647), .A4(n36646), .ZN(
        n36655) );
  AOI22_X1 U1404 ( .A1(n36794), .A2(\REGISTERS[11][3] ), .B1(n36793), .B2(
        \REGISTERS[29][3] ), .ZN(n36653) );
  AOI22_X1 U1405 ( .A1(n36796), .A2(\REGISTERS[1][3] ), .B1(n36795), .B2(
        \REGISTERS[16][3] ), .ZN(n36652) );
  AOI22_X1 U1406 ( .A1(n36798), .A2(\REGISTERS[12][3] ), .B1(n36797), .B2(
        \REGISTERS[24][3] ), .ZN(n36651) );
  AOI22_X1 U1407 ( .A1(n36800), .A2(\REGISTERS[20][3] ), .B1(n36799), .B2(
        \REGISTERS[15][3] ), .ZN(n36650) );
  NAND4_X1 U1408 ( .A1(n36653), .A2(n36652), .A3(n36651), .A4(n36650), .ZN(
        n36654) );
  AOI22_X1 U1409 ( .A1(n36759), .A2(\REGISTERS[5][4] ), .B1(n36758), .B2(
        \REGISTERS[22][4] ), .ZN(n36661) );
  AOI22_X1 U1410 ( .A1(n36761), .A2(\REGISTERS[25][4] ), .B1(n36760), .B2(
        \REGISTERS[21][4] ), .ZN(n36660) );
  AOI22_X1 U1411 ( .A1(n36763), .A2(\REGISTERS[17][4] ), .B1(n36762), .B2(
        \REGISTERS[23][4] ), .ZN(n36659) );
  NAND2_X1 U1412 ( .A1(n36764), .A2(\REGISTERS[19][4] ), .ZN(n36658) );
  NAND4_X1 U1413 ( .A1(n36661), .A2(n36660), .A3(n36659), .A4(n36658), .ZN(
        n36677) );
  AOI22_X1 U1414 ( .A1(n36770), .A2(\REGISTERS[14][4] ), .B1(n36769), .B2(
        \REGISTERS[13][4] ), .ZN(n36665) );
  AOI22_X1 U1415 ( .A1(n36772), .A2(\REGISTERS[27][4] ), .B1(n36771), .B2(
        \REGISTERS[4][4] ), .ZN(n36664) );
  AOI22_X1 U1416 ( .A1(n36774), .A2(\REGISTERS[6][4] ), .B1(n36773), .B2(
        \REGISTERS[28][4] ), .ZN(n36663) );
  AOI22_X1 U1417 ( .A1(n36776), .A2(\REGISTERS[26][4] ), .B1(n36775), .B2(
        \REGISTERS[7][4] ), .ZN(n36662) );
  NAND4_X1 U1418 ( .A1(n36665), .A2(n36664), .A3(n36663), .A4(n36662), .ZN(
        n36676) );
  AOI22_X1 U1419 ( .A1(n36782), .A2(\REGISTERS[10][4] ), .B1(n36781), .B2(
        \REGISTERS[9][4] ), .ZN(n36669) );
  AOI22_X1 U1420 ( .A1(n36784), .A2(\REGISTERS[2][4] ), .B1(n36783), .B2(
        \REGISTERS[18][4] ), .ZN(n36668) );
  AOI22_X1 U1421 ( .A1(n36786), .A2(\REGISTERS[3][4] ), .B1(n36785), .B2(
        \REGISTERS[31][4] ), .ZN(n36667) );
  AOI22_X1 U1422 ( .A1(n36788), .A2(\REGISTERS[30][4] ), .B1(n36787), .B2(
        \REGISTERS[8][4] ), .ZN(n36666) );
  NAND4_X1 U1423 ( .A1(n36669), .A2(n36668), .A3(n36667), .A4(n36666), .ZN(
        n36675) );
  AOI22_X1 U1424 ( .A1(n36794), .A2(\REGISTERS[11][4] ), .B1(n36793), .B2(
        \REGISTERS[29][4] ), .ZN(n36673) );
  AOI22_X1 U1425 ( .A1(n36796), .A2(\REGISTERS[1][4] ), .B1(n36795), .B2(
        \REGISTERS[16][4] ), .ZN(n36672) );
  AOI22_X1 U1426 ( .A1(n36798), .A2(\REGISTERS[12][4] ), .B1(n36797), .B2(
        \REGISTERS[24][4] ), .ZN(n36671) );
  AOI22_X1 U1427 ( .A1(n36800), .A2(\REGISTERS[20][4] ), .B1(n36799), .B2(
        \REGISTERS[15][4] ), .ZN(n36670) );
  NAND4_X1 U1428 ( .A1(n36673), .A2(n36672), .A3(n36671), .A4(n36670), .ZN(
        n36674) );
  AOI22_X1 U1429 ( .A1(n36759), .A2(\REGISTERS[5][5] ), .B1(n36758), .B2(
        \REGISTERS[22][5] ), .ZN(n36681) );
  AOI22_X1 U1430 ( .A1(n36761), .A2(\REGISTERS[25][5] ), .B1(n36760), .B2(
        \REGISTERS[21][5] ), .ZN(n36680) );
  AOI22_X1 U1431 ( .A1(n36763), .A2(\REGISTERS[17][5] ), .B1(n36762), .B2(
        \REGISTERS[23][5] ), .ZN(n36679) );
  NAND2_X1 U1432 ( .A1(n36764), .A2(\REGISTERS[19][5] ), .ZN(n36678) );
  NAND4_X1 U1433 ( .A1(n36681), .A2(n36680), .A3(n36679), .A4(n36678), .ZN(
        n36697) );
  AOI22_X1 U1434 ( .A1(n36770), .A2(\REGISTERS[14][5] ), .B1(n36769), .B2(
        \REGISTERS[13][5] ), .ZN(n36685) );
  AOI22_X1 U1435 ( .A1(n36772), .A2(\REGISTERS[27][5] ), .B1(n36771), .B2(
        \REGISTERS[4][5] ), .ZN(n36684) );
  AOI22_X1 U1436 ( .A1(n36774), .A2(\REGISTERS[6][5] ), .B1(n36773), .B2(
        \REGISTERS[28][5] ), .ZN(n36683) );
  AOI22_X1 U1437 ( .A1(n36776), .A2(\REGISTERS[26][5] ), .B1(n36775), .B2(
        \REGISTERS[7][5] ), .ZN(n36682) );
  NAND4_X1 U1438 ( .A1(n36685), .A2(n36684), .A3(n36683), .A4(n36682), .ZN(
        n36696) );
  AOI22_X1 U1439 ( .A1(n36782), .A2(\REGISTERS[10][5] ), .B1(n36781), .B2(
        \REGISTERS[9][5] ), .ZN(n36689) );
  AOI22_X1 U1440 ( .A1(n36784), .A2(\REGISTERS[2][5] ), .B1(n36783), .B2(
        \REGISTERS[18][5] ), .ZN(n36688) );
  AOI22_X1 U1441 ( .A1(n36786), .A2(\REGISTERS[3][5] ), .B1(n36785), .B2(
        \REGISTERS[31][5] ), .ZN(n36687) );
  AOI22_X1 U1442 ( .A1(n36788), .A2(\REGISTERS[30][5] ), .B1(n36787), .B2(
        \REGISTERS[8][5] ), .ZN(n36686) );
  NAND4_X1 U1443 ( .A1(n36689), .A2(n36688), .A3(n36687), .A4(n36686), .ZN(
        n36695) );
  AOI22_X1 U1444 ( .A1(n36794), .A2(\REGISTERS[11][5] ), .B1(n36793), .B2(
        \REGISTERS[29][5] ), .ZN(n36693) );
  AOI22_X1 U1445 ( .A1(n36796), .A2(\REGISTERS[1][5] ), .B1(n36795), .B2(
        \REGISTERS[16][5] ), .ZN(n36692) );
  AOI22_X1 U1446 ( .A1(n36798), .A2(\REGISTERS[12][5] ), .B1(n36797), .B2(
        \REGISTERS[24][5] ), .ZN(n36691) );
  AOI22_X1 U1447 ( .A1(n36800), .A2(\REGISTERS[20][5] ), .B1(n36799), .B2(
        \REGISTERS[15][5] ), .ZN(n36690) );
  NAND4_X1 U1448 ( .A1(n36693), .A2(n36692), .A3(n36691), .A4(n36690), .ZN(
        n36694) );
  AOI22_X1 U1449 ( .A1(n36759), .A2(\REGISTERS[5][6] ), .B1(n36758), .B2(
        \REGISTERS[22][6] ), .ZN(n36701) );
  AOI22_X1 U1450 ( .A1(n36761), .A2(\REGISTERS[25][6] ), .B1(n36760), .B2(
        \REGISTERS[21][6] ), .ZN(n36700) );
  AOI22_X1 U1451 ( .A1(n36763), .A2(\REGISTERS[17][6] ), .B1(n36762), .B2(
        \REGISTERS[23][6] ), .ZN(n36699) );
  NAND2_X1 U1452 ( .A1(n36764), .A2(\REGISTERS[19][6] ), .ZN(n36698) );
  NAND4_X1 U1453 ( .A1(n36701), .A2(n36700), .A3(n36699), .A4(n36698), .ZN(
        n36717) );
  AOI22_X1 U1454 ( .A1(n36770), .A2(\REGISTERS[14][6] ), .B1(n36769), .B2(
        \REGISTERS[13][6] ), .ZN(n36705) );
  AOI22_X1 U1455 ( .A1(n36772), .A2(\REGISTERS[27][6] ), .B1(n36771), .B2(
        \REGISTERS[4][6] ), .ZN(n36704) );
  AOI22_X1 U1456 ( .A1(n36774), .A2(\REGISTERS[6][6] ), .B1(n36773), .B2(
        \REGISTERS[28][6] ), .ZN(n36703) );
  AOI22_X1 U1457 ( .A1(n36776), .A2(\REGISTERS[26][6] ), .B1(n36775), .B2(
        \REGISTERS[7][6] ), .ZN(n36702) );
  NAND4_X1 U1458 ( .A1(n36705), .A2(n36704), .A3(n36703), .A4(n36702), .ZN(
        n36716) );
  AOI22_X1 U1459 ( .A1(n36782), .A2(\REGISTERS[10][6] ), .B1(n36781), .B2(
        \REGISTERS[9][6] ), .ZN(n36709) );
  AOI22_X1 U1460 ( .A1(n36784), .A2(\REGISTERS[2][6] ), .B1(n36783), .B2(
        \REGISTERS[18][6] ), .ZN(n36708) );
  AOI22_X1 U1461 ( .A1(n36786), .A2(\REGISTERS[3][6] ), .B1(n36785), .B2(
        \REGISTERS[31][6] ), .ZN(n36707) );
  AOI22_X1 U1462 ( .A1(n36788), .A2(\REGISTERS[30][6] ), .B1(n36787), .B2(
        \REGISTERS[8][6] ), .ZN(n36706) );
  NAND4_X1 U1463 ( .A1(n36709), .A2(n36708), .A3(n36707), .A4(n36706), .ZN(
        n36715) );
  AOI22_X1 U1464 ( .A1(n36794), .A2(\REGISTERS[11][6] ), .B1(n36793), .B2(
        \REGISTERS[29][6] ), .ZN(n36713) );
  AOI22_X1 U1465 ( .A1(n36796), .A2(\REGISTERS[1][6] ), .B1(n36795), .B2(
        \REGISTERS[16][6] ), .ZN(n36712) );
  AOI22_X1 U1466 ( .A1(n36798), .A2(\REGISTERS[12][6] ), .B1(n36797), .B2(
        \REGISTERS[24][6] ), .ZN(n36711) );
  AOI22_X1 U1467 ( .A1(n36800), .A2(\REGISTERS[20][6] ), .B1(n36799), .B2(
        \REGISTERS[15][6] ), .ZN(n36710) );
  NAND4_X1 U1468 ( .A1(n36713), .A2(n36712), .A3(n36711), .A4(n36710), .ZN(
        n36714) );
  AOI22_X1 U1469 ( .A1(n36269), .A2(\REGISTERS[5][7] ), .B1(n36268), .B2(
        \REGISTERS[22][7] ), .ZN(n36721) );
  AOI22_X1 U1470 ( .A1(n36271), .A2(\REGISTERS[25][7] ), .B1(n36270), .B2(
        \REGISTERS[21][7] ), .ZN(n36720) );
  AOI22_X1 U1471 ( .A1(n36273), .A2(\REGISTERS[17][7] ), .B1(n36272), .B2(
        \REGISTERS[23][7] ), .ZN(n36719) );
  NAND2_X1 U1472 ( .A1(n36764), .A2(\REGISTERS[19][7] ), .ZN(n36718) );
  NAND4_X1 U1473 ( .A1(n36721), .A2(n36720), .A3(n36719), .A4(n36718), .ZN(
        n36737) );
  AOI22_X1 U1474 ( .A1(n36276), .A2(\REGISTERS[14][7] ), .B1(n36275), .B2(
        \REGISTERS[13][7] ), .ZN(n36725) );
  AOI22_X1 U1475 ( .A1(n36278), .A2(\REGISTERS[27][7] ), .B1(n36277), .B2(
        \REGISTERS[4][7] ), .ZN(n36724) );
  AOI22_X1 U1476 ( .A1(n36280), .A2(\REGISTERS[6][7] ), .B1(n36279), .B2(
        \REGISTERS[28][7] ), .ZN(n36723) );
  AOI22_X1 U1477 ( .A1(n36282), .A2(\REGISTERS[26][7] ), .B1(n36281), .B2(
        \REGISTERS[7][7] ), .ZN(n36722) );
  NAND4_X1 U1478 ( .A1(n36725), .A2(n36724), .A3(n36723), .A4(n36722), .ZN(
        n36736) );
  AOI22_X1 U1479 ( .A1(n36284), .A2(\REGISTERS[10][7] ), .B1(n36283), .B2(
        \REGISTERS[9][7] ), .ZN(n36729) );
  AOI22_X1 U1480 ( .A1(n36286), .A2(\REGISTERS[2][7] ), .B1(n36285), .B2(
        \REGISTERS[18][7] ), .ZN(n36728) );
  AOI22_X1 U1481 ( .A1(n36288), .A2(\REGISTERS[3][7] ), .B1(n36287), .B2(
        \REGISTERS[31][7] ), .ZN(n36727) );
  AOI22_X1 U1482 ( .A1(n36290), .A2(\REGISTERS[30][7] ), .B1(n36289), .B2(
        \REGISTERS[8][7] ), .ZN(n36726) );
  NAND4_X1 U1483 ( .A1(n36729), .A2(n36728), .A3(n36727), .A4(n36726), .ZN(
        n36735) );
  AOI22_X1 U1484 ( .A1(n36292), .A2(\REGISTERS[11][7] ), .B1(n36291), .B2(
        \REGISTERS[29][7] ), .ZN(n36733) );
  AOI22_X1 U1485 ( .A1(n36294), .A2(\REGISTERS[1][7] ), .B1(n36293), .B2(
        \REGISTERS[16][7] ), .ZN(n36732) );
  AOI22_X1 U1486 ( .A1(n36296), .A2(\REGISTERS[12][7] ), .B1(n36295), .B2(
        \REGISTERS[24][7] ), .ZN(n36731) );
  AOI22_X1 U1487 ( .A1(n36298), .A2(\REGISTERS[20][7] ), .B1(n36297), .B2(
        \REGISTERS[15][7] ), .ZN(n36730) );
  NAND4_X1 U1488 ( .A1(n36733), .A2(n36732), .A3(n36731), .A4(n36730), .ZN(
        n36734) );
  AOI22_X1 U1489 ( .A1(n36759), .A2(\REGISTERS[5][8] ), .B1(n36268), .B2(
        \REGISTERS[22][8] ), .ZN(n36741) );
  AOI22_X1 U1490 ( .A1(n36761), .A2(\REGISTERS[25][8] ), .B1(n36760), .B2(
        \REGISTERS[21][8] ), .ZN(n36740) );
  AOI22_X1 U1491 ( .A1(n36763), .A2(\REGISTERS[17][8] ), .B1(n36762), .B2(
        \REGISTERS[23][8] ), .ZN(n36739) );
  NAND2_X1 U1492 ( .A1(n36274), .A2(\REGISTERS[19][8] ), .ZN(n36738) );
  NAND4_X1 U1493 ( .A1(n36741), .A2(n36740), .A3(n36739), .A4(n36738), .ZN(
        n36757) );
  AOI22_X1 U1494 ( .A1(n36770), .A2(\REGISTERS[14][8] ), .B1(n36769), .B2(
        \REGISTERS[13][8] ), .ZN(n36745) );
  AOI22_X1 U1495 ( .A1(n36772), .A2(\REGISTERS[27][8] ), .B1(n36277), .B2(
        \REGISTERS[4][8] ), .ZN(n36744) );
  AOI22_X1 U1496 ( .A1(n36774), .A2(\REGISTERS[6][8] ), .B1(n36773), .B2(
        \REGISTERS[28][8] ), .ZN(n36743) );
  AOI22_X1 U1497 ( .A1(n36776), .A2(\REGISTERS[26][8] ), .B1(n36775), .B2(
        \REGISTERS[7][8] ), .ZN(n36742) );
  NAND4_X1 U1498 ( .A1(n36745), .A2(n36744), .A3(n36743), .A4(n36742), .ZN(
        n36756) );
  AOI22_X1 U1499 ( .A1(n36782), .A2(\REGISTERS[10][8] ), .B1(n36781), .B2(
        \REGISTERS[9][8] ), .ZN(n36749) );
  AOI22_X1 U1500 ( .A1(n36286), .A2(\REGISTERS[2][8] ), .B1(n36783), .B2(
        \REGISTERS[18][8] ), .ZN(n36748) );
  AOI22_X1 U1501 ( .A1(n36786), .A2(\REGISTERS[3][8] ), .B1(n36785), .B2(
        \REGISTERS[31][8] ), .ZN(n36747) );
  AOI22_X1 U1502 ( .A1(n36788), .A2(\REGISTERS[30][8] ), .B1(n36787), .B2(
        \REGISTERS[8][8] ), .ZN(n36746) );
  NAND4_X1 U1503 ( .A1(n36749), .A2(n36748), .A3(n36747), .A4(n36746), .ZN(
        n36755) );
  AOI22_X1 U1504 ( .A1(n36794), .A2(\REGISTERS[11][8] ), .B1(n36793), .B2(
        \REGISTERS[29][8] ), .ZN(n36753) );
  AOI22_X1 U1505 ( .A1(n36796), .A2(\REGISTERS[1][8] ), .B1(n36795), .B2(
        \REGISTERS[16][8] ), .ZN(n36752) );
  AOI22_X1 U1506 ( .A1(n36798), .A2(\REGISTERS[12][8] ), .B1(n36797), .B2(
        \REGISTERS[24][8] ), .ZN(n36751) );
  AOI22_X1 U1507 ( .A1(n36800), .A2(\REGISTERS[20][8] ), .B1(n36799), .B2(
        \REGISTERS[15][8] ), .ZN(n36750) );
  NAND4_X1 U1508 ( .A1(n36753), .A2(n36752), .A3(n36751), .A4(n36750), .ZN(
        n36754) );
  AOI22_X1 U1509 ( .A1(n36759), .A2(\REGISTERS[5][9] ), .B1(n36758), .B2(
        \REGISTERS[22][9] ), .ZN(n36768) );
  AOI22_X1 U1510 ( .A1(n36761), .A2(\REGISTERS[25][9] ), .B1(n36760), .B2(
        \REGISTERS[21][9] ), .ZN(n36767) );
  AOI22_X1 U1511 ( .A1(n36763), .A2(\REGISTERS[17][9] ), .B1(n36762), .B2(
        \REGISTERS[23][9] ), .ZN(n36766) );
  NAND2_X1 U1512 ( .A1(n36274), .A2(\REGISTERS[19][9] ), .ZN(n36765) );
  NAND4_X1 U1513 ( .A1(n36768), .A2(n36767), .A3(n36766), .A4(n36765), .ZN(
        n36808) );
  AOI22_X1 U1514 ( .A1(n36770), .A2(\REGISTERS[14][9] ), .B1(n36769), .B2(
        \REGISTERS[13][9] ), .ZN(n36780) );
  AOI22_X1 U1515 ( .A1(n36772), .A2(\REGISTERS[27][9] ), .B1(n36277), .B2(
        \REGISTERS[4][9] ), .ZN(n36779) );
  AOI22_X1 U1516 ( .A1(n36774), .A2(\REGISTERS[6][9] ), .B1(n36773), .B2(
        \REGISTERS[28][9] ), .ZN(n36778) );
  AOI22_X1 U1517 ( .A1(n36776), .A2(\REGISTERS[26][9] ), .B1(n36775), .B2(
        \REGISTERS[7][9] ), .ZN(n36777) );
  NAND4_X1 U1518 ( .A1(n36780), .A2(n36779), .A3(n36778), .A4(n36777), .ZN(
        n36807) );
  AOI22_X1 U1519 ( .A1(n36782), .A2(\REGISTERS[10][9] ), .B1(n36781), .B2(
        \REGISTERS[9][9] ), .ZN(n36792) );
  AOI22_X1 U1520 ( .A1(n36286), .A2(\REGISTERS[2][9] ), .B1(n36285), .B2(
        \REGISTERS[18][9] ), .ZN(n36791) );
  AOI22_X1 U1521 ( .A1(n36786), .A2(\REGISTERS[3][9] ), .B1(n36287), .B2(
        \REGISTERS[31][9] ), .ZN(n36790) );
  AOI22_X1 U1522 ( .A1(n36788), .A2(\REGISTERS[30][9] ), .B1(n36787), .B2(
        \REGISTERS[8][9] ), .ZN(n36789) );
  NAND4_X1 U1523 ( .A1(n36792), .A2(n36791), .A3(n36790), .A4(n36789), .ZN(
        n36806) );
  AOI22_X1 U1524 ( .A1(n36794), .A2(\REGISTERS[11][9] ), .B1(n36793), .B2(
        \REGISTERS[29][9] ), .ZN(n36804) );
  AOI22_X1 U1525 ( .A1(n36796), .A2(\REGISTERS[1][9] ), .B1(n36795), .B2(
        \REGISTERS[16][9] ), .ZN(n36803) );
  AOI22_X1 U1526 ( .A1(n36798), .A2(\REGISTERS[12][9] ), .B1(n36797), .B2(
        \REGISTERS[24][9] ), .ZN(n36802) );
  AOI22_X1 U1527 ( .A1(n36800), .A2(\REGISTERS[20][9] ), .B1(n36799), .B2(
        \REGISTERS[15][9] ), .ZN(n36801) );
  NAND4_X1 U1528 ( .A1(n36804), .A2(n36803), .A3(n36802), .A4(n36801), .ZN(
        n36805) );
  NAND3_X1 U1529 ( .A1(ADD_RDB[0]), .A2(ADD_RDB[4]), .A3(n36810), .ZN(n36816)
         );
  INV_X1 U1530 ( .A(ADD_RDB[1]), .ZN(n36820) );
  NAND3_X1 U1531 ( .A1(ADD_RDB[2]), .A2(RESET), .A3(n36820), .ZN(n36827) );
  NOR2_X1 U1532 ( .A1(n36816), .A2(n36827), .ZN(n36829) );
  INV_X1 U1533 ( .A(ADD_RDB[2]), .ZN(n36814) );
  NAND3_X1 U1534 ( .A1(RESET), .A2(ADD_RDB[1]), .A3(n36814), .ZN(n36821) );
  INV_X1 U1535 ( .A(ADD_RDB[0]), .ZN(n36809) );
  NAND3_X1 U1536 ( .A1(ADD_RDB[3]), .A2(ADD_RDB[4]), .A3(n36809), .ZN(n36813)
         );
  NOR2_X1 U1537 ( .A1(n36821), .A2(n36813), .ZN(n36828) );
  INV_X1 U1538 ( .A(ADD_RDB[4]), .ZN(n36817) );
  NAND3_X1 U1539 ( .A1(ADD_RDB[0]), .A2(n36810), .A3(n36817), .ZN(n36815) );
  NAND3_X1 U1540 ( .A1(RESET), .A2(ADD_RDB[2]), .A3(ADD_RDB[1]), .ZN(n36823)
         );
  NOR2_X1 U1541 ( .A1(n36815), .A2(n36823), .ZN(n36831) );
  NAND3_X1 U1542 ( .A1(RESET), .A2(n36814), .A3(n36820), .ZN(n36825) );
  NOR2_X1 U1543 ( .A1(n36815), .A2(n36825), .ZN(n36830) );
  NOR2_X1 U1544 ( .A1(n36827), .A2(n36815), .ZN(n36833) );
  NAND3_X1 U1545 ( .A1(ADD_RDB[4]), .A2(n36810), .A3(n36809), .ZN(n36818) );
  NOR2_X1 U1546 ( .A1(n36818), .A2(n36827), .ZN(n36832) );
  NOR2_X1 U1547 ( .A1(n36821), .A2(n36818), .ZN(n36834) );
  NOR2_X1 U1548 ( .A1(n36821), .A2(n36816), .ZN(n36836) );
  NOR2_X1 U1549 ( .A1(n36813), .A2(n36827), .ZN(n36835) );
  NOR2_X1 U1550 ( .A1(n36816), .A2(n36823), .ZN(n36838) );
  NAND2_X1 U1551 ( .A1(ADD_RDB[2]), .A2(ADD_RDB[1]), .ZN(n36811) );
  NOR2_X1 U1552 ( .A1(ADD_RDB[0]), .A2(ADD_RDB[4]), .ZN(n36812) );
  NAND3_X1 U1553 ( .A1(RESET), .A2(n36812), .A3(n36810), .ZN(n36819) );
  NOR2_X1 U1554 ( .A1(n36811), .A2(n36819), .ZN(n36837) );
  NAND2_X1 U1555 ( .A1(ADD_RDB[3]), .A2(n36812), .ZN(n36824) );
  NOR2_X1 U1556 ( .A1(n36821), .A2(n36824), .ZN(n36840) );
  NOR2_X1 U1557 ( .A1(n36813), .A2(n36825), .ZN(n36839) );
  NAND3_X1 U1558 ( .A1(ADD_RDB[3]), .A2(ADD_RDB[0]), .A3(ADD_RDB[4]), .ZN(
        n36826) );
  NOR2_X1 U1559 ( .A1(n36821), .A2(n36826), .ZN(n36842) );
  NOR2_X1 U1560 ( .A1(n36827), .A2(n36824), .ZN(n36841) );
  NOR2_X1 U1561 ( .A1(n36823), .A2(n36824), .ZN(n36844) );
  NOR2_X1 U1562 ( .A1(n36813), .A2(n36823), .ZN(n36843) );
  NOR3_X1 U1563 ( .A1(ADD_RDB[1]), .A2(n36814), .A3(n36819), .ZN(n36846) );
  NOR2_X1 U1564 ( .A1(n36821), .A2(n36815), .ZN(n36845) );
  NOR2_X1 U1565 ( .A1(n36818), .A2(n36823), .ZN(n36848) );
  NOR2_X1 U1566 ( .A1(n36816), .A2(n36825), .ZN(n36847) );
  NAND3_X1 U1567 ( .A1(ADD_RDB[0]), .A2(ADD_RDB[3]), .A3(n36817), .ZN(n36822)
         );
  NOR2_X1 U1568 ( .A1(n36825), .A2(n36822), .ZN(n36850) );
  NOR2_X1 U1569 ( .A1(n36823), .A2(n36822), .ZN(n36849) );
  NOR2_X1 U1570 ( .A1(n36825), .A2(n36826), .ZN(n36852) );
  NOR2_X1 U1571 ( .A1(n36818), .A2(n36825), .ZN(n36851) );
  NOR3_X1 U1572 ( .A1(ADD_RDB[2]), .A2(n36820), .A3(n36819), .ZN(n36854) );
  NOR2_X1 U1573 ( .A1(n36821), .A2(n36822), .ZN(n36853) );
  NOR2_X1 U1574 ( .A1(n36827), .A2(n36822), .ZN(n36856) );
  NOR2_X1 U1575 ( .A1(n36825), .A2(n36824), .ZN(n36858) );
  NOR2_X1 U1576 ( .A1(n36827), .A2(n36826), .ZN(n36857) );
endmodule


module branch_predictor ( RST, PC_IN, PC_FAIL, IR_IN, IR_FAIL, WRONG_PRE, 
        RIGHT_PRE, NPC_OUT, LINK_ADD, SEL, TAKEN );
  input [31:0] PC_IN;
  input [31:0] PC_FAIL;
  input [31:0] IR_IN;
  input [15:0] IR_FAIL;
  output [31:0] NPC_OUT;
  output [31:0] LINK_ADD;
  input RST, WRONG_PRE, RIGHT_PRE;
  output SEL, TAKEN;
  wire   \CACHE_mem[0][1] , \CACHE_mem[0][0] , \CACHE_mem[1][1] ,
         \CACHE_mem[1][0] , \CACHE_mem[2][1] , \CACHE_mem[2][0] ,
         \CACHE_mem[3][1] , \CACHE_mem[3][0] , \CACHE_mem[4][1] ,
         \CACHE_mem[4][0] , \CACHE_mem[5][1] , \CACHE_mem[5][0] ,
         \CACHE_mem[6][1] , \CACHE_mem[6][0] , \CACHE_mem[7][1] ,
         \CACHE_mem[7][0] , \CACHE_mem[8][1] , \CACHE_mem[8][0] ,
         \CACHE_mem[9][1] , \CACHE_mem[9][0] , \CACHE_mem[10][1] ,
         \CACHE_mem[10][0] , \CACHE_mem[11][1] , \CACHE_mem[11][0] ,
         \CACHE_mem[12][1] , \CACHE_mem[12][0] , \CACHE_mem[13][1] ,
         \CACHE_mem[13][0] , \CACHE_mem[14][1] , \CACHE_mem[14][0] ,
         \CACHE_mem[15][1] , \CACHE_mem[15][0] , \CACHE_mem[16][1] ,
         \CACHE_mem[16][0] , \CACHE_mem[17][1] , \CACHE_mem[17][0] ,
         \CACHE_mem[18][1] , \CACHE_mem[18][0] , \CACHE_mem[19][1] ,
         \CACHE_mem[19][0] , \CACHE_mem[20][1] , \CACHE_mem[20][0] ,
         \CACHE_mem[21][1] , \CACHE_mem[21][0] , \CACHE_mem[22][1] ,
         \CACHE_mem[22][0] , \CACHE_mem[23][1] , \CACHE_mem[23][0] ,
         \CACHE_mem[24][1] , \CACHE_mem[24][0] , \CACHE_mem[25][1] ,
         \CACHE_mem[25][0] , \CACHE_mem[26][1] , \CACHE_mem[26][0] ,
         \CACHE_mem[27][1] , \CACHE_mem[27][0] , \CACHE_mem[28][1] ,
         \CACHE_mem[28][0] , \CACHE_mem[29][1] , \CACHE_mem[29][0] ,
         \CACHE_mem[30][1] , \CACHE_mem[30][0] , \CACHE_mem[31][1] ,
         \CACHE_mem[31][0] , N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N323, N356, N357, N358, N362, N387, N388, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n60,
         \add_65/carry[31] , \add_65/carry[30] , \add_65/carry[29] ,
         \add_65/carry[28] , \add_65/carry[27] , \add_65/carry[26] ,
         \add_65/carry[25] , \add_65/carry[24] , \add_65/carry[23] ,
         \add_65/carry[22] , \add_65/carry[21] , \add_65/carry[20] ,
         \add_65/carry[19] , \add_65/carry[18] , \add_65/carry[17] ,
         \add_65/carry[16] , \add_65/carry[15] , \add_65/carry[14] ,
         \add_65/carry[13] , \add_65/carry[12] , \add_65/carry[11] ,
         \add_65/carry[10] , \add_65/carry[9] , \add_65/carry[8] ,
         \add_65/carry[7] , \add_65/carry[6] , \add_65/carry[5] ,
         \add_65/carry[4] , \add_65/carry[3] , \add_65/carry[2] , \add_59/n1 ,
         \add_59/carry[31] , \add_59/carry[30] , \add_59/carry[29] ,
         \add_59/carry[28] , \add_59/carry[27] , \add_59/carry[26] ,
         \add_59/carry[25] , \add_59/carry[24] , \add_59/carry[23] ,
         \add_59/carry[22] , \add_59/carry[21] , \add_59/carry[20] ,
         \add_59/carry[19] , \add_59/carry[18] , \add_59/carry[17] ,
         \add_59/carry[16] , \add_59/carry[15] , \add_59/carry[14] ,
         \add_59/carry[13] , \add_59/carry[12] , \add_59/carry[11] ,
         \add_59/carry[10] , \add_59/carry[9] , \add_59/carry[8] ,
         \add_59/carry[7] , \add_59/carry[6] , \add_59/carry[5] ,
         \add_59/carry[4] , \add_59/carry[3] , \add_59/carry[2] ,
         \add_53_aco/n2 , \add_53_aco/carry[31] , \add_53_aco/carry[30] ,
         \add_53_aco/carry[29] , \add_53_aco/carry[28] ,
         \add_53_aco/carry[27] , \add_53_aco/carry[26] ,
         \add_53_aco/carry[25] , \add_53_aco/carry[24] ,
         \add_53_aco/carry[23] , \add_53_aco/carry[22] ,
         \add_53_aco/carry[21] , \add_53_aco/carry[20] ,
         \add_53_aco/carry[19] , \add_53_aco/carry[18] ,
         \add_53_aco/carry[17] , \add_53_aco/carry[16] ,
         \add_53_aco/carry[15] , \add_53_aco/carry[14] ,
         \add_53_aco/carry[13] , \add_53_aco/carry[12] ,
         \add_53_aco/carry[11] , \add_53_aco/carry[10] , \add_53_aco/carry[9] ,
         \add_53_aco/carry[8] , \add_53_aco/carry[7] , \add_53_aco/carry[6] ,
         \add_53_aco/carry[5] , \add_53_aco/carry[4] , \add_53_aco/carry[3] ,
         \add_53_aco/carry[2] , n62, n286, n291, n59, n1, n2, n3, n4, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n61, n281, n282, n283, n284,
         n285, n287, n288, n289, n290, n292, n293, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318;
  assign N113 = PC_IN[0];
  assign N114 = PC_IN[1];

  DLH_X1 \NPC_OUT_reg[31]  ( .G(N323), .D(n1), .Q(NPC_OUT[31]) );
  DLH_X1 \NPC_OUT_reg[30]  ( .G(N323), .D(n2), .Q(NPC_OUT[30]) );
  DLH_X1 \NPC_OUT_reg[29]  ( .G(N323), .D(n3), .Q(NPC_OUT[29]) );
  DLH_X1 \NPC_OUT_reg[28]  ( .G(N323), .D(n4), .Q(NPC_OUT[28]) );
  DLH_X1 \NPC_OUT_reg[27]  ( .G(N323), .D(n20), .Q(NPC_OUT[27]) );
  DLH_X1 \NPC_OUT_reg[26]  ( .G(N323), .D(n21), .Q(NPC_OUT[26]) );
  DLH_X1 \NPC_OUT_reg[25]  ( .G(N323), .D(n22), .Q(NPC_OUT[25]) );
  DLH_X1 \NPC_OUT_reg[24]  ( .G(N323), .D(n23), .Q(NPC_OUT[24]) );
  DLH_X1 \NPC_OUT_reg[23]  ( .G(N323), .D(n24), .Q(NPC_OUT[23]) );
  DLH_X1 \NPC_OUT_reg[22]  ( .G(N323), .D(n25), .Q(NPC_OUT[22]) );
  DLH_X1 \NPC_OUT_reg[21]  ( .G(N323), .D(n26), .Q(NPC_OUT[21]) );
  DLH_X1 \NPC_OUT_reg[20]  ( .G(N323), .D(n27), .Q(NPC_OUT[20]) );
  DLH_X1 \NPC_OUT_reg[19]  ( .G(N323), .D(n28), .Q(NPC_OUT[19]) );
  DLH_X1 \NPC_OUT_reg[18]  ( .G(N323), .D(n29), .Q(NPC_OUT[18]) );
  DLH_X1 \NPC_OUT_reg[17]  ( .G(N323), .D(n30), .Q(NPC_OUT[17]) );
  DLH_X1 \NPC_OUT_reg[16]  ( .G(N323), .D(n31), .Q(NPC_OUT[16]) );
  DLH_X1 \NPC_OUT_reg[15]  ( .G(N323), .D(n32), .Q(NPC_OUT[15]) );
  DLH_X1 \NPC_OUT_reg[14]  ( .G(N323), .D(n33), .Q(NPC_OUT[14]) );
  DLH_X1 \NPC_OUT_reg[13]  ( .G(N323), .D(n34), .Q(NPC_OUT[13]) );
  DLH_X1 \NPC_OUT_reg[12]  ( .G(N323), .D(n35), .Q(NPC_OUT[12]) );
  DLH_X1 \NPC_OUT_reg[11]  ( .G(N323), .D(n36), .Q(NPC_OUT[11]) );
  DLH_X1 \NPC_OUT_reg[10]  ( .G(N323), .D(n37), .Q(NPC_OUT[10]) );
  DLH_X1 \NPC_OUT_reg[9]  ( .G(N323), .D(n38), .Q(NPC_OUT[9]) );
  DLH_X1 \NPC_OUT_reg[8]  ( .G(N323), .D(n39), .Q(NPC_OUT[8]) );
  DLH_X1 \NPC_OUT_reg[7]  ( .G(N323), .D(n40), .Q(NPC_OUT[7]) );
  DLH_X1 \NPC_OUT_reg[6]  ( .G(N323), .D(n41), .Q(NPC_OUT[6]) );
  DLH_X1 \NPC_OUT_reg[5]  ( .G(N323), .D(n42), .Q(NPC_OUT[5]) );
  DLH_X1 \NPC_OUT_reg[4]  ( .G(N323), .D(n43), .Q(NPC_OUT[4]) );
  DLH_X1 \NPC_OUT_reg[3]  ( .G(N323), .D(n44), .Q(NPC_OUT[3]) );
  DLH_X1 \NPC_OUT_reg[2]  ( .G(N323), .D(n45), .Q(NPC_OUT[2]) );
  DLH_X1 \NPC_OUT_reg[1]  ( .G(N323), .D(n46), .Q(NPC_OUT[1]) );
  DLH_X1 \NPC_OUT_reg[0]  ( .G(N323), .D(n60), .Q(NPC_OUT[0]) );
  DLH_X1 \LINK_ADD_reg[31]  ( .G(N356), .D(N388), .Q(LINK_ADD[31]) );
  DLH_X1 \LINK_ADD_reg[30]  ( .G(N356), .D(N387), .Q(LINK_ADD[30]) );
  DLH_X1 \LINK_ADD_reg[29]  ( .G(n5092), .D(n48), .Q(LINK_ADD[29]) );
  DLH_X1 \LINK_ADD_reg[28]  ( .G(n5092), .D(n287), .Q(LINK_ADD[28]) );
  DLH_X1 \LINK_ADD_reg[27]  ( .G(n5092), .D(n49), .Q(LINK_ADD[27]) );
  DLH_X1 \LINK_ADD_reg[26]  ( .G(n5092), .D(n283), .Q(LINK_ADD[26]) );
  DLH_X1 \LINK_ADD_reg[25]  ( .G(n5092), .D(n50), .Q(LINK_ADD[25]) );
  DLH_X1 \LINK_ADD_reg[24]  ( .G(n5092), .D(n293), .Q(LINK_ADD[24]) );
  DLH_X1 \LINK_ADD_reg[23]  ( .G(n5092), .D(n51), .Q(LINK_ADD[23]) );
  DLH_X1 \LINK_ADD_reg[22]  ( .G(n5092), .D(n290), .Q(LINK_ADD[22]) );
  DLH_X1 \LINK_ADD_reg[21]  ( .G(n5092), .D(n52), .Q(LINK_ADD[21]) );
  DLH_X1 \LINK_ADD_reg[20]  ( .G(n5092), .D(n289), .Q(LINK_ADD[20]) );
  DLH_X1 \LINK_ADD_reg[19]  ( .G(n5092), .D(n53), .Q(LINK_ADD[19]) );
  DLH_X1 \LINK_ADD_reg[18]  ( .G(n5092), .D(n288), .Q(LINK_ADD[18]) );
  DLH_X1 \LINK_ADD_reg[17]  ( .G(n5092), .D(n54), .Q(LINK_ADD[17]) );
  DLH_X1 \LINK_ADD_reg[16]  ( .G(n5092), .D(n285), .Q(LINK_ADD[16]) );
  DLH_X1 \LINK_ADD_reg[15]  ( .G(n5092), .D(n55), .Q(LINK_ADD[15]) );
  DLH_X1 \LINK_ADD_reg[14]  ( .G(n5092), .D(n284), .Q(LINK_ADD[14]) );
  DLH_X1 \LINK_ADD_reg[13]  ( .G(n5092), .D(n56), .Q(LINK_ADD[13]) );
  DLH_X1 \LINK_ADD_reg[12]  ( .G(n5092), .D(n292), .Q(LINK_ADD[12]) );
  DLH_X1 \LINK_ADD_reg[11]  ( .G(n5092), .D(n57), .Q(LINK_ADD[11]) );
  DLH_X1 \LINK_ADD_reg[10]  ( .G(n5092), .D(n281), .Q(LINK_ADD[10]) );
  DLH_X1 \LINK_ADD_reg[9]  ( .G(n5092), .D(n58), .Q(LINK_ADD[9]) );
  DLH_X1 \LINK_ADD_reg[8]  ( .G(n5092), .D(n282), .Q(LINK_ADD[8]) );
  DLH_X1 \LINK_ADD_reg[7]  ( .G(N356), .D(n61), .Q(LINK_ADD[7]) );
  DLH_X1 \LINK_ADD_reg[6]  ( .G(N356), .D(n291), .Q(LINK_ADD[6]) );
  DLH_X1 \LINK_ADD_reg[5]  ( .G(N356), .D(N362), .Q(LINK_ADD[5]) );
  DLH_X1 \LINK_ADD_reg[4]  ( .G(N356), .D(n286), .Q(LINK_ADD[4]) );
  DLH_X1 \LINK_ADD_reg[3]  ( .G(N356), .D(n59), .Q(LINK_ADD[3]) );
  DLH_X1 \LINK_ADD_reg[2]  ( .G(N356), .D(n62), .Q(LINK_ADD[2]) );
  DLH_X1 \LINK_ADD_reg[1]  ( .G(N356), .D(N358), .Q(LINK_ADD[1]) );
  DLH_X1 \LINK_ADD_reg[0]  ( .G(N356), .D(N357), .Q(LINK_ADD[0]) );
  DLH_X1 \CACHE_mem_reg[0][1]  ( .G(N643), .D(N645), .Q(\CACHE_mem[0][1] ) );
  DLH_X1 \CACHE_mem_reg[0][0]  ( .G(N643), .D(N644), .Q(\CACHE_mem[0][0] ) );
  DLH_X1 \CACHE_mem_reg[1][1]  ( .G(N642), .D(N645), .Q(\CACHE_mem[1][1] ) );
  DLH_X1 \CACHE_mem_reg[1][0]  ( .G(N642), .D(N644), .Q(\CACHE_mem[1][0] ) );
  DLH_X1 \CACHE_mem_reg[2][1]  ( .G(N641), .D(N645), .Q(\CACHE_mem[2][1] ) );
  DLH_X1 \CACHE_mem_reg[2][0]  ( .G(N641), .D(N644), .Q(\CACHE_mem[2][0] ) );
  DLH_X1 \CACHE_mem_reg[3][1]  ( .G(N640), .D(N645), .Q(\CACHE_mem[3][1] ) );
  DLH_X1 \CACHE_mem_reg[3][0]  ( .G(N640), .D(N644), .Q(\CACHE_mem[3][0] ) );
  DLH_X1 \CACHE_mem_reg[4][1]  ( .G(N639), .D(N645), .Q(\CACHE_mem[4][1] ) );
  DLH_X1 \CACHE_mem_reg[4][0]  ( .G(N639), .D(N644), .Q(\CACHE_mem[4][0] ) );
  DLH_X1 \CACHE_mem_reg[5][1]  ( .G(N638), .D(N645), .Q(\CACHE_mem[5][1] ) );
  DLH_X1 \CACHE_mem_reg[5][0]  ( .G(N638), .D(N644), .Q(\CACHE_mem[5][0] ) );
  DLH_X1 \CACHE_mem_reg[6][1]  ( .G(N637), .D(N645), .Q(\CACHE_mem[6][1] ) );
  DLH_X1 \CACHE_mem_reg[6][0]  ( .G(N637), .D(N644), .Q(\CACHE_mem[6][0] ) );
  DLH_X1 \CACHE_mem_reg[7][1]  ( .G(N636), .D(N645), .Q(\CACHE_mem[7][1] ) );
  DLH_X1 \CACHE_mem_reg[7][0]  ( .G(N636), .D(N644), .Q(\CACHE_mem[7][0] ) );
  DLH_X1 \CACHE_mem_reg[8][1]  ( .G(N635), .D(N645), .Q(\CACHE_mem[8][1] ) );
  DLH_X1 \CACHE_mem_reg[8][0]  ( .G(N635), .D(N644), .Q(\CACHE_mem[8][0] ) );
  DLH_X1 \CACHE_mem_reg[9][1]  ( .G(N634), .D(N645), .Q(\CACHE_mem[9][1] ) );
  DLH_X1 \CACHE_mem_reg[9][0]  ( .G(N634), .D(N644), .Q(\CACHE_mem[9][0] ) );
  DLH_X1 \CACHE_mem_reg[10][1]  ( .G(N633), .D(N645), .Q(\CACHE_mem[10][1] )
         );
  DLH_X1 \CACHE_mem_reg[10][0]  ( .G(N633), .D(N644), .Q(\CACHE_mem[10][0] )
         );
  DLH_X1 \CACHE_mem_reg[11][1]  ( .G(N632), .D(N645), .Q(\CACHE_mem[11][1] )
         );
  DLH_X1 \CACHE_mem_reg[11][0]  ( .G(N632), .D(N644), .Q(\CACHE_mem[11][0] )
         );
  DLH_X1 \CACHE_mem_reg[12][1]  ( .G(N631), .D(N645), .Q(\CACHE_mem[12][1] )
         );
  DLH_X1 \CACHE_mem_reg[12][0]  ( .G(N631), .D(N644), .Q(\CACHE_mem[12][0] )
         );
  DLH_X1 \CACHE_mem_reg[13][1]  ( .G(N630), .D(N645), .Q(\CACHE_mem[13][1] )
         );
  DLH_X1 \CACHE_mem_reg[13][0]  ( .G(N630), .D(N644), .Q(\CACHE_mem[13][0] )
         );
  DLH_X1 \CACHE_mem_reg[14][1]  ( .G(N629), .D(N645), .Q(\CACHE_mem[14][1] )
         );
  DLH_X1 \CACHE_mem_reg[14][0]  ( .G(N629), .D(N644), .Q(\CACHE_mem[14][0] )
         );
  DLH_X1 \CACHE_mem_reg[15][1]  ( .G(N628), .D(N645), .Q(\CACHE_mem[15][1] )
         );
  DLH_X1 \CACHE_mem_reg[15][0]  ( .G(N628), .D(N644), .Q(\CACHE_mem[15][0] )
         );
  DLH_X1 \CACHE_mem_reg[16][1]  ( .G(N627), .D(N645), .Q(\CACHE_mem[16][1] )
         );
  DLH_X1 \CACHE_mem_reg[16][0]  ( .G(N627), .D(N644), .Q(\CACHE_mem[16][0] )
         );
  DLH_X1 \CACHE_mem_reg[17][1]  ( .G(N626), .D(N645), .Q(\CACHE_mem[17][1] )
         );
  DLH_X1 \CACHE_mem_reg[17][0]  ( .G(N626), .D(N644), .Q(\CACHE_mem[17][0] )
         );
  DLH_X1 \CACHE_mem_reg[18][1]  ( .G(N625), .D(N645), .Q(\CACHE_mem[18][1] )
         );
  DLH_X1 \CACHE_mem_reg[18][0]  ( .G(N625), .D(N644), .Q(\CACHE_mem[18][0] )
         );
  DLH_X1 \CACHE_mem_reg[19][1]  ( .G(N624), .D(N645), .Q(\CACHE_mem[19][1] )
         );
  DLH_X1 \CACHE_mem_reg[19][0]  ( .G(N624), .D(N644), .Q(\CACHE_mem[19][0] )
         );
  DLH_X1 \CACHE_mem_reg[20][1]  ( .G(N623), .D(N645), .Q(\CACHE_mem[20][1] )
         );
  DLH_X1 \CACHE_mem_reg[20][0]  ( .G(N623), .D(N644), .Q(\CACHE_mem[20][0] )
         );
  DLH_X1 \CACHE_mem_reg[21][1]  ( .G(N622), .D(N645), .Q(\CACHE_mem[21][1] )
         );
  DLH_X1 \CACHE_mem_reg[21][0]  ( .G(N622), .D(N644), .Q(\CACHE_mem[21][0] )
         );
  DLH_X1 \CACHE_mem_reg[22][1]  ( .G(N621), .D(N645), .Q(\CACHE_mem[22][1] )
         );
  DLH_X1 \CACHE_mem_reg[22][0]  ( .G(N621), .D(N644), .Q(\CACHE_mem[22][0] )
         );
  DLH_X1 \CACHE_mem_reg[23][1]  ( .G(N620), .D(N645), .Q(\CACHE_mem[23][1] )
         );
  DLH_X1 \CACHE_mem_reg[23][0]  ( .G(N620), .D(N644), .Q(\CACHE_mem[23][0] )
         );
  DLH_X1 \CACHE_mem_reg[24][1]  ( .G(N619), .D(N645), .Q(\CACHE_mem[24][1] )
         );
  DLH_X1 \CACHE_mem_reg[24][0]  ( .G(N619), .D(N644), .Q(\CACHE_mem[24][0] )
         );
  DLH_X1 \CACHE_mem_reg[25][1]  ( .G(N618), .D(N645), .Q(\CACHE_mem[25][1] )
         );
  DLH_X1 \CACHE_mem_reg[25][0]  ( .G(N618), .D(N644), .Q(\CACHE_mem[25][0] )
         );
  DLH_X1 \CACHE_mem_reg[26][1]  ( .G(N617), .D(N645), .Q(\CACHE_mem[26][1] )
         );
  DLH_X1 \CACHE_mem_reg[26][0]  ( .G(N617), .D(N644), .Q(\CACHE_mem[26][0] )
         );
  DLH_X1 \CACHE_mem_reg[27][1]  ( .G(N616), .D(N645), .Q(\CACHE_mem[27][1] )
         );
  DLH_X1 \CACHE_mem_reg[27][0]  ( .G(N616), .D(N644), .Q(\CACHE_mem[27][0] )
         );
  DLH_X1 \CACHE_mem_reg[28][1]  ( .G(N615), .D(N645), .Q(\CACHE_mem[28][1] )
         );
  DLH_X1 \CACHE_mem_reg[28][0]  ( .G(N615), .D(N644), .Q(\CACHE_mem[28][0] )
         );
  DLH_X1 \CACHE_mem_reg[29][1]  ( .G(N614), .D(N645), .Q(\CACHE_mem[29][1] )
         );
  DLH_X1 \CACHE_mem_reg[29][0]  ( .G(N614), .D(N644), .Q(\CACHE_mem[29][0] )
         );
  DLH_X1 \CACHE_mem_reg[30][1]  ( .G(N613), .D(N645), .Q(\CACHE_mem[30][1] )
         );
  DLH_X1 \CACHE_mem_reg[30][0]  ( .G(N613), .D(N644), .Q(\CACHE_mem[30][0] )
         );
  DLH_X1 \CACHE_mem_reg[31][1]  ( .G(N612), .D(N645), .Q(\CACHE_mem[31][1] )
         );
  DLH_X1 \CACHE_mem_reg[31][0]  ( .G(N612), .D(N644), .Q(\CACHE_mem[31][0] )
         );
  FA_X1 \add_65/U1_1  ( .A(N114), .B(IR_IN[1]), .CI(\add_59/n1 ), .CO(
        \add_65/carry[2] ), .S(N220) );
  FA_X1 \add_65/U1_2  ( .A(PC_IN[2]), .B(IR_IN[2]), .CI(\add_65/carry[2] ), 
        .CO(\add_65/carry[3] ), .S(N221) );
  FA_X1 \add_65/U1_3  ( .A(PC_IN[3]), .B(IR_IN[3]), .CI(\add_65/carry[3] ), 
        .CO(\add_65/carry[4] ), .S(N222) );
  FA_X1 \add_65/U1_4  ( .A(PC_IN[4]), .B(IR_IN[4]), .CI(\add_65/carry[4] ), 
        .CO(\add_65/carry[5] ), .S(N223) );
  FA_X1 \add_65/U1_5  ( .A(PC_IN[5]), .B(IR_IN[5]), .CI(\add_65/carry[5] ), 
        .CO(\add_65/carry[6] ), .S(N224) );
  FA_X1 \add_65/U1_6  ( .A(PC_IN[6]), .B(IR_IN[6]), .CI(\add_65/carry[6] ), 
        .CO(\add_65/carry[7] ), .S(N225) );
  FA_X1 \add_65/U1_7  ( .A(PC_IN[7]), .B(IR_IN[7]), .CI(\add_65/carry[7] ), 
        .CO(\add_65/carry[8] ), .S(N226) );
  FA_X1 \add_65/U1_8  ( .A(PC_IN[8]), .B(IR_IN[8]), .CI(\add_65/carry[8] ), 
        .CO(\add_65/carry[9] ), .S(N227) );
  FA_X1 \add_65/U1_9  ( .A(PC_IN[9]), .B(IR_IN[9]), .CI(\add_65/carry[9] ), 
        .CO(\add_65/carry[10] ), .S(N228) );
  FA_X1 \add_65/U1_10  ( .A(PC_IN[10]), .B(IR_IN[10]), .CI(\add_65/carry[10] ), 
        .CO(\add_65/carry[11] ), .S(N229) );
  FA_X1 \add_65/U1_11  ( .A(PC_IN[11]), .B(IR_IN[11]), .CI(\add_65/carry[11] ), 
        .CO(\add_65/carry[12] ), .S(N230) );
  FA_X1 \add_65/U1_12  ( .A(PC_IN[12]), .B(IR_IN[12]), .CI(\add_65/carry[12] ), 
        .CO(\add_65/carry[13] ), .S(N231) );
  FA_X1 \add_65/U1_13  ( .A(PC_IN[13]), .B(IR_IN[13]), .CI(\add_65/carry[13] ), 
        .CO(\add_65/carry[14] ), .S(N232) );
  FA_X1 \add_65/U1_14  ( .A(PC_IN[14]), .B(IR_IN[14]), .CI(\add_65/carry[14] ), 
        .CO(\add_65/carry[15] ), .S(N233) );
  FA_X1 \add_65/U1_15  ( .A(PC_IN[15]), .B(IR_IN[15]), .CI(\add_65/carry[15] ), 
        .CO(\add_65/carry[16] ), .S(N234) );
  FA_X1 \add_65/U1_16  ( .A(PC_IN[16]), .B(IR_IN[15]), .CI(\add_65/carry[16] ), 
        .CO(\add_65/carry[17] ), .S(N235) );
  FA_X1 \add_65/U1_17  ( .A(PC_IN[17]), .B(IR_IN[15]), .CI(\add_65/carry[17] ), 
        .CO(\add_65/carry[18] ), .S(N236) );
  FA_X1 \add_65/U1_18  ( .A(PC_IN[18]), .B(IR_IN[15]), .CI(\add_65/carry[18] ), 
        .CO(\add_65/carry[19] ), .S(N237) );
  FA_X1 \add_65/U1_19  ( .A(PC_IN[19]), .B(IR_IN[15]), .CI(\add_65/carry[19] ), 
        .CO(\add_65/carry[20] ), .S(N238) );
  FA_X1 \add_65/U1_20  ( .A(PC_IN[20]), .B(IR_IN[15]), .CI(\add_65/carry[20] ), 
        .CO(\add_65/carry[21] ), .S(N239) );
  FA_X1 \add_65/U1_21  ( .A(PC_IN[21]), .B(IR_IN[15]), .CI(\add_65/carry[21] ), 
        .CO(\add_65/carry[22] ), .S(N240) );
  FA_X1 \add_65/U1_22  ( .A(PC_IN[22]), .B(IR_IN[15]), .CI(\add_65/carry[22] ), 
        .CO(\add_65/carry[23] ), .S(N241) );
  FA_X1 \add_65/U1_23  ( .A(PC_IN[23]), .B(IR_IN[15]), .CI(\add_65/carry[23] ), 
        .CO(\add_65/carry[24] ), .S(N242) );
  FA_X1 \add_65/U1_24  ( .A(PC_IN[24]), .B(IR_IN[15]), .CI(\add_65/carry[24] ), 
        .CO(\add_65/carry[25] ), .S(N243) );
  FA_X1 \add_65/U1_25  ( .A(PC_IN[25]), .B(IR_IN[15]), .CI(\add_65/carry[25] ), 
        .CO(\add_65/carry[26] ), .S(N244) );
  FA_X1 \add_65/U1_26  ( .A(PC_IN[26]), .B(IR_IN[15]), .CI(\add_65/carry[26] ), 
        .CO(\add_65/carry[27] ), .S(N245) );
  FA_X1 \add_65/U1_27  ( .A(PC_IN[27]), .B(IR_IN[15]), .CI(\add_65/carry[27] ), 
        .CO(\add_65/carry[28] ), .S(N246) );
  FA_X1 \add_65/U1_28  ( .A(PC_IN[28]), .B(IR_IN[15]), .CI(\add_65/carry[28] ), 
        .CO(\add_65/carry[29] ), .S(N247) );
  FA_X1 \add_65/U1_29  ( .A(PC_IN[29]), .B(IR_IN[15]), .CI(\add_65/carry[29] ), 
        .CO(\add_65/carry[30] ), .S(N248) );
  FA_X1 \add_65/U1_30  ( .A(PC_IN[30]), .B(IR_IN[15]), .CI(\add_65/carry[30] ), 
        .CO(\add_65/carry[31] ), .S(N249) );
  FA_X1 \add_65/U1_31  ( .A(PC_IN[31]), .B(IR_IN[15]), .CI(\add_65/carry[31] ), 
        .S(N250) );
  FA_X1 \add_59/U1_1  ( .A(N114), .B(IR_IN[1]), .CI(\add_59/n1 ), .CO(
        \add_59/carry[2] ), .S(N82) );
  FA_X1 \add_59/U1_2  ( .A(PC_IN[2]), .B(IR_IN[2]), .CI(\add_59/carry[2] ), 
        .CO(\add_59/carry[3] ), .S(N83) );
  FA_X1 \add_59/U1_3  ( .A(PC_IN[3]), .B(IR_IN[3]), .CI(\add_59/carry[3] ), 
        .CO(\add_59/carry[4] ), .S(N84) );
  FA_X1 \add_59/U1_4  ( .A(PC_IN[4]), .B(IR_IN[4]), .CI(\add_59/carry[4] ), 
        .CO(\add_59/carry[5] ), .S(N85) );
  FA_X1 \add_59/U1_5  ( .A(PC_IN[5]), .B(IR_IN[5]), .CI(\add_59/carry[5] ), 
        .CO(\add_59/carry[6] ), .S(N86) );
  FA_X1 \add_59/U1_6  ( .A(PC_IN[6]), .B(IR_IN[6]), .CI(\add_59/carry[6] ), 
        .CO(\add_59/carry[7] ), .S(N87) );
  FA_X1 \add_59/U1_7  ( .A(PC_IN[7]), .B(IR_IN[7]), .CI(\add_59/carry[7] ), 
        .CO(\add_59/carry[8] ), .S(N88) );
  FA_X1 \add_59/U1_8  ( .A(PC_IN[8]), .B(IR_IN[8]), .CI(\add_59/carry[8] ), 
        .CO(\add_59/carry[9] ), .S(N89) );
  FA_X1 \add_59/U1_9  ( .A(PC_IN[9]), .B(IR_IN[9]), .CI(\add_59/carry[9] ), 
        .CO(\add_59/carry[10] ), .S(N90) );
  FA_X1 \add_59/U1_10  ( .A(PC_IN[10]), .B(IR_IN[10]), .CI(\add_59/carry[10] ), 
        .CO(\add_59/carry[11] ), .S(N91) );
  FA_X1 \add_59/U1_11  ( .A(PC_IN[11]), .B(IR_IN[11]), .CI(\add_59/carry[11] ), 
        .CO(\add_59/carry[12] ), .S(N92) );
  FA_X1 \add_59/U1_12  ( .A(PC_IN[12]), .B(IR_IN[12]), .CI(\add_59/carry[12] ), 
        .CO(\add_59/carry[13] ), .S(N93) );
  FA_X1 \add_59/U1_13  ( .A(PC_IN[13]), .B(IR_IN[13]), .CI(\add_59/carry[13] ), 
        .CO(\add_59/carry[14] ), .S(N94) );
  FA_X1 \add_59/U1_14  ( .A(PC_IN[14]), .B(IR_IN[14]), .CI(\add_59/carry[14] ), 
        .CO(\add_59/carry[15] ), .S(N95) );
  FA_X1 \add_59/U1_15  ( .A(PC_IN[15]), .B(IR_IN[15]), .CI(\add_59/carry[15] ), 
        .CO(\add_59/carry[16] ), .S(N96) );
  FA_X1 \add_59/U1_16  ( .A(PC_IN[16]), .B(IR_IN[16]), .CI(\add_59/carry[16] ), 
        .CO(\add_59/carry[17] ), .S(N97) );
  FA_X1 \add_59/U1_17  ( .A(PC_IN[17]), .B(IR_IN[17]), .CI(\add_59/carry[17] ), 
        .CO(\add_59/carry[18] ), .S(N98) );
  FA_X1 \add_59/U1_18  ( .A(PC_IN[18]), .B(IR_IN[18]), .CI(\add_59/carry[18] ), 
        .CO(\add_59/carry[19] ), .S(N99) );
  FA_X1 \add_59/U1_19  ( .A(PC_IN[19]), .B(IR_IN[19]), .CI(\add_59/carry[19] ), 
        .CO(\add_59/carry[20] ), .S(N100) );
  FA_X1 \add_59/U1_20  ( .A(PC_IN[20]), .B(IR_IN[20]), .CI(\add_59/carry[20] ), 
        .CO(\add_59/carry[21] ), .S(N101) );
  FA_X1 \add_59/U1_21  ( .A(PC_IN[21]), .B(IR_IN[21]), .CI(\add_59/carry[21] ), 
        .CO(\add_59/carry[22] ), .S(N102) );
  FA_X1 \add_59/U1_22  ( .A(PC_IN[22]), .B(IR_IN[22]), .CI(\add_59/carry[22] ), 
        .CO(\add_59/carry[23] ), .S(N103) );
  FA_X1 \add_59/U1_23  ( .A(PC_IN[23]), .B(IR_IN[23]), .CI(\add_59/carry[23] ), 
        .CO(\add_59/carry[24] ), .S(N104) );
  FA_X1 \add_59/U1_24  ( .A(PC_IN[24]), .B(IR_IN[24]), .CI(\add_59/carry[24] ), 
        .CO(\add_59/carry[25] ), .S(N105) );
  FA_X1 \add_59/U1_25  ( .A(PC_IN[25]), .B(IR_IN[25]), .CI(\add_59/carry[25] ), 
        .CO(\add_59/carry[26] ), .S(N106) );
  FA_X1 \add_59/U1_26  ( .A(PC_IN[26]), .B(IR_IN[25]), .CI(\add_59/carry[26] ), 
        .CO(\add_59/carry[27] ), .S(N107) );
  FA_X1 \add_59/U1_27  ( .A(PC_IN[27]), .B(IR_IN[25]), .CI(\add_59/carry[27] ), 
        .CO(\add_59/carry[28] ), .S(N108) );
  FA_X1 \add_59/U1_28  ( .A(PC_IN[28]), .B(IR_IN[25]), .CI(\add_59/carry[28] ), 
        .CO(\add_59/carry[29] ), .S(N109) );
  FA_X1 \add_59/U1_29  ( .A(PC_IN[29]), .B(IR_IN[25]), .CI(\add_59/carry[29] ), 
        .CO(\add_59/carry[30] ), .S(N110) );
  FA_X1 \add_59/U1_30  ( .A(PC_IN[30]), .B(IR_IN[25]), .CI(\add_59/carry[30] ), 
        .CO(\add_59/carry[31] ), .S(N111) );
  FA_X1 \add_59/U1_31  ( .A(PC_IN[31]), .B(IR_IN[25]), .CI(\add_59/carry[31] ), 
        .S(N112) );
  FA_X1 \add_53_aco/U1_1  ( .A(PC_FAIL[1]), .B(n6), .CI(\add_53_aco/n2 ), .CO(
        \add_53_aco/carry[2] ), .S(N47) );
  FA_X1 \add_53_aco/U1_2  ( .A(PC_FAIL[2]), .B(n8), .CI(\add_53_aco/carry[2] ), 
        .CO(\add_53_aco/carry[3] ), .S(N48) );
  FA_X1 \add_53_aco/U1_3  ( .A(PC_FAIL[3]), .B(n9), .CI(\add_53_aco/carry[3] ), 
        .CO(\add_53_aco/carry[4] ), .S(N49) );
  FA_X1 \add_53_aco/U1_4  ( .A(PC_FAIL[4]), .B(n10), .CI(\add_53_aco/carry[4] ), .CO(\add_53_aco/carry[5] ), .S(N50) );
  FA_X1 \add_53_aco/U1_5  ( .A(PC_FAIL[5]), .B(n7), .CI(\add_53_aco/carry[5] ), 
        .CO(\add_53_aco/carry[6] ), .S(N51) );
  FA_X1 \add_53_aco/U1_6  ( .A(PC_FAIL[6]), .B(n11), .CI(\add_53_aco/carry[6] ), .CO(\add_53_aco/carry[7] ), .S(N52) );
  FA_X1 \add_53_aco/U1_7  ( .A(PC_FAIL[7]), .B(n12), .CI(\add_53_aco/carry[7] ), .CO(\add_53_aco/carry[8] ), .S(N53) );
  FA_X1 \add_53_aco/U1_8  ( .A(PC_FAIL[8]), .B(n13), .CI(\add_53_aco/carry[8] ), .CO(\add_53_aco/carry[9] ), .S(N54) );
  FA_X1 \add_53_aco/U1_9  ( .A(PC_FAIL[9]), .B(n14), .CI(\add_53_aco/carry[9] ), .CO(\add_53_aco/carry[10] ), .S(N55) );
  FA_X1 \add_53_aco/U1_10  ( .A(PC_FAIL[10]), .B(n15), .CI(
        \add_53_aco/carry[10] ), .CO(\add_53_aco/carry[11] ), .S(N56) );
  FA_X1 \add_53_aco/U1_11  ( .A(PC_FAIL[11]), .B(n16), .CI(
        \add_53_aco/carry[11] ), .CO(\add_53_aco/carry[12] ), .S(N57) );
  FA_X1 \add_53_aco/U1_12  ( .A(PC_FAIL[12]), .B(n17), .CI(
        \add_53_aco/carry[12] ), .CO(\add_53_aco/carry[13] ), .S(N58) );
  FA_X1 \add_53_aco/U1_13  ( .A(PC_FAIL[13]), .B(n18), .CI(
        \add_53_aco/carry[13] ), .CO(\add_53_aco/carry[14] ), .S(N59) );
  FA_X1 \add_53_aco/U1_14  ( .A(PC_FAIL[14]), .B(n19), .CI(
        \add_53_aco/carry[14] ), .CO(\add_53_aco/carry[15] ), .S(N60) );
  FA_X1 \add_53_aco/U1_15  ( .A(PC_FAIL[15]), .B(n5), .CI(
        \add_53_aco/carry[15] ), .CO(\add_53_aco/carry[16] ), .S(N61) );
  FA_X1 \add_53_aco/U1_16  ( .A(PC_FAIL[16]), .B(n5), .CI(
        \add_53_aco/carry[16] ), .CO(\add_53_aco/carry[17] ), .S(N62) );
  FA_X1 \add_53_aco/U1_17  ( .A(PC_FAIL[17]), .B(n5), .CI(
        \add_53_aco/carry[17] ), .CO(\add_53_aco/carry[18] ), .S(N63) );
  FA_X1 \add_53_aco/U1_18  ( .A(PC_FAIL[18]), .B(n5), .CI(
        \add_53_aco/carry[18] ), .CO(\add_53_aco/carry[19] ), .S(N64) );
  FA_X1 \add_53_aco/U1_19  ( .A(PC_FAIL[19]), .B(n5), .CI(
        \add_53_aco/carry[19] ), .CO(\add_53_aco/carry[20] ), .S(N65) );
  FA_X1 \add_53_aco/U1_20  ( .A(PC_FAIL[20]), .B(n5), .CI(
        \add_53_aco/carry[20] ), .CO(\add_53_aco/carry[21] ), .S(N66) );
  FA_X1 \add_53_aco/U1_21  ( .A(PC_FAIL[21]), .B(n5), .CI(
        \add_53_aco/carry[21] ), .CO(\add_53_aco/carry[22] ), .S(N67) );
  FA_X1 \add_53_aco/U1_22  ( .A(PC_FAIL[22]), .B(n5), .CI(
        \add_53_aco/carry[22] ), .CO(\add_53_aco/carry[23] ), .S(N68) );
  FA_X1 \add_53_aco/U1_23  ( .A(PC_FAIL[23]), .B(n5), .CI(
        \add_53_aco/carry[23] ), .CO(\add_53_aco/carry[24] ), .S(N69) );
  FA_X1 \add_53_aco/U1_24  ( .A(PC_FAIL[24]), .B(n5), .CI(
        \add_53_aco/carry[24] ), .CO(\add_53_aco/carry[25] ), .S(N70) );
  FA_X1 \add_53_aco/U1_25  ( .A(PC_FAIL[25]), .B(n5), .CI(
        \add_53_aco/carry[25] ), .CO(\add_53_aco/carry[26] ), .S(N71) );
  FA_X1 \add_53_aco/U1_26  ( .A(PC_FAIL[26]), .B(n5), .CI(
        \add_53_aco/carry[26] ), .CO(\add_53_aco/carry[27] ), .S(N72) );
  FA_X1 \add_53_aco/U1_27  ( .A(PC_FAIL[27]), .B(n5), .CI(
        \add_53_aco/carry[27] ), .CO(\add_53_aco/carry[28] ), .S(N73) );
  FA_X1 \add_53_aco/U1_28  ( .A(PC_FAIL[28]), .B(n5), .CI(
        \add_53_aco/carry[28] ), .CO(\add_53_aco/carry[29] ), .S(N74) );
  FA_X1 \add_53_aco/U1_29  ( .A(PC_FAIL[29]), .B(n5), .CI(
        \add_53_aco/carry[29] ), .CO(\add_53_aco/carry[30] ), .S(N75) );
  FA_X1 \add_53_aco/U1_30  ( .A(PC_FAIL[30]), .B(n5), .CI(
        \add_53_aco/carry[30] ), .CO(\add_53_aco/carry[31] ), .S(N76) );
  FA_X1 \add_53_aco/U1_31  ( .A(PC_FAIL[31]), .B(n5), .CI(
        \add_53_aco/carry[31] ), .S(N77) );
  NAND2_X1 U3 ( .A1(n5317), .A2(n5225), .ZN(N323) );
  INV_X2 U4 ( .A(n5224), .ZN(n5317) );
  NOR2_X2 U5 ( .A1(n5222), .A2(n5090), .ZN(N644) );
  INV_X2 U6 ( .A(n5090), .ZN(n5089) );
  NOR3_X2 U7 ( .A1(PC_FAIL[4]), .A2(n5143), .A3(n5145), .ZN(n5205) );
  AOI211_X1 U8 ( .C1(n5202), .C2(\CACHE_mem[26][1] ), .A(n5192), .B(n5191), 
        .ZN(n5216) );
  NOR3_X2 U9 ( .A1(PC_FAIL[2]), .A2(PC_FAIL[4]), .A3(n5145), .ZN(n5202) );
  NOR3_X2 U10 ( .A1(PC_FAIL[4]), .A2(PC_FAIL[3]), .A3(n5143), .ZN(n5203) );
  NOR3_X2 U11 ( .A1(PC_FAIL[2]), .A2(PC_FAIL[4]), .A3(PC_FAIL[3]), .ZN(n5207)
         );
  AOI211_X4 U12 ( .C1(n5218), .C2(n5217), .A(n5216), .B(n5215), .ZN(n5236) );
  INV_X1 U13 ( .A(n5202), .ZN(n5178) );
  INV_X1 U14 ( .A(n5203), .ZN(n5179) );
  INV_X1 U15 ( .A(n5207), .ZN(n5181) );
  BUF_X1 U16 ( .A(N356), .Z(n5092) );
  OAI221_X1 U17 ( .B1(n5093), .B2(n5284), .C1(n5093), .C2(n5225), .A(n5090), 
        .ZN(SEL) );
  INV_X1 U18 ( .A(RST), .ZN(n5093) );
  BUF_X1 U19 ( .A(n5316), .Z(n5091) );
  NOR2_X1 U20 ( .A1(n5285), .A2(n5284), .ZN(n5316) );
  OR2_X1 U21 ( .A1(n5094), .A2(n5219), .ZN(n5090) );
  AND2_X1 U22 ( .A1(RST), .A2(n5223), .ZN(N645) );
  INV_X1 U23 ( .A(n5205), .ZN(n5187) );
  INV_X1 U24 ( .A(PC_FAIL[5]), .ZN(n5199) );
  INV_X1 U25 ( .A(RST), .ZN(n5094) );
  INV_X1 U26 ( .A(IR_IN[28]), .ZN(n5095) );
  INV_X1 U27 ( .A(PC_IN[6]), .ZN(n5229) );
  INV_X1 U28 ( .A(PC_IN[3]), .ZN(n5233) );
  AND2_X2 U29 ( .A1(n5236), .A2(IR_FAIL[15]), .ZN(n5) );
  INV_X1 U30 ( .A(PC_FAIL[6]), .ZN(n5200) );
  NOR2_X1 U31 ( .A1(PC_FAIL[2]), .A2(n5144), .ZN(n5206) );
  NOR3_X1 U32 ( .A1(IR_IN[29]), .A2(IR_IN[30]), .A3(IR_IN[31]), .ZN(n5135) );
  NAND3_X1 U33 ( .A1(n5135), .A2(IR_IN[27]), .A3(n5095), .ZN(n5284) );
  INV_X1 U34 ( .A(WRONG_PRE), .ZN(n5219) );
  NAND2_X1 U35 ( .A1(RST), .A2(n5219), .ZN(n5285) );
  INV_X1 U36 ( .A(n5285), .ZN(n5096) );
  NAND2_X1 U37 ( .A1(n5284), .A2(n5096), .ZN(n5224) );
  INV_X1 U38 ( .A(PC_IN[2]), .ZN(n5232) );
  NOR2_X1 U39 ( .A1(n5233), .A2(n5232), .ZN(n5231) );
  INV_X1 U40 ( .A(PC_IN[5]), .ZN(n5138) );
  INV_X1 U41 ( .A(PC_IN[4]), .ZN(n5226) );
  NOR2_X1 U42 ( .A1(n5138), .A2(n5226), .ZN(n5121) );
  NAND2_X1 U43 ( .A1(n5231), .A2(n5121), .ZN(n5230) );
  NOR2_X1 U44 ( .A1(n5230), .A2(n5229), .ZN(n5228) );
  AOI21_X1 U45 ( .B1(\CACHE_mem[31][1] ), .B2(n5228), .A(IR_IN[27]), .ZN(n5134) );
  NAND2_X1 U46 ( .A1(PC_IN[5]), .A2(n5226), .ZN(n5123) );
  INV_X1 U47 ( .A(\CACHE_mem[27][1] ), .ZN(n5186) );
  NOR2_X1 U48 ( .A1(PC_IN[5]), .A2(PC_IN[4]), .ZN(n5126) );
  NOR2_X1 U49 ( .A1(PC_IN[5]), .A2(n5226), .ZN(n5120) );
  AOI22_X1 U50 ( .A1(\CACHE_mem[19][1] ), .A2(n5126), .B1(\CACHE_mem[23][1] ), 
        .B2(n5120), .ZN(n5097) );
  OAI211_X1 U51 ( .C1(n5123), .C2(n5186), .A(PC_IN[6]), .B(n5097), .ZN(n5132)
         );
  INV_X1 U52 ( .A(n5231), .ZN(n5227) );
  INV_X1 U53 ( .A(\CACHE_mem[11][1] ), .ZN(n5099) );
  AOI22_X1 U54 ( .A1(\CACHE_mem[3][1] ), .A2(n5126), .B1(\CACHE_mem[7][1] ), 
        .B2(n5120), .ZN(n5098) );
  OAI211_X1 U55 ( .C1(n5099), .C2(n5123), .A(n5098), .B(n5229), .ZN(n5100) );
  AOI21_X1 U56 ( .B1(\CACHE_mem[15][1] ), .B2(n5121), .A(n5100), .ZN(n5101) );
  NOR2_X1 U57 ( .A1(n5227), .A2(n5101), .ZN(n5131) );
  AOI22_X1 U58 ( .A1(n5121), .A2(\CACHE_mem[30][1] ), .B1(\CACHE_mem[22][1] ), 
        .B2(n5120), .ZN(n5103) );
  INV_X1 U59 ( .A(n5123), .ZN(n5110) );
  AOI22_X1 U60 ( .A1(\CACHE_mem[26][1] ), .A2(n5110), .B1(\CACHE_mem[18][1] ), 
        .B2(n5126), .ZN(n5102) );
  AOI21_X1 U61 ( .B1(n5103), .B2(n5102), .A(n5233), .ZN(n5107) );
  AOI22_X1 U62 ( .A1(n5121), .A2(\CACHE_mem[28][1] ), .B1(\CACHE_mem[20][1] ), 
        .B2(n5120), .ZN(n5105) );
  AOI22_X1 U63 ( .A1(\CACHE_mem[24][1] ), .A2(n5110), .B1(\CACHE_mem[16][1] ), 
        .B2(n5126), .ZN(n5104) );
  AOI21_X1 U64 ( .B1(n5105), .B2(n5104), .A(PC_IN[3]), .ZN(n5106) );
  OAI21_X1 U65 ( .B1(n5107), .B2(n5106), .A(PC_IN[6]), .ZN(n5116) );
  AOI22_X1 U66 ( .A1(n5121), .A2(\CACHE_mem[14][1] ), .B1(\CACHE_mem[6][1] ), 
        .B2(n5120), .ZN(n5109) );
  AOI22_X1 U67 ( .A1(\CACHE_mem[10][1] ), .A2(n5110), .B1(\CACHE_mem[2][1] ), 
        .B2(n5126), .ZN(n5108) );
  AOI21_X1 U68 ( .B1(n5109), .B2(n5108), .A(n5233), .ZN(n5114) );
  AOI22_X1 U69 ( .A1(n5121), .A2(\CACHE_mem[12][1] ), .B1(\CACHE_mem[4][1] ), 
        .B2(n5120), .ZN(n5112) );
  AOI22_X1 U70 ( .A1(\CACHE_mem[8][1] ), .A2(n5110), .B1(\CACHE_mem[0][1] ), 
        .B2(n5126), .ZN(n5111) );
  AOI21_X1 U71 ( .B1(n5112), .B2(n5111), .A(PC_IN[3]), .ZN(n5113) );
  OAI21_X1 U72 ( .B1(n5114), .B2(n5113), .A(n5229), .ZN(n5115) );
  AOI21_X1 U73 ( .B1(n5116), .B2(n5115), .A(PC_IN[2]), .ZN(n5130) );
  INV_X1 U74 ( .A(\CACHE_mem[25][1] ), .ZN(n5118) );
  AOI22_X1 U75 ( .A1(n5121), .A2(\CACHE_mem[29][1] ), .B1(\CACHE_mem[21][1] ), 
        .B2(n5120), .ZN(n5117) );
  OAI211_X1 U76 ( .C1(n5123), .C2(n5118), .A(PC_IN[6]), .B(n5117), .ZN(n5119)
         );
  AOI21_X1 U77 ( .B1(\CACHE_mem[17][1] ), .B2(n5126), .A(n5119), .ZN(n5128) );
  INV_X1 U78 ( .A(\CACHE_mem[9][1] ), .ZN(n5124) );
  AOI22_X1 U79 ( .A1(n5121), .A2(\CACHE_mem[13][1] ), .B1(\CACHE_mem[5][1] ), 
        .B2(n5120), .ZN(n5122) );
  OAI211_X1 U80 ( .C1(n5124), .C2(n5123), .A(n5122), .B(n5229), .ZN(n5125) );
  AOI21_X1 U81 ( .B1(\CACHE_mem[1][1] ), .B2(n5126), .A(n5125), .ZN(n5127) );
  NOR4_X1 U82 ( .A1(PC_IN[3]), .A2(n5128), .A3(n5127), .A4(n5232), .ZN(n5129)
         );
  AOI211_X1 U83 ( .C1(n5132), .C2(n5131), .A(n5130), .B(n5129), .ZN(n5133) );
  NAND4_X1 U84 ( .A1(n5135), .A2(IR_IN[28]), .A3(n5134), .A4(n5133), .ZN(n5225) );
  OAI21_X1 U85 ( .B1(WRONG_PRE), .B2(n5284), .A(RST), .ZN(N356) );
  AND2_X1 U86 ( .A1(RST), .A2(N113), .ZN(N357) );
  AND2_X1 U87 ( .A1(RST), .A2(N114), .ZN(N358) );
  NAND2_X1 U88 ( .A1(n5231), .A2(PC_IN[4]), .ZN(n5137) );
  INV_X1 U89 ( .A(n5230), .ZN(n5136) );
  AOI211_X1 U90 ( .C1(n5138), .C2(n5137), .A(n5136), .B(n5094), .ZN(N362) );
  INV_X1 U91 ( .A(n5228), .ZN(n5250) );
  INV_X1 U92 ( .A(PC_IN[7]), .ZN(n5249) );
  NOR2_X1 U93 ( .A1(n5250), .A2(n5249), .ZN(n5248) );
  NAND2_X1 U94 ( .A1(n5248), .A2(PC_IN[8]), .ZN(n5253) );
  INV_X1 U95 ( .A(PC_IN[9]), .ZN(n5252) );
  NOR2_X1 U96 ( .A1(n5253), .A2(n5252), .ZN(n5251) );
  NAND2_X1 U97 ( .A1(n5251), .A2(PC_IN[10]), .ZN(n5256) );
  INV_X1 U98 ( .A(PC_IN[11]), .ZN(n5255) );
  NOR2_X1 U99 ( .A1(n5256), .A2(n5255), .ZN(n5254) );
  NAND2_X1 U100 ( .A1(n5254), .A2(PC_IN[12]), .ZN(n5259) );
  INV_X1 U101 ( .A(PC_IN[13]), .ZN(n5258) );
  NOR2_X1 U102 ( .A1(n5259), .A2(n5258), .ZN(n5257) );
  NAND2_X1 U103 ( .A1(n5257), .A2(PC_IN[14]), .ZN(n5262) );
  INV_X1 U104 ( .A(PC_IN[15]), .ZN(n5261) );
  NOR2_X1 U105 ( .A1(n5262), .A2(n5261), .ZN(n5260) );
  NAND2_X1 U106 ( .A1(n5260), .A2(PC_IN[16]), .ZN(n5265) );
  INV_X1 U107 ( .A(PC_IN[17]), .ZN(n5264) );
  NOR2_X1 U108 ( .A1(n5265), .A2(n5264), .ZN(n5263) );
  NAND2_X1 U109 ( .A1(n5263), .A2(PC_IN[18]), .ZN(n5268) );
  INV_X1 U110 ( .A(PC_IN[19]), .ZN(n5267) );
  NOR2_X1 U111 ( .A1(n5268), .A2(n5267), .ZN(n5266) );
  NAND2_X1 U112 ( .A1(n5266), .A2(PC_IN[20]), .ZN(n5271) );
  INV_X1 U113 ( .A(PC_IN[21]), .ZN(n5270) );
  NOR2_X1 U114 ( .A1(n5271), .A2(n5270), .ZN(n5269) );
  NAND2_X1 U115 ( .A1(n5269), .A2(PC_IN[22]), .ZN(n5274) );
  INV_X1 U116 ( .A(PC_IN[23]), .ZN(n5273) );
  NOR2_X1 U117 ( .A1(n5274), .A2(n5273), .ZN(n5272) );
  NAND2_X1 U118 ( .A1(n5272), .A2(PC_IN[24]), .ZN(n5277) );
  INV_X1 U119 ( .A(PC_IN[25]), .ZN(n5276) );
  NOR2_X1 U120 ( .A1(n5277), .A2(n5276), .ZN(n5275) );
  NAND2_X1 U121 ( .A1(n5275), .A2(PC_IN[26]), .ZN(n5280) );
  INV_X1 U122 ( .A(PC_IN[27]), .ZN(n5279) );
  NOR2_X1 U123 ( .A1(n5280), .A2(n5279), .ZN(n5278) );
  NAND2_X1 U124 ( .A1(n5278), .A2(PC_IN[28]), .ZN(n5283) );
  INV_X1 U125 ( .A(PC_IN[29]), .ZN(n5282) );
  NOR2_X1 U126 ( .A1(n5283), .A2(n5282), .ZN(n5281) );
  INV_X1 U127 ( .A(n5281), .ZN(n5140) );
  INV_X1 U128 ( .A(PC_IN[30]), .ZN(n5139) );
  NOR2_X1 U129 ( .A1(n5140), .A2(n5139), .ZN(n5142) );
  AOI211_X1 U130 ( .C1(n5140), .C2(n5139), .A(n5142), .B(n5093), .ZN(N387) );
  OAI21_X1 U131 ( .B1(PC_IN[31]), .B2(n5142), .A(RST), .ZN(n5141) );
  AOI21_X1 U132 ( .B1(PC_IN[31]), .B2(n5142), .A(n5141), .ZN(N388) );
  NAND3_X1 U133 ( .A1(PC_FAIL[2]), .A2(PC_FAIL[4]), .A3(PC_FAIL[3]), .ZN(n5174) );
  INV_X1 U134 ( .A(PC_FAIL[2]), .ZN(n5143) );
  INV_X1 U135 ( .A(PC_FAIL[3]), .ZN(n5145) );
  AOI22_X1 U136 ( .A1(n5203), .A2(\CACHE_mem[9][0] ), .B1(n5202), .B2(
        \CACHE_mem[10][0] ), .ZN(n5155) );
  NAND3_X1 U137 ( .A1(n5143), .A2(n5145), .A3(PC_FAIL[4]), .ZN(n5177) );
  INV_X1 U138 ( .A(n5177), .ZN(n5204) );
  AOI22_X1 U139 ( .A1(n5205), .A2(\CACHE_mem[11][0] ), .B1(n5204), .B2(
        \CACHE_mem[12][0] ), .ZN(n5148) );
  NAND2_X1 U140 ( .A1(PC_FAIL[4]), .A2(PC_FAIL[3]), .ZN(n5144) );
  AOI22_X1 U141 ( .A1(n5207), .A2(\CACHE_mem[8][0] ), .B1(n5206), .B2(
        \CACHE_mem[14][0] ), .ZN(n5147) );
  INV_X1 U142 ( .A(n5174), .ZN(n5198) );
  NAND3_X1 U143 ( .A1(n5145), .A2(PC_FAIL[4]), .A3(PC_FAIL[2]), .ZN(n5176) );
  INV_X1 U144 ( .A(n5176), .ZN(n5197) );
  AOI22_X1 U145 ( .A1(n5198), .A2(\CACHE_mem[15][0] ), .B1(n5197), .B2(
        \CACHE_mem[13][0] ), .ZN(n5146) );
  AND4_X1 U146 ( .A1(PC_FAIL[5]), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(
        n5154) );
  AOI22_X1 U147 ( .A1(n5203), .A2(\CACHE_mem[1][0] ), .B1(n5202), .B2(
        \CACHE_mem[2][0] ), .ZN(n5153) );
  AOI22_X1 U148 ( .A1(n5205), .A2(\CACHE_mem[3][0] ), .B1(n5204), .B2(
        \CACHE_mem[4][0] ), .ZN(n5151) );
  AOI22_X1 U149 ( .A1(n5207), .A2(\CACHE_mem[0][0] ), .B1(n5206), .B2(
        \CACHE_mem[6][0] ), .ZN(n5150) );
  AOI22_X1 U150 ( .A1(n5198), .A2(\CACHE_mem[7][0] ), .B1(n5197), .B2(
        \CACHE_mem[5][0] ), .ZN(n5149) );
  AND4_X1 U151 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5199), .ZN(n5152) );
  AOI22_X1 U152 ( .A1(n5155), .A2(n5154), .B1(n5153), .B2(n5152), .ZN(n5167)
         );
  AOI22_X1 U153 ( .A1(n5203), .A2(\CACHE_mem[25][0] ), .B1(n5202), .B2(
        \CACHE_mem[26][0] ), .ZN(n5165) );
  AOI22_X1 U154 ( .A1(n5205), .A2(\CACHE_mem[27][0] ), .B1(n5204), .B2(
        \CACHE_mem[28][0] ), .ZN(n5158) );
  AOI22_X1 U155 ( .A1(n5207), .A2(\CACHE_mem[24][0] ), .B1(n5206), .B2(
        \CACHE_mem[30][0] ), .ZN(n5157) );
  AOI22_X1 U156 ( .A1(n5198), .A2(\CACHE_mem[31][0] ), .B1(n5197), .B2(
        \CACHE_mem[29][0] ), .ZN(n5156) );
  AND4_X1 U157 ( .A1(PC_FAIL[5]), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(
        n5164) );
  AOI22_X1 U158 ( .A1(n5203), .A2(\CACHE_mem[17][0] ), .B1(n5202), .B2(
        \CACHE_mem[18][0] ), .ZN(n5163) );
  AOI22_X1 U159 ( .A1(n5205), .A2(\CACHE_mem[19][0] ), .B1(n5204), .B2(
        \CACHE_mem[20][0] ), .ZN(n5161) );
  AOI22_X1 U160 ( .A1(n5207), .A2(\CACHE_mem[16][0] ), .B1(n5206), .B2(
        \CACHE_mem[22][0] ), .ZN(n5160) );
  AOI22_X1 U161 ( .A1(n5198), .A2(\CACHE_mem[23][0] ), .B1(n5197), .B2(
        \CACHE_mem[21][0] ), .ZN(n5159) );
  AND4_X1 U162 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5199), .ZN(n5162) );
  AOI22_X1 U163 ( .A1(n5165), .A2(n5164), .B1(n5163), .B2(n5162), .ZN(n5166)
         );
  MUX2_X1 U164 ( .A(n5167), .B(n5166), .S(PC_FAIL[6]), .Z(n5222) );
  AOI21_X1 U165 ( .B1(n5222), .B2(RIGHT_PRE), .A(n5089), .ZN(n5169) );
  NOR2_X1 U166 ( .A1(n5169), .A2(n5199), .ZN(n5171) );
  NAND2_X1 U167 ( .A1(PC_FAIL[6]), .A2(n5171), .ZN(n5168) );
  OAI21_X1 U168 ( .B1(n5174), .B2(n5168), .A(RST), .ZN(N612) );
  INV_X1 U169 ( .A(n5206), .ZN(n5175) );
  OAI21_X1 U170 ( .B1(n5175), .B2(n5168), .A(RST), .ZN(N613) );
  OAI21_X1 U171 ( .B1(n5176), .B2(n5168), .A(RST), .ZN(N614) );
  OAI21_X1 U172 ( .B1(n5177), .B2(n5168), .A(RST), .ZN(N615) );
  OAI21_X1 U173 ( .B1(n5187), .B2(n5168), .A(RST), .ZN(N616) );
  OAI21_X1 U174 ( .B1(n5178), .B2(n5168), .A(RST), .ZN(N617) );
  OAI21_X1 U175 ( .B1(n5179), .B2(n5168), .A(RST), .ZN(N618) );
  OAI21_X1 U176 ( .B1(n5181), .B2(n5168), .A(RST), .ZN(N619) );
  NOR2_X1 U177 ( .A1(PC_FAIL[5]), .A2(n5169), .ZN(n5173) );
  NAND2_X1 U178 ( .A1(PC_FAIL[6]), .A2(n5173), .ZN(n5170) );
  OAI21_X1 U179 ( .B1(n5174), .B2(n5170), .A(RST), .ZN(N620) );
  OAI21_X1 U180 ( .B1(n5175), .B2(n5170), .A(RST), .ZN(N621) );
  OAI21_X1 U181 ( .B1(n5176), .B2(n5170), .A(RST), .ZN(N622) );
  OAI21_X1 U182 ( .B1(n5177), .B2(n5170), .A(RST), .ZN(N623) );
  OAI21_X1 U183 ( .B1(n5187), .B2(n5170), .A(RST), .ZN(N624) );
  OAI21_X1 U184 ( .B1(n5178), .B2(n5170), .A(RST), .ZN(N625) );
  OAI21_X1 U185 ( .B1(n5179), .B2(n5170), .A(RST), .ZN(N626) );
  OAI21_X1 U186 ( .B1(n5181), .B2(n5170), .A(RST), .ZN(N627) );
  NAND2_X1 U187 ( .A1(n5171), .A2(n5200), .ZN(n5172) );
  OAI21_X1 U188 ( .B1(n5174), .B2(n5172), .A(RST), .ZN(N628) );
  OAI21_X1 U189 ( .B1(n5175), .B2(n5172), .A(RST), .ZN(N629) );
  OAI21_X1 U190 ( .B1(n5176), .B2(n5172), .A(RST), .ZN(N630) );
  OAI21_X1 U191 ( .B1(n5177), .B2(n5172), .A(RST), .ZN(N631) );
  OAI21_X1 U192 ( .B1(n5187), .B2(n5172), .A(RST), .ZN(N632) );
  OAI21_X1 U193 ( .B1(n5178), .B2(n5172), .A(RST), .ZN(N633) );
  OAI21_X1 U194 ( .B1(n5179), .B2(n5172), .A(RST), .ZN(N634) );
  OAI21_X1 U195 ( .B1(n5181), .B2(n5172), .A(RST), .ZN(N635) );
  NAND2_X1 U196 ( .A1(n5173), .A2(n5200), .ZN(n5180) );
  OAI21_X1 U197 ( .B1(n5174), .B2(n5180), .A(RST), .ZN(N636) );
  OAI21_X1 U198 ( .B1(n5175), .B2(n5180), .A(RST), .ZN(N637) );
  OAI21_X1 U199 ( .B1(n5176), .B2(n5180), .A(RST), .ZN(N638) );
  OAI21_X1 U200 ( .B1(n5177), .B2(n5180), .A(RST), .ZN(N639) );
  OAI21_X1 U201 ( .B1(n5187), .B2(n5180), .A(RST), .ZN(N640) );
  OAI21_X1 U202 ( .B1(n5178), .B2(n5180), .A(RST), .ZN(N641) );
  OAI21_X1 U203 ( .B1(n5179), .B2(n5180), .A(RST), .ZN(N642) );
  OAI21_X1 U204 ( .B1(n5181), .B2(n5180), .A(RST), .ZN(N643) );
  AOI22_X1 U205 ( .A1(n5203), .A2(\CACHE_mem[9][1] ), .B1(n5202), .B2(
        \CACHE_mem[10][1] ), .ZN(n5218) );
  NOR2_X1 U206 ( .A1(PC_FAIL[6]), .A2(n5199), .ZN(n5185) );
  AOI22_X1 U207 ( .A1(n5205), .A2(\CACHE_mem[11][1] ), .B1(n5206), .B2(
        \CACHE_mem[14][1] ), .ZN(n5184) );
  AOI22_X1 U208 ( .A1(n5198), .A2(\CACHE_mem[15][1] ), .B1(n5207), .B2(
        \CACHE_mem[8][1] ), .ZN(n5183) );
  AOI22_X1 U209 ( .A1(n5204), .A2(\CACHE_mem[12][1] ), .B1(n5197), .B2(
        \CACHE_mem[13][1] ), .ZN(n5182) );
  AND4_X1 U210 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n5217) );
  OAI211_X1 U211 ( .C1(n5187), .C2(n5186), .A(PC_FAIL[5]), .B(PC_FAIL[6]), 
        .ZN(n5192) );
  AOI22_X1 U212 ( .A1(n5203), .A2(\CACHE_mem[25][1] ), .B1(n5207), .B2(
        \CACHE_mem[24][1] ), .ZN(n5190) );
  AOI22_X1 U213 ( .A1(n5204), .A2(\CACHE_mem[28][1] ), .B1(n5206), .B2(
        \CACHE_mem[30][1] ), .ZN(n5189) );
  AOI22_X1 U214 ( .A1(n5198), .A2(\CACHE_mem[31][1] ), .B1(n5197), .B2(
        \CACHE_mem[29][1] ), .ZN(n5188) );
  NAND3_X1 U215 ( .A1(n5190), .A2(n5189), .A3(n5188), .ZN(n5191) );
  AOI22_X1 U216 ( .A1(n5202), .A2(\CACHE_mem[18][1] ), .B1(n5207), .B2(
        \CACHE_mem[16][1] ), .ZN(n5193) );
  NAND3_X1 U217 ( .A1(PC_FAIL[6]), .A2(n5193), .A3(n5199), .ZN(n5214) );
  AOI22_X1 U218 ( .A1(n5203), .A2(\CACHE_mem[17][1] ), .B1(n5197), .B2(
        \CACHE_mem[21][1] ), .ZN(n5196) );
  AOI22_X1 U219 ( .A1(n5205), .A2(\CACHE_mem[19][1] ), .B1(n5204), .B2(
        \CACHE_mem[20][1] ), .ZN(n5195) );
  AOI22_X1 U220 ( .A1(n5198), .A2(\CACHE_mem[23][1] ), .B1(n5206), .B2(
        \CACHE_mem[22][1] ), .ZN(n5194) );
  NAND3_X1 U221 ( .A1(n5196), .A2(n5195), .A3(n5194), .ZN(n5213) );
  AOI22_X1 U222 ( .A1(n5198), .A2(\CACHE_mem[7][1] ), .B1(n5197), .B2(
        \CACHE_mem[5][1] ), .ZN(n5201) );
  NAND3_X1 U223 ( .A1(n5201), .A2(n5200), .A3(n5199), .ZN(n5212) );
  AOI22_X1 U224 ( .A1(n5203), .A2(\CACHE_mem[1][1] ), .B1(n5202), .B2(
        \CACHE_mem[2][1] ), .ZN(n5210) );
  AOI22_X1 U225 ( .A1(n5205), .A2(\CACHE_mem[3][1] ), .B1(n5204), .B2(
        \CACHE_mem[4][1] ), .ZN(n5209) );
  AOI22_X1 U226 ( .A1(n5207), .A2(\CACHE_mem[0][1] ), .B1(n5206), .B2(
        \CACHE_mem[6][1] ), .ZN(n5208) );
  NAND3_X1 U227 ( .A1(n5210), .A2(n5209), .A3(n5208), .ZN(n5211) );
  OAI22_X1 U228 ( .A1(n5214), .A2(n5213), .B1(n5212), .B2(n5211), .ZN(n5215)
         );
  NOR2_X1 U229 ( .A1(n5236), .A2(n5219), .ZN(n5221) );
  AOI22_X1 U230 ( .A1(n5236), .A2(n5219), .B1(n5222), .B2(n5221), .ZN(n5220)
         );
  OAI21_X1 U231 ( .B1(n5222), .B2(n5221), .A(n5220), .ZN(n5223) );
  NOR2_X1 U232 ( .A1(n5225), .A2(n5224), .ZN(TAKEN) );
  AND3_X1 U233 ( .A1(n5236), .A2(IR_FAIL[0]), .A3(PC_FAIL[0]), .ZN(
        \add_53_aco/n2 ) );
  AND2_X1 U234 ( .A1(N113), .A2(IR_IN[0]), .ZN(\add_59/n1 ) );
  AND2_X1 U235 ( .A1(n5236), .A2(IR_FAIL[4]), .ZN(n10) );
  AND2_X1 U236 ( .A1(n5236), .A2(IR_FAIL[6]), .ZN(n11) );
  AND2_X1 U237 ( .A1(n5236), .A2(IR_FAIL[7]), .ZN(n12) );
  AND2_X1 U238 ( .A1(n5236), .A2(IR_FAIL[8]), .ZN(n13) );
  AND2_X1 U239 ( .A1(n5236), .A2(IR_FAIL[9]), .ZN(n14) );
  AND2_X1 U240 ( .A1(n5236), .A2(IR_FAIL[10]), .ZN(n15) );
  AND2_X1 U241 ( .A1(n5236), .A2(IR_FAIL[11]), .ZN(n16) );
  AND2_X1 U242 ( .A1(n5236), .A2(IR_FAIL[12]), .ZN(n17) );
  AND2_X1 U243 ( .A1(n5236), .A2(IR_FAIL[13]), .ZN(n18) );
  AND2_X1 U244 ( .A1(n5236), .A2(IR_FAIL[14]), .ZN(n19) );
  AOI221_X1 U245 ( .B1(n5231), .B2(PC_IN[4]), .C1(n5227), .C2(n5226), .A(n5094), .ZN(n286) );
  AOI211_X1 U246 ( .C1(n5230), .C2(n5229), .A(n5228), .B(n5093), .ZN(n291) );
  AOI211_X1 U247 ( .C1(n5233), .C2(n5232), .A(n5231), .B(n5093), .ZN(n59) );
  AND2_X1 U248 ( .A1(n5236), .A2(IR_FAIL[1]), .ZN(n6) );
  NOR2_X1 U249 ( .A1(N113), .A2(IR_IN[0]), .ZN(n5235) );
  AOI21_X1 U250 ( .B1(IR_FAIL[0]), .B2(n5236), .A(PC_FAIL[0]), .ZN(n5234) );
  OAI33_X1 U251 ( .A1(n5285), .A2(\add_59/n1 ), .A3(n5235), .B1(n5090), .B2(
        n5234), .B3(\add_53_aco/n2 ), .ZN(n60) );
  NOR2_X1 U252 ( .A1(PC_IN[2]), .A2(n5093), .ZN(n62) );
  AND2_X1 U253 ( .A1(n5236), .A2(IR_FAIL[5]), .ZN(n7) );
  AND2_X1 U254 ( .A1(n5236), .A2(IR_FAIL[2]), .ZN(n8) );
  AND2_X1 U255 ( .A1(n5236), .A2(IR_FAIL[3]), .ZN(n9) );
  OAI211_X1 U256 ( .C1(n5272), .C2(PC_IN[24]), .A(n5277), .B(RST), .ZN(n5237)
         );
  INV_X1 U257 ( .A(n5237), .ZN(n293) );
  OAI211_X1 U258 ( .C1(n5254), .C2(PC_IN[12]), .A(n5259), .B(RST), .ZN(n5238)
         );
  INV_X1 U259 ( .A(n5238), .ZN(n292) );
  OAI211_X1 U260 ( .C1(n5269), .C2(PC_IN[22]), .A(n5274), .B(RST), .ZN(n5239)
         );
  INV_X1 U261 ( .A(n5239), .ZN(n290) );
  OAI211_X1 U262 ( .C1(n5266), .C2(PC_IN[20]), .A(n5271), .B(RST), .ZN(n5240)
         );
  INV_X1 U263 ( .A(n5240), .ZN(n289) );
  OAI211_X1 U264 ( .C1(n5263), .C2(PC_IN[18]), .A(n5268), .B(RST), .ZN(n5241)
         );
  INV_X1 U265 ( .A(n5241), .ZN(n288) );
  OAI211_X1 U266 ( .C1(n5278), .C2(PC_IN[28]), .A(n5283), .B(RST), .ZN(n5242)
         );
  INV_X1 U267 ( .A(n5242), .ZN(n287) );
  OAI211_X1 U268 ( .C1(n5260), .C2(PC_IN[16]), .A(n5265), .B(RST), .ZN(n5243)
         );
  INV_X1 U269 ( .A(n5243), .ZN(n285) );
  OAI211_X1 U270 ( .C1(n5257), .C2(PC_IN[14]), .A(n5262), .B(RST), .ZN(n5244)
         );
  INV_X1 U271 ( .A(n5244), .ZN(n284) );
  OAI211_X1 U272 ( .C1(n5275), .C2(PC_IN[26]), .A(n5280), .B(RST), .ZN(n5245)
         );
  INV_X1 U273 ( .A(n5245), .ZN(n283) );
  OAI211_X1 U274 ( .C1(n5248), .C2(PC_IN[8]), .A(n5253), .B(RST), .ZN(n5246)
         );
  INV_X1 U275 ( .A(n5246), .ZN(n282) );
  OAI211_X1 U276 ( .C1(n5251), .C2(PC_IN[10]), .A(n5256), .B(RST), .ZN(n5247)
         );
  INV_X1 U277 ( .A(n5247), .ZN(n281) );
  AOI211_X1 U278 ( .C1(n5250), .C2(n5249), .A(n5248), .B(n5093), .ZN(n61) );
  AOI211_X1 U279 ( .C1(n5253), .C2(n5252), .A(n5251), .B(n5093), .ZN(n58) );
  AOI211_X1 U280 ( .C1(n5256), .C2(n5255), .A(n5254), .B(n5093), .ZN(n57) );
  AOI211_X1 U281 ( .C1(n5259), .C2(n5258), .A(n5257), .B(n5093), .ZN(n56) );
  AOI211_X1 U282 ( .C1(n5262), .C2(n5261), .A(n5260), .B(n5093), .ZN(n55) );
  AOI211_X1 U283 ( .C1(n5265), .C2(n5264), .A(n5263), .B(n5094), .ZN(n54) );
  AOI211_X1 U284 ( .C1(n5268), .C2(n5267), .A(n5266), .B(n5094), .ZN(n53) );
  AOI211_X1 U285 ( .C1(n5271), .C2(n5270), .A(n5269), .B(n5094), .ZN(n52) );
  AOI211_X1 U286 ( .C1(n5274), .C2(n5273), .A(n5272), .B(n5094), .ZN(n51) );
  AOI211_X1 U287 ( .C1(n5277), .C2(n5276), .A(n5275), .B(n5094), .ZN(n50) );
  AOI211_X1 U288 ( .C1(n5280), .C2(n5279), .A(n5278), .B(n5094), .ZN(n49) );
  AOI211_X1 U289 ( .C1(n5283), .C2(n5282), .A(n5281), .B(n5093), .ZN(n48) );
  AOI222_X1 U290 ( .A1(n5089), .A2(N47), .B1(n5317), .B2(N220), .C1(n5316), 
        .C2(N82), .ZN(n5286) );
  INV_X1 U291 ( .A(n5286), .ZN(n46) );
  AOI222_X1 U292 ( .A1(n5089), .A2(N48), .B1(n5317), .B2(N221), .C1(n5091), 
        .C2(N83), .ZN(n5287) );
  INV_X1 U293 ( .A(n5287), .ZN(n45) );
  AOI222_X1 U294 ( .A1(n5089), .A2(N49), .B1(n5317), .B2(N222), .C1(n5316), 
        .C2(N84), .ZN(n5288) );
  INV_X1 U295 ( .A(n5288), .ZN(n44) );
  AOI222_X1 U296 ( .A1(n5089), .A2(N50), .B1(n5317), .B2(N223), .C1(n5091), 
        .C2(N85), .ZN(n5289) );
  INV_X1 U297 ( .A(n5289), .ZN(n43) );
  AOI222_X1 U298 ( .A1(n5089), .A2(N51), .B1(n5317), .B2(N224), .C1(n5316), 
        .C2(N86), .ZN(n5290) );
  INV_X1 U299 ( .A(n5290), .ZN(n42) );
  AOI222_X1 U300 ( .A1(n5089), .A2(N52), .B1(n5317), .B2(N225), .C1(n5091), 
        .C2(N87), .ZN(n5291) );
  INV_X1 U301 ( .A(n5291), .ZN(n41) );
  AOI222_X1 U302 ( .A1(n5089), .A2(N53), .B1(n5317), .B2(N226), .C1(n5316), 
        .C2(N88), .ZN(n5292) );
  INV_X1 U303 ( .A(n5292), .ZN(n40) );
  AOI222_X1 U304 ( .A1(n5089), .A2(N54), .B1(n5317), .B2(N227), .C1(n5316), 
        .C2(N89), .ZN(n5293) );
  INV_X1 U305 ( .A(n5293), .ZN(n39) );
  AOI222_X1 U306 ( .A1(n5089), .A2(N55), .B1(n5317), .B2(N228), .C1(n5316), 
        .C2(N90), .ZN(n5294) );
  INV_X1 U307 ( .A(n5294), .ZN(n38) );
  AOI222_X1 U308 ( .A1(n5089), .A2(N56), .B1(n5317), .B2(N229), .C1(n5316), 
        .C2(N91), .ZN(n5295) );
  INV_X1 U309 ( .A(n5295), .ZN(n37) );
  AOI222_X1 U310 ( .A1(n5089), .A2(N57), .B1(n5317), .B2(N230), .C1(n5316), 
        .C2(N92), .ZN(n5296) );
  INV_X1 U311 ( .A(n5296), .ZN(n36) );
  AOI222_X1 U312 ( .A1(n5089), .A2(N58), .B1(n5317), .B2(N231), .C1(n5316), 
        .C2(N93), .ZN(n5297) );
  INV_X1 U313 ( .A(n5297), .ZN(n35) );
  AOI222_X1 U314 ( .A1(n5089), .A2(N59), .B1(n5317), .B2(N232), .C1(n5091), 
        .C2(N94), .ZN(n5298) );
  INV_X1 U315 ( .A(n5298), .ZN(n34) );
  AOI222_X1 U316 ( .A1(n5089), .A2(N60), .B1(n5317), .B2(N233), .C1(n5091), 
        .C2(N95), .ZN(n5299) );
  INV_X1 U317 ( .A(n5299), .ZN(n33) );
  AOI222_X1 U318 ( .A1(n5089), .A2(N61), .B1(n5317), .B2(N234), .C1(n5091), 
        .C2(N96), .ZN(n5300) );
  INV_X1 U319 ( .A(n5300), .ZN(n32) );
  AOI222_X1 U320 ( .A1(n5089), .A2(N62), .B1(n5317), .B2(N235), .C1(n5091), 
        .C2(N97), .ZN(n5301) );
  INV_X1 U321 ( .A(n5301), .ZN(n31) );
  AOI222_X1 U322 ( .A1(n5089), .A2(N63), .B1(n5317), .B2(N236), .C1(n5091), 
        .C2(N98), .ZN(n5302) );
  INV_X1 U323 ( .A(n5302), .ZN(n30) );
  AOI222_X1 U324 ( .A1(n5089), .A2(N64), .B1(n5317), .B2(N237), .C1(n5091), 
        .C2(N99), .ZN(n5303) );
  INV_X1 U325 ( .A(n5303), .ZN(n29) );
  AOI222_X1 U326 ( .A1(n5089), .A2(N65), .B1(n5317), .B2(N238), .C1(n5091), 
        .C2(N100), .ZN(n5304) );
  INV_X1 U327 ( .A(n5304), .ZN(n28) );
  AOI222_X1 U328 ( .A1(n5089), .A2(N66), .B1(n5317), .B2(N239), .C1(n5316), 
        .C2(N101), .ZN(n5305) );
  INV_X1 U329 ( .A(n5305), .ZN(n27) );
  AOI222_X1 U330 ( .A1(n5089), .A2(N67), .B1(n5317), .B2(N240), .C1(n5091), 
        .C2(N102), .ZN(n5306) );
  INV_X1 U331 ( .A(n5306), .ZN(n26) );
  AOI222_X1 U332 ( .A1(n5089), .A2(N68), .B1(n5317), .B2(N241), .C1(n5316), 
        .C2(N103), .ZN(n5307) );
  INV_X1 U333 ( .A(n5307), .ZN(n25) );
  AOI222_X1 U334 ( .A1(n5089), .A2(N69), .B1(n5317), .B2(N242), .C1(n5091), 
        .C2(N104), .ZN(n5308) );
  INV_X1 U335 ( .A(n5308), .ZN(n24) );
  AOI222_X1 U336 ( .A1(n5089), .A2(N70), .B1(n5317), .B2(N243), .C1(n5316), 
        .C2(N105), .ZN(n5309) );
  INV_X1 U337 ( .A(n5309), .ZN(n23) );
  AOI222_X1 U338 ( .A1(n5089), .A2(N71), .B1(n5317), .B2(N244), .C1(n5091), 
        .C2(N106), .ZN(n5310) );
  INV_X1 U339 ( .A(n5310), .ZN(n22) );
  AOI222_X1 U340 ( .A1(n5089), .A2(N72), .B1(n5317), .B2(N245), .C1(n5091), 
        .C2(N107), .ZN(n5311) );
  INV_X1 U341 ( .A(n5311), .ZN(n21) );
  AOI222_X1 U342 ( .A1(n5089), .A2(N73), .B1(n5317), .B2(N246), .C1(n5091), 
        .C2(N108), .ZN(n5312) );
  INV_X1 U343 ( .A(n5312), .ZN(n20) );
  AOI222_X1 U344 ( .A1(n5089), .A2(N74), .B1(n5317), .B2(N247), .C1(n5091), 
        .C2(N109), .ZN(n5313) );
  INV_X1 U345 ( .A(n5313), .ZN(n4) );
  AOI222_X1 U346 ( .A1(n5089), .A2(N75), .B1(n5317), .B2(N248), .C1(n5091), 
        .C2(N110), .ZN(n5314) );
  INV_X1 U347 ( .A(n5314), .ZN(n3) );
  AOI222_X1 U348 ( .A1(n5089), .A2(N76), .B1(n5317), .B2(N249), .C1(n5091), 
        .C2(N111), .ZN(n5315) );
  INV_X1 U349 ( .A(n5315), .ZN(n2) );
  AOI222_X1 U350 ( .A1(n5089), .A2(N77), .B1(n5317), .B2(N250), .C1(n5091), 
        .C2(N112), .ZN(n5318) );
  INV_X1 U351 ( .A(n5318), .ZN(n1) );
endmodule


module DLX_syn ( Clk, Rst, IRAM_DATA_OUT, DRAM_DATA_OUT, DRAM_DATA_IN, 
        DRAM_ADDRESS, DRAM_ENABLE, DRAM_RW, DRAM_SEL, IRAM_ADDRESS );
  input [31:0] IRAM_DATA_OUT;
  input [31:0] DRAM_DATA_OUT;
  output [31:0] DRAM_DATA_IN;
  output [11:0] DRAM_ADDRESS;
  output [2:0] DRAM_SEL;
  output [7:0] IRAM_ADDRESS;
  input Clk, Rst;
  output DRAM_ENABLE, DRAM_RW;
  wire   IR_CU_31, IR_CU_28, IR_CU_27, IR_CU_26, BR_EN_i, \WB_MUX_SEL_i[1] ,
         RF_WE_i, \CU_I/aluOpcode_i[4] , \CU_I/aluOpcode_i[3] ,
         \CU_I/aluOpcode_i[2] , \CU_I/aluOpcode_i[1] , \CU_I/aluOpcode_i[0] ,
         \CU_I/cw2[1] , \CU_I/cw[10] , \CU_I/cw[7] , \CU_I/cw[6] ,
         \CU_I/cw[4] , \CU_I/cw[3] , \CU_I/cw[1] , \CU_I/cw[0] ,
         \DataP/LMD_out[31] , \DataP/LMD_out[30] , \DataP/LMD_out[29] ,
         \DataP/LMD_out[28] , \DataP/LMD_out[27] , \DataP/LMD_out[26] ,
         \DataP/LMD_out[25] , \DataP/LMD_out[24] , \DataP/LMD_out[23] ,
         \DataP/LMD_out[22] , \DataP/LMD_out[21] , \DataP/LMD_out[20] ,
         \DataP/LMD_out[19] , \DataP/LMD_out[18] , \DataP/LMD_out[17] ,
         \DataP/LMD_out[16] , \DataP/LMD_out[15] , \DataP/LMD_out[14] ,
         \DataP/LMD_out[13] , \DataP/LMD_out[12] , \DataP/LMD_out[11] ,
         \DataP/LMD_out[10] , \DataP/LMD_out[9] , \DataP/LMD_out[8] ,
         \DataP/LMD_out[7] , \DataP/LMD_out[6] , \DataP/LMD_out[5] ,
         \DataP/LMD_out[4] , \DataP/LMD_out[3] , \DataP/LMD_out[2] ,
         \DataP/LMD_out[1] , \DataP/LMD_out[0] , \DataP/link_addr_W[31] ,
         \DataP/link_addr_W[30] , \DataP/link_addr_W[29] ,
         \DataP/link_addr_W[28] , \DataP/link_addr_W[27] ,
         \DataP/link_addr_W[26] , \DataP/link_addr_W[25] ,
         \DataP/link_addr_W[24] , \DataP/link_addr_W[23] ,
         \DataP/link_addr_W[22] , \DataP/link_addr_W[21] ,
         \DataP/link_addr_W[20] , \DataP/link_addr_W[19] ,
         \DataP/link_addr_W[18] , \DataP/link_addr_W[17] ,
         \DataP/link_addr_W[16] , \DataP/link_addr_W[15] ,
         \DataP/link_addr_W[14] , \DataP/link_addr_W[13] ,
         \DataP/link_addr_W[12] , \DataP/link_addr_W[11] ,
         \DataP/link_addr_W[10] , \DataP/link_addr_W[9] ,
         \DataP/link_addr_W[8] , \DataP/link_addr_W[7] ,
         \DataP/link_addr_W[6] , \DataP/link_addr_W[5] ,
         \DataP/link_addr_W[4] , \DataP/link_addr_W[3] ,
         \DataP/link_addr_W[2] , \DataP/link_addr_W[1] ,
         \DataP/link_addr_W[0] , \DataP/FWD_MUX_BR_S[1] ,
         \DataP/FWD_MUX_BR_S[0] , \DataP/alu_b_in[31] , \DataP/alu_b_in[30] ,
         \DataP/alu_b_in[29] , \DataP/alu_b_in[28] , \DataP/alu_b_in[27] ,
         \DataP/alu_b_in[26] , \DataP/alu_b_in[24] , \DataP/alu_b_in[23] ,
         \DataP/alu_b_in[22] , \DataP/alu_b_in[21] , \DataP/alu_b_in[20] ,
         \DataP/alu_b_in[19] , \DataP/alu_b_in[18] , \DataP/alu_b_in[17] ,
         \DataP/alu_b_in[16] , \DataP/alu_b_in[15] , \DataP/alu_b_in[13] ,
         \DataP/alu_b_in[12] , \DataP/alu_b_in[11] , \DataP/alu_b_in[10] ,
         \DataP/alu_b_in[9] , \DataP/alu_b_in[8] , \DataP/alu_b_in[7] ,
         \DataP/alu_b_in[6] , \DataP/alu_b_in[3] , \DataP/alu_b_in[2] ,
         \DataP/alu_b_in[1] , \DataP/alu_b_in[0] , \DataP/alu_a_in[31] ,
         \DataP/alu_a_in[30] , \DataP/alu_a_in[29] , \DataP/alu_a_in[28] ,
         \DataP/alu_a_in[27] , \DataP/alu_a_in[26] , \DataP/alu_a_in[25] ,
         \DataP/alu_a_in[24] , \DataP/alu_a_in[23] , \DataP/alu_a_in[22] ,
         \DataP/alu_a_in[21] , \DataP/alu_a_in[20] , \DataP/alu_a_in[19] ,
         \DataP/alu_a_in[18] , \DataP/alu_a_in[17] , \DataP/alu_a_in[16] ,
         \DataP/alu_a_in[15] , \DataP/alu_a_in[14] , \DataP/alu_a_in[13] ,
         \DataP/alu_a_in[12] , \DataP/alu_a_in[11] , \DataP/alu_a_in[10] ,
         \DataP/alu_a_in[9] , \DataP/alu_a_in[8] , \DataP/alu_a_in[7] ,
         \DataP/alu_a_in[6] , \DataP/alu_a_in[5] , \DataP/alu_a_in[4] ,
         \DataP/alu_a_in[3] , \DataP/alu_a_in[2] , \DataP/alu_a_in[0] ,
         \DataP/alu_out_W[0] , \DataP/alu_out_W[1] , \DataP/alu_out_W[2] ,
         \DataP/alu_out_W[3] , \DataP/alu_out_W[4] , \DataP/alu_out_W[5] ,
         \DataP/alu_out_W[6] , \DataP/alu_out_W[7] , \DataP/alu_out_W[8] ,
         \DataP/alu_out_W[9] , \DataP/alu_out_W[10] , \DataP/alu_out_W[11] ,
         \DataP/alu_out_W[12] , \DataP/alu_out_W[13] , \DataP/alu_out_W[14] ,
         \DataP/alu_out_W[15] , \DataP/alu_out_W[16] , \DataP/alu_out_W[17] ,
         \DataP/alu_out_W[18] , \DataP/alu_out_W[19] , \DataP/alu_out_W[20] ,
         \DataP/alu_out_W[21] , \DataP/alu_out_W[22] , \DataP/alu_out_W[23] ,
         \DataP/alu_out_W[24] , \DataP/alu_out_W[25] , \DataP/alu_out_W[26] ,
         \DataP/alu_out_W[27] , \DataP/alu_out_W[28] , \DataP/alu_out_W[29] ,
         \DataP/alu_out_W[30] , \DataP/alu_out_W[31] , \DataP/alu_out_M[12] ,
         \DataP/alu_out_M[13] , \DataP/alu_out_M[14] , \DataP/alu_out_M[15] ,
         \DataP/alu_out_M[16] , \DataP/alu_out_M[17] , \DataP/alu_out_M[18] ,
         \DataP/alu_out_M[19] , \DataP/alu_out_M[20] , \DataP/alu_out_M[21] ,
         \DataP/alu_out_M[22] , \DataP/alu_out_M[23] , \DataP/alu_out_M[24] ,
         \DataP/alu_out_M[25] , \DataP/alu_out_M[26] , \DataP/alu_out_M[27] ,
         \DataP/alu_out_M[28] , \DataP/alu_out_M[29] , \DataP/alu_out_M[30] ,
         \DataP/alu_out_M[31] , \DataP/opcode_W[0] , \DataP/opcode_W[1] ,
         \DataP/opcode_W[2] , \DataP/opcode_W[3] , \DataP/opcode_W[4] ,
         \DataP/opcode_W[5] , \DataP/opcode_M[0] , \DataP/opcode_M[1] ,
         \DataP/opcode_M[2] , \DataP/opcode_M[3] , \DataP/opcode_M[4] ,
         \DataP/dest_M[0] , \DataP/dest_M[1] , \DataP/dest_M[2] ,
         \DataP/dest_M[3] , \DataP/dest_M[4] , \DataP/pr_E ,
         \DataP/opcode_E[0] , \DataP/opcode_E[1] , \DataP/opcode_E[3] ,
         \DataP/opcode_E[4] , \DataP/Rs2[4] , \DataP/Rs2[3] , \DataP/Rs2[2] ,
         \DataP/Rs2[1] , \DataP/Rs2[0] , \DataP/Rs1[1] , \DataP/Rs1[2] ,
         \DataP/IMM_s[30] , \DataP/IMM_s[24] , \DataP/IMM_s[23] ,
         \DataP/IMM_s[22] , \DataP/IMM_s[21] , \DataP/IMM_s[20] ,
         \DataP/IMM_s[19] , \DataP/IMM_s[18] , \DataP/IMM_s[17] ,
         \DataP/IMM_s[16] , \DataP/IMM_s[15] , \DataP/IMM_s[14] ,
         \DataP/IMM_s[13] , \DataP/IMM_s[12] , \DataP/IMM_s[11] ,
         \DataP/IMM_s[10] , \DataP/IMM_s[9] , \DataP/IMM_s[8] ,
         \DataP/IMM_s[7] , \DataP/IMM_s[6] , \DataP/IMM_s[5] ,
         \DataP/IMM_s[4] , \DataP/IMM_s[3] , \DataP/IMM_s[2] ,
         \DataP/IMM_s[1] , \DataP/IMM_s[0] , \DataP/B_s[0] , \DataP/B_s[1] ,
         \DataP/B_s[2] , \DataP/B_s[3] , \DataP/B_s[4] , \DataP/B_s[5] ,
         \DataP/B_s[6] , \DataP/B_s[7] , \DataP/B_s[8] , \DataP/B_s[9] ,
         \DataP/B_s[10] , \DataP/B_s[11] , \DataP/B_s[12] , \DataP/B_s[13] ,
         \DataP/B_s[14] , \DataP/B_s[15] , \DataP/B_s[16] , \DataP/B_s[17] ,
         \DataP/B_s[18] , \DataP/B_s[19] , \DataP/B_s[20] , \DataP/B_s[21] ,
         \DataP/B_s[22] , \DataP/B_s[23] , \DataP/B_s[24] , \DataP/B_s[25] ,
         \DataP/B_s[26] , \DataP/B_s[27] , \DataP/B_s[28] , \DataP/B_s[29] ,
         \DataP/B_s[30] , \DataP/B_s[31] , \DataP/A_s[0] , \DataP/A_s[1] ,
         \DataP/A_s[2] , \DataP/A_s[3] , \DataP/A_s[4] , \DataP/A_s[5] ,
         \DataP/A_s[6] , \DataP/A_s[7] , \DataP/A_s[8] , \DataP/A_s[9] ,
         \DataP/A_s[10] , \DataP/A_s[11] , \DataP/A_s[12] , \DataP/A_s[13] ,
         \DataP/A_s[14] , \DataP/A_s[15] , \DataP/A_s[16] , \DataP/A_s[17] ,
         \DataP/A_s[18] , \DataP/A_s[19] , \DataP/A_s[20] , \DataP/A_s[21] ,
         \DataP/A_s[22] , \DataP/A_s[23] , \DataP/A_s[24] , \DataP/A_s[25] ,
         \DataP/A_s[26] , \DataP/A_s[27] , \DataP/A_s[28] , \DataP/A_s[29] ,
         \DataP/A_s[30] , \DataP/A_s[31] , \DataP/npc_E[9] ,
         \DataP/imm_out[31] , \DataP/imm_out[24] , \DataP/imm_out[23] ,
         \DataP/imm_out[22] , \DataP/imm_out[21] , \DataP/imm_out[20] ,
         \DataP/imm_out[19] , \DataP/imm_out[18] , \DataP/imm_out[17] ,
         \DataP/imm_out[16] , \DataP/b_out[31] , \DataP/b_out[30] ,
         \DataP/b_out[29] , \DataP/b_out[28] , \DataP/b_out[27] ,
         \DataP/b_out[26] , \DataP/b_out[25] , \DataP/b_out[24] ,
         \DataP/b_out[23] , \DataP/b_out[22] , \DataP/b_out[21] ,
         \DataP/b_out[20] , \DataP/b_out[19] , \DataP/b_out[18] ,
         \DataP/b_out[17] , \DataP/b_out[16] , \DataP/b_out[15] ,
         \DataP/b_out[14] , \DataP/b_out[13] , \DataP/b_out[12] ,
         \DataP/b_out[11] , \DataP/b_out[10] , \DataP/b_out[9] ,
         \DataP/b_out[8] , \DataP/b_out[7] , \DataP/b_out[6] ,
         \DataP/b_out[5] , \DataP/b_out[4] , \DataP/b_out[3] ,
         \DataP/b_out[2] , \DataP/b_out[1] , \DataP/b_out[0] ,
         \DataP/a_out[31] , \DataP/a_out[30] , \DataP/a_out[29] ,
         \DataP/a_out[28] , \DataP/a_out[27] , \DataP/a_out[26] ,
         \DataP/a_out[25] , \DataP/a_out[24] , \DataP/a_out[23] ,
         \DataP/a_out[22] , \DataP/a_out[21] , \DataP/a_out[20] ,
         \DataP/a_out[19] , \DataP/a_out[18] , \DataP/a_out[17] ,
         \DataP/a_out[16] , \DataP/a_out[15] , \DataP/a_out[14] ,
         \DataP/a_out[13] , \DataP/a_out[12] , \DataP/a_out[11] ,
         \DataP/a_out[10] , \DataP/a_out[9] , \DataP/a_out[8] ,
         \DataP/a_out[7] , \DataP/a_out[6] , \DataP/a_out[5] ,
         \DataP/a_out[4] , \DataP/a_out[3] , \DataP/a_out[2] ,
         \DataP/a_out[1] , \DataP/a_out[0] , \DataP/WB[31] , \DataP/WB[30] ,
         \DataP/WB[29] , \DataP/WB[28] , \DataP/WB[27] , \DataP/WB[26] ,
         \DataP/WB[25] , \DataP/WB[24] , \DataP/WB[23] , \DataP/WB[22] ,
         \DataP/WB[21] , \DataP/WB[20] , \DataP/WB[19] , \DataP/WB[18] ,
         \DataP/WB[17] , \DataP/WB[16] , \DataP/WB[15] , \DataP/WB[14] ,
         \DataP/WB[13] , \DataP/WB[12] , \DataP/WB[11] , \DataP/WB[10] ,
         \DataP/WB[9] , \DataP/WB[8] , \DataP/WB[7] , \DataP/WB[6] ,
         \DataP/WB[5] , \DataP/WB[4] , \DataP/WB[3] , \DataP/WB[2] ,
         \DataP/WB[1] , \DataP/WB[0] , \DataP/add_D[0] , \DataP/add_D[1] ,
         \DataP/add_D[2] , \DataP/add_D[3] , \DataP/add_D[4] ,
         \DataP/dest_D[4] , \DataP/dest_D[3] , \DataP/dest_D[2] ,
         \DataP/dest_D[1] , \DataP/dest_D[0] , \DataP/add_S2[0] ,
         \DataP/add_S2[1] , \DataP/add_S2[2] , \DataP/add_S2[3] ,
         \DataP/add_S2[4] , \DataP/pr_D , \DataP/link_addr_D[31] ,
         \DataP/link_addr_D[30] , \DataP/link_addr_D[29] ,
         \DataP/link_addr_D[28] , \DataP/link_addr_D[27] ,
         \DataP/link_addr_D[26] , \DataP/link_addr_D[25] ,
         \DataP/link_addr_D[24] , \DataP/link_addr_D[23] ,
         \DataP/link_addr_D[22] , \DataP/link_addr_D[21] ,
         \DataP/link_addr_D[20] , \DataP/link_addr_D[19] ,
         \DataP/link_addr_D[18] , \DataP/link_addr_D[17] ,
         \DataP/link_addr_D[16] , \DataP/link_addr_D[15] ,
         \DataP/link_addr_D[14] , \DataP/link_addr_D[13] ,
         \DataP/link_addr_D[12] , \DataP/link_addr_D[11] ,
         \DataP/link_addr_D[10] , \DataP/link_addr_D[9] ,
         \DataP/link_addr_D[8] , \DataP/link_addr_D[7] ,
         \DataP/link_addr_D[6] , \DataP/link_addr_D[5] ,
         \DataP/link_addr_D[4] , \DataP/link_addr_D[3] ,
         \DataP/link_addr_D[2] , \DataP/link_addr_D[1] ,
         \DataP/link_addr_D[0] , \DataP/prediction , \DataP/npc_mux_sel ,
         \DataP/link_addr_F[31] , \DataP/link_addr_F[30] ,
         \DataP/link_addr_F[29] , \DataP/link_addr_F[28] ,
         \DataP/link_addr_F[27] , \DataP/link_addr_F[26] ,
         \DataP/link_addr_F[25] , \DataP/link_addr_F[24] ,
         \DataP/link_addr_F[23] , \DataP/link_addr_F[22] ,
         \DataP/link_addr_F[21] , \DataP/link_addr_F[20] ,
         \DataP/link_addr_F[19] , \DataP/link_addr_F[18] ,
         \DataP/link_addr_F[17] , \DataP/link_addr_F[16] ,
         \DataP/link_addr_F[15] , \DataP/link_addr_F[14] ,
         \DataP/link_addr_F[13] , \DataP/link_addr_F[12] ,
         \DataP/link_addr_F[11] , \DataP/link_addr_F[10] ,
         \DataP/link_addr_F[9] , \DataP/link_addr_F[8] ,
         \DataP/link_addr_F[7] , \DataP/link_addr_F[6] ,
         \DataP/link_addr_F[5] , \DataP/link_addr_F[4] ,
         \DataP/link_addr_F[3] , \DataP/link_addr_F[2] ,
         \DataP/link_addr_F[1] , \DataP/link_addr_F[0] , \DataP/npc_pre[31] ,
         \DataP/npc_pre[30] , \DataP/npc_pre[29] , \DataP/npc_pre[28] ,
         \DataP/npc_pre[27] , \DataP/npc_pre[26] , \DataP/npc_pre[25] ,
         \DataP/npc_pre[24] , \DataP/npc_pre[23] , \DataP/npc_pre[22] ,
         \DataP/npc_pre[21] , \DataP/npc_pre[20] , \DataP/npc_pre[19] ,
         \DataP/npc_pre[18] , \DataP/npc_pre[17] , \DataP/npc_pre[16] ,
         \DataP/npc_pre[15] , \DataP/npc_pre[14] , \DataP/npc_pre[13] ,
         \DataP/npc_pre[12] , \DataP/npc_pre[11] , \DataP/npc_pre[10] ,
         \DataP/npc_pre[9] , \DataP/npc_pre[8] , \DataP/npc_pre[7] ,
         \DataP/npc_pre[6] , \DataP/npc_pre[5] , \DataP/npc_pre[4] ,
         \DataP/npc_pre[3] , \DataP/npc_pre[2] , \DataP/npc_pre[1] ,
         \DataP/npc_pre[0] , \DataP/right_br , \DataP/wrong_br ,
         \DataP/npc_M[31] , \DataP/npc_M[30] , \DataP/npc_M[29] ,
         \DataP/npc_M[28] , \DataP/npc_M[27] , \DataP/npc_M[26] ,
         \DataP/npc_M[25] , \DataP/npc_M[24] , \DataP/npc_M[23] ,
         \DataP/npc_M[22] , \DataP/npc_M[21] , \DataP/npc_M[20] ,
         \DataP/npc_M[19] , \DataP/npc_M[18] , \DataP/npc_M[17] ,
         \DataP/npc_M[16] , \DataP/npc_M[15] , \DataP/npc_M[14] ,
         \DataP/npc_M[13] , \DataP/npc_M[12] , \DataP/npc_M[11] ,
         \DataP/npc_M[10] , \DataP/npc_M[9] , \DataP/npc_M[8] ,
         \DataP/npc_M[7] , \DataP/npc_M[6] , \DataP/npc_M[5] ,
         \DataP/npc_M[4] , \DataP/npc_M[3] , \DataP/npc_M[2] ,
         \DataP/npc_M[1] , \DataP/npc_M[0] , \DataP/pc_out_0 ,
         \DataP/pc_out_1 , \DataP/pc_out[10] , \DataP/pc_out[11] ,
         \DataP/pc_out[12] , \DataP/pc_out[13] , \DataP/pc_out[14] ,
         \DataP/pc_out[15] , \DataP/pc_out[16] , \DataP/pc_out[17] ,
         \DataP/pc_out[18] , \DataP/pc_out[19] , \DataP/pc_out[20] ,
         \DataP/pc_out[21] , \DataP/pc_out[22] , \DataP/pc_out[23] ,
         \DataP/pc_out[24] , \DataP/pc_out[25] , \DataP/pc_out[26] ,
         \DataP/pc_out[27] , \DataP/pc_out[28] , \DataP/pc_out[29] ,
         \DataP/pc_out[30] , \DataP/pc_out[31] , \DataP/npc[0] ,
         \DataP/npc[1] , \DataP/npc[2] , \DataP/npc[3] , \DataP/npc[4] ,
         \DataP/npc[5] , \DataP/npc[6] , \DataP/npc[7] , \DataP/npc[8] ,
         \DataP/npc[9] , \DataP/npc[10] , \DataP/npc[11] , \DataP/npc[12] ,
         \DataP/npc[13] , \DataP/npc[14] , \DataP/npc[15] , \DataP/npc[16] ,
         \DataP/npc[17] , \DataP/npc[18] , \DataP/npc[19] , \DataP/npc[20] ,
         \DataP/npc[21] , \DataP/npc[22] , \DataP/npc[23] , \DataP/npc[24] ,
         \DataP/npc[25] , \DataP/npc[26] , \DataP/npc[27] , \DataP/npc[28] ,
         \DataP/npc[29] , \DataP/npc[30] , \DataP/npc[31] , \DataP/IR1[11] ,
         \DataP/IR1[12] , \DataP/IR1[13] , \DataP/IR1[14] , \DataP/IR1[15] ,
         \DataP/IR1[21] , \DataP/IR1[22] , \DataP/IR1[23] , \DataP/IR1[24] ,
         \DataP/IR1[25] , \DataP/PC_reg/N33 , \DataP/PC_reg/N32 ,
         \DataP/PC_reg/N31 , \DataP/PC_reg/N30 , \DataP/PC_reg/N29 ,
         \DataP/PC_reg/N28 , \DataP/PC_reg/N27 , \DataP/PC_reg/N26 ,
         \DataP/PC_reg/N25 , \DataP/PC_reg/N24 , \DataP/PC_reg/N23 ,
         \DataP/PC_reg/N22 , \DataP/PC_reg/N21 , \DataP/PC_reg/N20 ,
         \DataP/PC_reg/N19 , \DataP/PC_reg/N18 , \DataP/PC_reg/N17 ,
         \DataP/PC_reg/N16 , \DataP/PC_reg/N15 , \DataP/PC_reg/N14 ,
         \DataP/PC_reg/N13 , \DataP/PC_reg/N12 , \DataP/PC_reg/N11 ,
         \DataP/PC_reg/N10 , \DataP/PC_reg/N9 , \DataP/PC_reg/N8 ,
         \DataP/PC_reg/N7 , \DataP/PC_reg/N6 , \DataP/PC_reg/N5 ,
         \DataP/PC_reg/N4 , \DataP/PC_reg/N3 , \DataP/PC_reg/N2 ,
         \DataP/NPC_add/N32 , \DataP/NPC_add/N31 , \DataP/NPC_add/N30 ,
         \DataP/NPC_add/N29 , \DataP/NPC_add/N28 , \DataP/NPC_add/N27 ,
         \DataP/NPC_add/N26 , \DataP/NPC_add/N25 , \DataP/NPC_add/N24 ,
         \DataP/NPC_add/N23 , \DataP/NPC_add/N22 , \DataP/NPC_add/N21 ,
         \DataP/NPC_add/N20 , \DataP/NPC_add/N19 , \DataP/NPC_add/N18 ,
         \DataP/NPC_add/N17 , \DataP/NPC_add/N16 , \DataP/NPC_add/N15 ,
         \DataP/NPC_add/N14 , \DataP/NPC_add/N13 , \DataP/NPC_add/N12 ,
         \DataP/NPC_add/N11 , \DataP/NPC_add/N10 , \DataP/NPC_add/N9 ,
         \DataP/NPC_add/N8 , \DataP/NPC_add/N7 , \DataP/NPC_add/N6 ,
         \DataP/NPC_add/N5 , \DataP/NPC_add/N4 , \DataP/NPC_add/N3 ,
         \DataP/NPC_add/N2 , \DataP/NPC_add/N1 , \DataP/NPC_add/N0 ,
         \DataP/FORWARDING_BR/N12 , \DataP/ALU_C/shifter/N108 ,
         \DataP/ALU_C/shifter/N107 , \DataP/ALU_C/shifter/N106 ,
         \DataP/ALU_C/shifter/N105 , \DataP/ALU_C/shifter/N104 ,
         \DataP/ALU_C/shifter/N103 , \DataP/ALU_C/shifter/N102 ,
         \DataP/ALU_C/shifter/N101 , \DataP/ALU_C/shifter/N100 ,
         \DataP/ALU_C/shifter/N99 , \DataP/ALU_C/shifter/N97 ,
         \DataP/ALU_C/shifter/N96 , \DataP/ALU_C/shifter/N93 ,
         \DataP/ALU_C/shifter/N84 , \DataP/ALU_C/shifter/N83 ,
         \DataP/ALU_C/shifter/N82 , \DataP/ALU_C/shifter/N81 ,
         \DataP/ALU_C/shifter/N80 , \DataP/ALU_C/shifter/N79 ,
         \DataP/ALU_C/shifter/N78 , \DataP/ALU_C/shifter/N77 ,
         \DataP/ALU_C/shifter/N76 , \DataP/ALU_C/shifter/N75 ,
         \DataP/ALU_C/shifter/N74 , \DataP/ALU_C/shifter/N73 ,
         \DataP/ALU_C/shifter/N72 , \DataP/ALU_C/shifter/N71 ,
         \DataP/ALU_C/shifter/N70 , \DataP/ALU_C/shifter/N69 ,
         \DataP/ALU_C/shifter/N67 , \DataP/ALU_C/shifter/N66 ,
         \DataP/ALU_C/shifter/N65 , \DataP/ALU_C/shifter/N64 ,
         \DataP/ALU_C/shifter/N61 , \DataP/ALU_C/shifter/N59 ,
         \DataP/ALU_C/shifter/N52 , \DataP/ALU_C/shifter/N51 ,
         \DataP/ALU_C/shifter/N50 , \DataP/ALU_C/shifter/N49 ,
         \DataP/ALU_C/shifter/N47 , \DataP/ALU_C/shifter/N46 ,
         \DataP/ALU_C/shifter/N45 , \DataP/ALU_C/shifter/N43 ,
         \DataP/ALU_C/shifter/N42 , \DataP/ALU_C/shifter/N41 ,
         \DataP/ALU_C/shifter/N40 , \DataP/ALU_C/shifter/N39 ,
         \DataP/ALU_C/shifter/N38 , \DataP/ALU_C/shifter/N37 ,
         \DataP/ALU_C/shifter/N36 , \DataP/ALU_C/shifter/N34 ,
         \DataP/ALU_C/shifter/N33 , \DataP/ALU_C/shifter/N32 ,
         \DataP/ALU_C/shifter/N29 , \DataP/ALU_C/shifter/N20 ,
         \DataP/ALU_C/shifter/N19 , \DataP/ALU_C/comp/N50 ,
         \DataP/ALU_C/comp/N24 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n294, n296, n297,
         n299, n300, n301, n303, n304, n308, n311, n313, n317, n319, n322,
         n323, n326, n330, n332, n333, n337, n340, n341, n345, n350, n353,
         n354, n355, n356, n357, n358, n399, n432, n443, n476, n477, n478,
         n479, n480, n482, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n497, n504, n514, n515, n516, n520, n521, n523,
         n524, n528, n529, n530, n536, n538, n540, n607, n1358, n1372, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, \sra_131/SH[4] , \lt_x_135/B[12] , \lt_x_135/B[5] ,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223;
  wire   [10:0] IR_CU;
  wire   [4:0] ALU_OPCODE_i;

  register_file_N32_addBit5 \DataP/Reg_F  ( .RESET(Rst), .RE(1'b1), .WE(
        RF_WE_i), .ADD_WR({n1629, n2146, \DataP/add_D[2] , n2229, 
        \DataP/add_D[0] }), .ADD_RDA({n494, n493, n492, n491, n490}), 
        .ADD_RDB({\DataP/add_S2[4] , \DataP/add_S2[3] , \DataP/add_S2[2] , 
        \DataP/add_S2[1] , \DataP/add_S2[0] }), .DATAIN({\DataP/WB[31] , 
        \DataP/WB[30] , \DataP/WB[29] , \DataP/WB[28] , \DataP/WB[27] , 
        \DataP/WB[26] , \DataP/WB[25] , \DataP/WB[24] , \DataP/WB[23] , 
        \DataP/WB[22] , \DataP/WB[21] , \DataP/WB[20] , \DataP/WB[19] , 
        \DataP/WB[18] , \DataP/WB[17] , \DataP/WB[16] , \DataP/WB[15] , 
        \DataP/WB[14] , \DataP/WB[13] , \DataP/WB[12] , \DataP/WB[11] , 
        \DataP/WB[10] , \DataP/WB[9] , \DataP/WB[8] , \DataP/WB[7] , 
        \DataP/WB[6] , \DataP/WB[5] , \DataP/WB[4] , \DataP/WB[3] , 
        \DataP/WB[2] , \DataP/WB[1] , \DataP/WB[0] }), .OUTA({
        \DataP/a_out[31] , \DataP/a_out[30] , \DataP/a_out[29] , 
        \DataP/a_out[28] , \DataP/a_out[27] , \DataP/a_out[26] , 
        \DataP/a_out[25] , \DataP/a_out[24] , \DataP/a_out[23] , 
        \DataP/a_out[22] , \DataP/a_out[21] , \DataP/a_out[20] , 
        \DataP/a_out[19] , \DataP/a_out[18] , \DataP/a_out[17] , 
        \DataP/a_out[16] , \DataP/a_out[15] , \DataP/a_out[14] , 
        \DataP/a_out[13] , \DataP/a_out[12] , \DataP/a_out[11] , 
        \DataP/a_out[10] , \DataP/a_out[9] , \DataP/a_out[8] , 
        \DataP/a_out[7] , \DataP/a_out[6] , \DataP/a_out[5] , \DataP/a_out[4] , 
        \DataP/a_out[3] , \DataP/a_out[2] , \DataP/a_out[1] , \DataP/a_out[0] }), .OUTB({\DataP/b_out[31] , \DataP/b_out[30] , \DataP/b_out[29] , 
        \DataP/b_out[28] , \DataP/b_out[27] , \DataP/b_out[26] , 
        \DataP/b_out[25] , \DataP/b_out[24] , \DataP/b_out[23] , 
        \DataP/b_out[22] , \DataP/b_out[21] , \DataP/b_out[20] , 
        \DataP/b_out[19] , \DataP/b_out[18] , \DataP/b_out[17] , 
        \DataP/b_out[16] , \DataP/b_out[15] , \DataP/b_out[14] , 
        \DataP/b_out[13] , \DataP/b_out[12] , \DataP/b_out[11] , 
        \DataP/b_out[10] , \DataP/b_out[9] , \DataP/b_out[8] , 
        \DataP/b_out[7] , \DataP/b_out[6] , \DataP/b_out[5] , \DataP/b_out[4] , 
        \DataP/b_out[3] , \DataP/b_out[2] , \DataP/b_out[1] , \DataP/b_out[0] }) );
  branch_predictor \DataP/BR_pred  ( .RST(Rst), .PC_IN({\DataP/pc_out[31] , 
        \DataP/pc_out[30] , \DataP/pc_out[29] , \DataP/pc_out[28] , 
        \DataP/pc_out[27] , \DataP/pc_out[26] , \DataP/pc_out[25] , 
        \DataP/pc_out[24] , \DataP/pc_out[23] , \DataP/pc_out[22] , 
        \DataP/pc_out[21] , \DataP/pc_out[20] , \DataP/pc_out[19] , 
        \DataP/pc_out[18] , \DataP/pc_out[17] , \DataP/pc_out[16] , 
        \DataP/pc_out[15] , \DataP/pc_out[14] , \DataP/pc_out[13] , 
        \DataP/pc_out[12] , \DataP/pc_out[11] , \DataP/pc_out[10] , 
        IRAM_ADDRESS, \DataP/pc_out_1 , \DataP/pc_out_0 }), .PC_FAIL({
        \DataP/npc_M[31] , \DataP/npc_M[30] , \DataP/npc_M[29] , 
        \DataP/npc_M[28] , \DataP/npc_M[27] , \DataP/npc_M[26] , 
        \DataP/npc_M[25] , \DataP/npc_M[24] , \DataP/npc_M[23] , 
        \DataP/npc_M[22] , \DataP/npc_M[21] , \DataP/npc_M[20] , 
        \DataP/npc_M[19] , \DataP/npc_M[18] , \DataP/npc_M[17] , 
        \DataP/npc_M[16] , \DataP/npc_M[15] , \DataP/npc_M[14] , 
        \DataP/npc_M[13] , \DataP/npc_M[12] , \DataP/npc_M[11] , 
        \DataP/npc_M[10] , \DataP/npc_M[9] , \DataP/npc_M[8] , 
        \DataP/npc_M[7] , \DataP/npc_M[6] , \DataP/npc_M[5] , \DataP/npc_M[4] , 
        \DataP/npc_M[3] , \DataP/npc_M[2] , \DataP/npc_M[1] , \DataP/npc_M[0] }), .IR_IN({IRAM_DATA_OUT[31:27], 1'b0, IRAM_DATA_OUT[25:0]}), .IR_FAIL({
        \DataP/IMM_s[15] , \DataP/IMM_s[14] , \DataP/IMM_s[13] , 
        \DataP/IMM_s[12] , \DataP/IMM_s[11] , \DataP/IMM_s[10] , 
        \DataP/IMM_s[9] , \DataP/IMM_s[8] , \DataP/IMM_s[7] , \DataP/IMM_s[6] , 
        \DataP/IMM_s[5] , \DataP/IMM_s[4] , \DataP/IMM_s[3] , \DataP/IMM_s[2] , 
        \DataP/IMM_s[1] , \DataP/IMM_s[0] }), .WRONG_PRE(\DataP/wrong_br ), 
        .RIGHT_PRE(\DataP/right_br ), .NPC_OUT({\DataP/npc_pre[31] , 
        \DataP/npc_pre[30] , \DataP/npc_pre[29] , \DataP/npc_pre[28] , 
        \DataP/npc_pre[27] , \DataP/npc_pre[26] , \DataP/npc_pre[25] , 
        \DataP/npc_pre[24] , \DataP/npc_pre[23] , \DataP/npc_pre[22] , 
        \DataP/npc_pre[21] , \DataP/npc_pre[20] , \DataP/npc_pre[19] , 
        \DataP/npc_pre[18] , \DataP/npc_pre[17] , \DataP/npc_pre[16] , 
        \DataP/npc_pre[15] , \DataP/npc_pre[14] , \DataP/npc_pre[13] , 
        \DataP/npc_pre[12] , \DataP/npc_pre[11] , \DataP/npc_pre[10] , 
        \DataP/npc_pre[9] , \DataP/npc_pre[8] , \DataP/npc_pre[7] , 
        \DataP/npc_pre[6] , \DataP/npc_pre[5] , \DataP/npc_pre[4] , 
        \DataP/npc_pre[3] , \DataP/npc_pre[2] , \DataP/npc_pre[1] , 
        \DataP/npc_pre[0] }), .LINK_ADD({\DataP/link_addr_F[31] , 
        \DataP/link_addr_F[30] , \DataP/link_addr_F[29] , 
        \DataP/link_addr_F[28] , \DataP/link_addr_F[27] , 
        \DataP/link_addr_F[26] , \DataP/link_addr_F[25] , 
        \DataP/link_addr_F[24] , \DataP/link_addr_F[23] , 
        \DataP/link_addr_F[22] , \DataP/link_addr_F[21] , 
        \DataP/link_addr_F[20] , \DataP/link_addr_F[19] , 
        \DataP/link_addr_F[18] , \DataP/link_addr_F[17] , 
        \DataP/link_addr_F[16] , \DataP/link_addr_F[15] , 
        \DataP/link_addr_F[14] , \DataP/link_addr_F[13] , 
        \DataP/link_addr_F[12] , \DataP/link_addr_F[11] , 
        \DataP/link_addr_F[10] , \DataP/link_addr_F[9] , 
        \DataP/link_addr_F[8] , \DataP/link_addr_F[7] , \DataP/link_addr_F[6] , 
        \DataP/link_addr_F[5] , \DataP/link_addr_F[4] , \DataP/link_addr_F[3] , 
        \DataP/link_addr_F[2] , \DataP/link_addr_F[1] , \DataP/link_addr_F[0] }), .SEL(\DataP/npc_mux_sel ), .TAKEN(\DataP/prediction ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[0]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N1 ), .Q(\DataP/npc[0] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[1]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N2 ), .Q(\DataP/npc[1] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[2]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N3 ), .Q(\DataP/npc[2] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[3]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N4 ), .Q(\DataP/npc[3] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[4]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N5 ), .Q(\DataP/npc[4] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[5]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N6 ), .Q(\DataP/npc[5] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[6]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N7 ), .Q(\DataP/npc[6] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[7]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N8 ), .Q(\DataP/npc[7] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[8]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N9 ), .Q(\DataP/npc[8] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[9]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N10 ), .Q(\DataP/npc[9] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[10]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N11 ), .Q(\DataP/npc[10] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[11]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N12 ), .Q(\DataP/npc[11] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[12]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N13 ), .Q(\DataP/npc[12] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[13]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N14 ), .Q(\DataP/npc[13] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[14]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N15 ), .Q(\DataP/npc[14] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[15]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N16 ), .Q(\DataP/npc[15] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[16]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N17 ), .Q(\DataP/npc[16] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[17]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N18 ), .Q(\DataP/npc[17] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[18]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N19 ), .Q(\DataP/npc[18] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[19]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N20 ), .Q(\DataP/npc[19] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[20]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N21 ), .Q(\DataP/npc[20] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[21]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N22 ), .Q(\DataP/npc[21] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[22]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N23 ), .Q(\DataP/npc[22] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[23]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N24 ), .Q(\DataP/npc[23] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[24]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N25 ), .Q(\DataP/npc[24] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[25]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N26 ), .Q(\DataP/npc[25] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[26]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N27 ), .Q(\DataP/npc[26] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[27]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N28 ), .Q(\DataP/npc[27] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[28]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N29 ), .Q(\DataP/npc[28] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[29]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N30 ), .Q(\DataP/npc[29] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[30]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N31 ), .Q(\DataP/npc[30] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[31]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N32 ), .Q(\DataP/npc[31] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[0]  ( .D(DRAM_DATA_OUT[0]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[0] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[1]  ( .D(DRAM_DATA_OUT[1]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[1] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[2]  ( .D(DRAM_DATA_OUT[2]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[2] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[3]  ( .D(DRAM_DATA_OUT[3]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[3] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[4]  ( .D(DRAM_DATA_OUT[4]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[4] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[5]  ( .D(DRAM_DATA_OUT[5]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[5] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[6]  ( .D(DRAM_DATA_OUT[6]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[6] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[7]  ( .D(DRAM_DATA_OUT[7]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[7] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[8]  ( .D(DRAM_DATA_OUT[8]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[8] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[9]  ( .D(DRAM_DATA_OUT[9]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[9] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[10]  ( .D(DRAM_DATA_OUT[10]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[10] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[11]  ( .D(DRAM_DATA_OUT[11]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[11] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[12]  ( .D(DRAM_DATA_OUT[12]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[12] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[13]  ( .D(DRAM_DATA_OUT[13]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[13] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[14]  ( .D(DRAM_DATA_OUT[14]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[14] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[15]  ( .D(DRAM_DATA_OUT[15]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[15] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[16]  ( .D(DRAM_DATA_OUT[16]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[16] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[17]  ( .D(DRAM_DATA_OUT[17]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[17] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[18]  ( .D(DRAM_DATA_OUT[18]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[18] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[19]  ( .D(DRAM_DATA_OUT[19]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[19] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[20]  ( .D(DRAM_DATA_OUT[20]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[20] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[21]  ( .D(DRAM_DATA_OUT[21]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[21] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[22]  ( .D(DRAM_DATA_OUT[22]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[22] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[23]  ( .D(DRAM_DATA_OUT[23]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[23] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[24]  ( .D(DRAM_DATA_OUT[24]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[24] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[25]  ( .D(DRAM_DATA_OUT[25]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[25] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[26]  ( .D(DRAM_DATA_OUT[26]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[26] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[27]  ( .D(DRAM_DATA_OUT[27]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[27] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[28]  ( .D(DRAM_DATA_OUT[28]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[28] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[29]  ( .D(DRAM_DATA_OUT[29]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[29] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[30]  ( .D(DRAM_DATA_OUT[30]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[30] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[31]  ( .D(DRAM_DATA_OUT[31]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[31] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[31]  ( .D(n297), .CK(Clk), .SN(Rst), .Q(
        n2414), .QN(\DataP/alu_out_M[31] ) );
  DFF_X1 \DataP/PC_reg/O_reg[31]  ( .D(\DataP/PC_reg/N33 ), .CK(Clk), .Q(
        \DataP/pc_out[31] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[31]  ( .D(n1481), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[31] ) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[31]  ( .D(n292), .CK(Clk), .SN(Rst), 
        .Q(n291) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[31]  ( .D(n291), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[31] ) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[0]  ( .D(\DataP/b_out[0] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[0] ), .QN(n290) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[0]  ( .D(n290), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[0]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[1]  ( .D(\DataP/b_out[1] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[1] ), .QN(n289) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[1]  ( .D(n289), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[1]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[2]  ( .D(\DataP/b_out[2] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[2] ), .QN(n288) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[2]  ( .D(n288), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[2]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[3]  ( .D(\DataP/b_out[3] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[3] ), .QN(n287) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[3]  ( .D(n287), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[3]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[4]  ( .D(\DataP/b_out[4] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[4] ), .QN(n286) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[4]  ( .D(n286), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[4]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[5]  ( .D(\DataP/b_out[5] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[5] ), .QN(n285) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[5]  ( .D(n285), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[5]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[6]  ( .D(\DataP/b_out[6] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[6] ), .QN(n284) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[6]  ( .D(n284), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[6]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[7]  ( .D(\DataP/b_out[7] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[7] ), .QN(n283) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[7]  ( .D(n283), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[7]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[8]  ( .D(\DataP/b_out[8] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[8] ), .QN(n282) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[8]  ( .D(n282), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[8]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[9]  ( .D(\DataP/b_out[9] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[9] ), .QN(n281) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[9]  ( .D(n281), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[9]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[10]  ( .D(\DataP/b_out[10] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[10] ), .QN(n280) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[10]  ( .D(n280), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[10]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[11]  ( .D(\DataP/b_out[11] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[11] ), .QN(n279) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[11]  ( .D(n279), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[11]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[12]  ( .D(\DataP/b_out[12] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[12] ), .QN(n278) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[12]  ( .D(n278), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[12]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[13]  ( .D(\DataP/b_out[13] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[13] ), .QN(n277) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[13]  ( .D(n277), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[13]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[14]  ( .D(\DataP/b_out[14] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[14] ), .QN(n276) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[14]  ( .D(n276), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[14]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[15]  ( .D(\DataP/b_out[15] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[15] ), .QN(n275) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[15]  ( .D(n275), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[15]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[16]  ( .D(\DataP/b_out[16] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[16] ), .QN(n274) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[16]  ( .D(n274), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[16]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[17]  ( .D(\DataP/b_out[17] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[17] ), .QN(n273) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[17]  ( .D(n273), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[17]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[18]  ( .D(\DataP/b_out[18] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[18] ), .QN(n272) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[18]  ( .D(n272), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[18]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[19]  ( .D(\DataP/b_out[19] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[19] ), .QN(n271) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[19]  ( .D(n271), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[19]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[20]  ( .D(\DataP/b_out[20] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[20] ), .QN(n270) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[20]  ( .D(n270), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[20]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[21]  ( .D(\DataP/b_out[21] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[21] ), .QN(n269) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[21]  ( .D(n269), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[21]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[22]  ( .D(\DataP/b_out[22] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[22] ), .QN(n268) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[22]  ( .D(n268), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[22]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[23]  ( .D(\DataP/b_out[23] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[23] ), .QN(n267) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[23]  ( .D(n267), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[23]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[24]  ( .D(\DataP/b_out[24] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[24] ), .QN(n266) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[24]  ( .D(n266), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[24]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[25]  ( .D(\DataP/b_out[25] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[25] ), .QN(n265) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[25]  ( .D(n265), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[25]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[26]  ( .D(\DataP/b_out[26] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[26] ), .QN(n264) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[26]  ( .D(n264), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[26]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[27]  ( .D(\DataP/b_out[27] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[27] ), .QN(n263) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[27]  ( .D(n263), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[27]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[28]  ( .D(\DataP/b_out[28] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[28] ), .QN(n262) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[28]  ( .D(n262), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[28]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[29]  ( .D(\DataP/b_out[29] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[29] ), .QN(n261) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[29]  ( .D(n261), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[29]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[30]  ( .D(\DataP/b_out[30] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[30] ), .QN(n260) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[30]  ( .D(n260), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[30]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[31]  ( .D(\DataP/b_out[31] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[31] ), .QN(n259) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[31]  ( .D(n259), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[31]) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[2]  ( .D(\DataP/a_out[2] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[2] ), .QN(n2459) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[8]  ( .D(\DataP/a_out[8] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[8] ), .QN(n2467) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[9]  ( .D(\DataP/a_out[9] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[9] ), .QN(n2435) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[15]  ( .D(n330), .CK(Clk), .SN(Rst), .Q(
        n2433), .QN(\DataP/alu_out_M[15] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[19]  ( .D(n319), .CK(Clk), .SN(Rst), .Q(
        n2421), .QN(\DataP/alu_out_M[19] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[30]  ( .D(n2774), .CK(Clk), .SN(Rst), 
        .Q(n2417), .QN(\DataP/alu_out_M[30] ) );
  DFFR_X1 \DataP/IF_IDs/PR_OUT_reg  ( .D(n1449), .CK(Clk), .RN(Rst), .Q(
        \DataP/pr_D ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[30]  ( .D(n1450), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[30] ), .QN(n257) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[30]  ( .D(n257), .CK(Clk), .SN(Rst), .Q(
        n256) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[30]  ( .D(n256), .CK(Clk), .SN(Rst), 
        .Q(n255) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[30]  ( .D(n255), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[30] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[29]  ( .D(n1451), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[29] ), .QN(n254) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[29]  ( .D(n254), .CK(Clk), .SN(Rst), .Q(
        n253) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[29]  ( .D(n253), .CK(Clk), .SN(Rst), 
        .Q(n252) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[29]  ( .D(n252), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[29] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[28]  ( .D(n1452), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[28] ), .QN(n251) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[28]  ( .D(n251), .CK(Clk), .SN(Rst), .Q(
        n250) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[28]  ( .D(n250), .CK(Clk), .SN(Rst), 
        .Q(n249) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[28]  ( .D(n249), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[28] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[27]  ( .D(n1453), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[27] ), .QN(n248) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[27]  ( .D(n248), .CK(Clk), .SN(Rst), .Q(
        n247) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[27]  ( .D(n247), .CK(Clk), .SN(Rst), 
        .Q(n246) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[27]  ( .D(n246), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[27] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[26]  ( .D(n1454), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[26] ), .QN(n245) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[26]  ( .D(n245), .CK(Clk), .SN(Rst), .Q(
        n244) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[26]  ( .D(n244), .CK(Clk), .SN(Rst), 
        .Q(n243) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[26]  ( .D(n243), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[26] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[25]  ( .D(n1455), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[25] ), .QN(n242) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[25]  ( .D(n242), .CK(Clk), .SN(Rst), .Q(
        n241) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[25]  ( .D(n241), .CK(Clk), .SN(Rst), 
        .Q(n240) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[25]  ( .D(n240), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[25] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[24]  ( .D(n1456), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[24] ), .QN(n239) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[24]  ( .D(n239), .CK(Clk), .SN(Rst), .Q(
        n238) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[24]  ( .D(n238), .CK(Clk), .SN(Rst), 
        .Q(n237) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[24]  ( .D(n237), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[24] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[23]  ( .D(n1457), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[23] ), .QN(n236) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[23]  ( .D(n236), .CK(Clk), .SN(Rst), .Q(
        n235) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[23]  ( .D(n235), .CK(Clk), .SN(Rst), 
        .Q(n234) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[23]  ( .D(n234), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[23] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[22]  ( .D(n1458), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[22] ), .QN(n233) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[22]  ( .D(n233), .CK(Clk), .SN(Rst), .Q(
        n232) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[22]  ( .D(n232), .CK(Clk), .SN(Rst), 
        .Q(n231) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[22]  ( .D(n231), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[22] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[21]  ( .D(n1459), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[21] ), .QN(n230) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[21]  ( .D(n230), .CK(Clk), .SN(Rst), .Q(
        n229) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[21]  ( .D(n229), .CK(Clk), .SN(Rst), 
        .Q(n228) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[21]  ( .D(n228), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[21] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[20]  ( .D(n1460), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[20] ), .QN(n227) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[20]  ( .D(n227), .CK(Clk), .SN(Rst), .Q(
        n226) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[20]  ( .D(n226), .CK(Clk), .SN(Rst), 
        .Q(n225) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[20]  ( .D(n225), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[20] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[19]  ( .D(n1461), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[19] ), .QN(n224) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[19]  ( .D(n224), .CK(Clk), .SN(Rst), .Q(
        n223) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[19]  ( .D(n223), .CK(Clk), .SN(Rst), 
        .Q(n222) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[19]  ( .D(n222), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[19] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[18]  ( .D(n1462), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[18] ), .QN(n221) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[18]  ( .D(n221), .CK(Clk), .SN(Rst), .Q(
        n220) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[18]  ( .D(n220), .CK(Clk), .SN(Rst), 
        .Q(n219) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[18]  ( .D(n219), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[18] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[17]  ( .D(n1463), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[17] ), .QN(n218) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[17]  ( .D(n218), .CK(Clk), .SN(Rst), .Q(
        n217) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[17]  ( .D(n217), .CK(Clk), .SN(Rst), 
        .Q(n216) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[17]  ( .D(n216), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[17] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[16]  ( .D(n1464), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[16] ), .QN(n215) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[16]  ( .D(n215), .CK(Clk), .SN(Rst), .Q(
        n214) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[16]  ( .D(n214), .CK(Clk), .SN(Rst), 
        .Q(n213) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[16]  ( .D(n213), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[16] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[15]  ( .D(n1465), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[15] ), .QN(n212) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[15]  ( .D(n212), .CK(Clk), .SN(Rst), .Q(
        n211) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[15]  ( .D(n211), .CK(Clk), .SN(Rst), 
        .Q(n210) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[15]  ( .D(n210), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[15] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[14]  ( .D(n1466), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[14] ), .QN(n209) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[14]  ( .D(n209), .CK(Clk), .SN(Rst), .Q(
        n208) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[14]  ( .D(n208), .CK(Clk), .SN(Rst), 
        .Q(n207) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[14]  ( .D(n207), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[14] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[13]  ( .D(n1467), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[13] ), .QN(n206) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[13]  ( .D(n206), .CK(Clk), .SN(Rst), .Q(
        n205) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[13]  ( .D(n205), .CK(Clk), .SN(Rst), 
        .Q(n204) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[13]  ( .D(n204), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[13] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[12]  ( .D(n1468), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[12] ), .QN(n203) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[12]  ( .D(n203), .CK(Clk), .SN(Rst), .Q(
        n202) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[12]  ( .D(n202), .CK(Clk), .SN(Rst), 
        .Q(n201) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[12]  ( .D(n201), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[12] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[11]  ( .D(n1469), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[11] ), .QN(n200) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[11]  ( .D(n200), .CK(Clk), .SN(Rst), .Q(
        n199) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[11]  ( .D(n199), .CK(Clk), .SN(Rst), 
        .Q(n198) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[11]  ( .D(n198), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[11] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[10]  ( .D(n1470), .CK(Clk), .RN(Rst), 
        .Q(\DataP/link_addr_D[10] ), .QN(n197) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[10]  ( .D(n197), .CK(Clk), .SN(Rst), .Q(
        n196) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[10]  ( .D(n196), .CK(Clk), .SN(Rst), 
        .Q(n195) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[10]  ( .D(n195), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[10] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[9]  ( .D(n1471), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[9] ), .QN(n194) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[9]  ( .D(n194), .CK(Clk), .SN(Rst), .Q(
        n193) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[9]  ( .D(n193), .CK(Clk), .SN(Rst), 
        .Q(n192) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[9]  ( .D(n192), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[9] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[8]  ( .D(n1472), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[8] ), .QN(n191) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[8]  ( .D(n191), .CK(Clk), .SN(Rst), .Q(
        n190) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[8]  ( .D(n190), .CK(Clk), .SN(Rst), 
        .Q(n189) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[8]  ( .D(n189), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[8] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[7]  ( .D(n1473), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[7] ), .QN(n188) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[7]  ( .D(n188), .CK(Clk), .SN(Rst), .Q(
        n187) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[7]  ( .D(n187), .CK(Clk), .SN(Rst), 
        .Q(n186) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[7]  ( .D(n186), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[7] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[6]  ( .D(n1474), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[6] ), .QN(n185) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[6]  ( .D(n185), .CK(Clk), .SN(Rst), .Q(
        n184) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[6]  ( .D(n184), .CK(Clk), .SN(Rst), 
        .Q(n183) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[6]  ( .D(n183), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[6] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[5]  ( .D(n1475), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[5] ), .QN(n182) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[5]  ( .D(n182), .CK(Clk), .SN(Rst), .Q(
        n181) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[5]  ( .D(n181), .CK(Clk), .SN(Rst), 
        .Q(n180) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[5]  ( .D(n180), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[5] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[4]  ( .D(n1476), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[4] ), .QN(n179) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[4]  ( .D(n179), .CK(Clk), .SN(Rst), .Q(
        n178) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[4]  ( .D(n178), .CK(Clk), .SN(Rst), 
        .Q(n177) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[4]  ( .D(n177), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[4] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[3]  ( .D(n1477), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[3] ), .QN(n176) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[3]  ( .D(n176), .CK(Clk), .SN(Rst), .Q(
        n175) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[3]  ( .D(n175), .CK(Clk), .SN(Rst), 
        .Q(n174) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[3]  ( .D(n174), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[3] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[2]  ( .D(n1478), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[2] ), .QN(n173) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[2]  ( .D(n173), .CK(Clk), .SN(Rst), .Q(
        n172) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[2]  ( .D(n172), .CK(Clk), .SN(Rst), 
        .Q(n171) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[2]  ( .D(n171), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[2] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[1]  ( .D(n1479), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[1] ), .QN(n170) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[1]  ( .D(n170), .CK(Clk), .SN(Rst), .Q(
        n169) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[1]  ( .D(n169), .CK(Clk), .SN(Rst), 
        .Q(n168) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[1]  ( .D(n168), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[1] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[0]  ( .D(n1480), .CK(Clk), .RN(Rst), .Q(
        \DataP/link_addr_D[0] ), .QN(n167) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[0]  ( .D(n167), .CK(Clk), .SN(Rst), .Q(
        n166) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[0]  ( .D(n166), .CK(Clk), .SN(Rst), 
        .Q(n165) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[0]  ( .D(n165), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[0] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[31]  ( .D(\DataP/npc[31] ), .CK(Clk), 
        .RN(n162), .SN(n163), .QN(n164) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[31]  ( .D(n164), .CK(Clk), .SN(Rst), .Q(
        n161) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[31]  ( .D(n161), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[31] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[30]  ( .D(\DataP/npc[30] ), .CK(Clk), 
        .RN(n158), .SN(n159), .QN(n160) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[30]  ( .D(n160), .CK(Clk), .SN(Rst), .Q(
        n157) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[30]  ( .D(n157), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[30] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[29]  ( .D(\DataP/npc[29] ), .CK(Clk), 
        .RN(n154), .SN(n155), .QN(n156) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[29]  ( .D(n156), .CK(Clk), .SN(Rst), .Q(
        n153) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[29]  ( .D(n153), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[29] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[28]  ( .D(\DataP/npc[28] ), .CK(Clk), 
        .RN(n150), .SN(n151), .QN(n152) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[28]  ( .D(n152), .CK(Clk), .SN(Rst), .Q(
        n149) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[28]  ( .D(n149), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[28] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[27]  ( .D(\DataP/npc[27] ), .CK(Clk), 
        .RN(n146), .SN(n147), .QN(n148) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[27]  ( .D(n148), .CK(Clk), .SN(Rst), .Q(
        n145) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[27]  ( .D(n145), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[27] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[26]  ( .D(\DataP/npc[26] ), .CK(Clk), 
        .RN(n142), .SN(n143), .QN(n144) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[26]  ( .D(n144), .CK(Clk), .SN(Rst), .Q(
        n141) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[26]  ( .D(n141), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[26] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[25]  ( .D(\DataP/npc[25] ), .CK(Clk), 
        .RN(n138), .SN(n139), .QN(n140) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[25]  ( .D(n140), .CK(Clk), .SN(Rst), .Q(
        n137) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[25]  ( .D(n137), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[25] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[24]  ( .D(\DataP/npc[24] ), .CK(Clk), 
        .RN(n134), .SN(n135), .QN(n136) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[24]  ( .D(n136), .CK(Clk), .SN(Rst), .Q(
        n133) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[24]  ( .D(n133), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[24] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[23]  ( .D(\DataP/npc[23] ), .CK(Clk), 
        .RN(n130), .SN(n131), .QN(n132) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[23]  ( .D(n132), .CK(Clk), .SN(Rst), .Q(
        n129) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[23]  ( .D(n129), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[23] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[22]  ( .D(\DataP/npc[22] ), .CK(Clk), 
        .RN(n126), .SN(n127), .QN(n128) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[22]  ( .D(n128), .CK(Clk), .SN(Rst), .Q(
        n125) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[22]  ( .D(n125), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[22] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[21]  ( .D(\DataP/npc[21] ), .CK(Clk), 
        .RN(n122), .SN(n123), .QN(n124) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[21]  ( .D(n124), .CK(Clk), .SN(Rst), .Q(
        n121) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[21]  ( .D(n121), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[21] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[20]  ( .D(\DataP/npc[20] ), .CK(Clk), 
        .RN(n118), .SN(n119), .QN(n120) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[20]  ( .D(n120), .CK(Clk), .SN(Rst), .Q(
        n117) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[20]  ( .D(n117), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[20] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[19]  ( .D(\DataP/npc[19] ), .CK(Clk), 
        .RN(n114), .SN(n115), .QN(n116) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[19]  ( .D(n116), .CK(Clk), .SN(Rst), .Q(
        n113) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[19]  ( .D(n113), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[19] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[18]  ( .D(\DataP/npc[18] ), .CK(Clk), 
        .RN(n110), .SN(n111), .QN(n112) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[18]  ( .D(n112), .CK(Clk), .SN(Rst), .Q(
        n109) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[18]  ( .D(n109), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[18] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[17]  ( .D(\DataP/npc[17] ), .CK(Clk), 
        .RN(n106), .SN(n107), .QN(n108) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[17]  ( .D(n108), .CK(Clk), .SN(Rst), .Q(
        n105), .QN(n1606) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[17]  ( .D(n105), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[17] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[16]  ( .D(\DataP/npc[16] ), .CK(Clk), 
        .RN(n102), .SN(n103), .QN(n104) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[16]  ( .D(n104), .CK(Clk), .SN(Rst), .Q(
        n101) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[16]  ( .D(n101), .CK(Clk), .SN(Rst), 
        .QN(\DataP/npc_M[16] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[15]  ( .D(\DataP/npc[15] ), .CK(Clk), 
        .RN(n98), .SN(n99), .QN(n100) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[15]  ( .D(n100), .CK(Clk), .SN(Rst), .Q(
        n97) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[15]  ( .D(n97), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[15] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[14]  ( .D(\DataP/npc[14] ), .CK(Clk), 
        .RN(n94), .SN(n95), .QN(n96) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[14]  ( .D(n96), .CK(Clk), .SN(Rst), .Q(n93) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[14]  ( .D(n93), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[14] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[13]  ( .D(\DataP/npc[13] ), .CK(Clk), 
        .RN(n90), .SN(n91), .QN(n92) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[13]  ( .D(n92), .CK(Clk), .SN(Rst), .Q(n89) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[13]  ( .D(n89), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[13] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[12]  ( .D(\DataP/npc[12] ), .CK(Clk), 
        .RN(n86), .SN(n87), .QN(n88) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[12]  ( .D(n88), .CK(Clk), .SN(Rst), .Q(n85), .QN(n1969) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[12]  ( .D(n85), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[12] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[11]  ( .D(\DataP/npc[11] ), .CK(Clk), 
        .RN(n82), .SN(n83), .QN(n84) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[11]  ( .D(n84), .CK(Clk), .SN(Rst), .Q(n81) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[11]  ( .D(n81), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[11] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[10]  ( .D(\DataP/npc[10] ), .CK(Clk), 
        .RN(n78), .SN(n79), .QN(n80) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[10]  ( .D(n80), .CK(Clk), .SN(Rst), .Q(n77) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[10]  ( .D(n77), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[10] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[9]  ( .D(\DataP/npc[9] ), .CK(Clk), .RN(
        n74), .SN(n75), .QN(n76) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[9]  ( .D(n76), .CK(Clk), .SN(Rst), .Q(n73), 
        .QN(\DataP/npc_E[9] ) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[9]  ( .D(n73), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[9] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[8]  ( .D(\DataP/npc[8] ), .CK(Clk), .RN(
        n70), .SN(n71), .QN(n72) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[8]  ( .D(n72), .CK(Clk), .SN(Rst), .Q(n69)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[8]  ( .D(n69), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[8] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[7]  ( .D(\DataP/npc[7] ), .CK(Clk), .RN(
        n66), .SN(n67), .QN(n68) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[7]  ( .D(n68), .CK(Clk), .SN(Rst), .Q(n65)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[7]  ( .D(n65), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[7] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[6]  ( .D(\DataP/npc[6] ), .CK(Clk), .RN(
        n62), .SN(n63), .QN(n64) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[6]  ( .D(n64), .CK(Clk), .SN(Rst), .Q(n61)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[6]  ( .D(n61), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[6] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[5]  ( .D(\DataP/npc[5] ), .CK(Clk), .RN(
        n58), .SN(n59), .QN(n60) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[5]  ( .D(n60), .CK(Clk), .SN(Rst), .Q(n57)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[5]  ( .D(n57), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[5] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[4]  ( .D(\DataP/npc[4] ), .CK(Clk), .RN(
        n54), .SN(n55), .QN(n56) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[4]  ( .D(n56), .CK(Clk), .SN(Rst), .Q(n53)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[4]  ( .D(n53), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[4] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[3]  ( .D(\DataP/npc[3] ), .CK(Clk), .RN(
        n50), .SN(n51), .QN(n52) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[3]  ( .D(n52), .CK(Clk), .SN(Rst), .Q(n49)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[3]  ( .D(n49), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[3] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[2]  ( .D(\DataP/npc[2] ), .CK(Clk), .RN(
        n46), .SN(n47), .QN(n48) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[2]  ( .D(n48), .CK(Clk), .SN(Rst), .Q(n45)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[2]  ( .D(n45), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[2] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[1]  ( .D(\DataP/npc[1] ), .CK(Clk), .RN(
        n42), .SN(n43), .QN(n44) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[1]  ( .D(n44), .CK(Clk), .SN(Rst), .Q(n41)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[1]  ( .D(n41), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[1] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[0]  ( .D(\DataP/npc[0] ), .CK(Clk), .RN(
        n38), .SN(n39), .QN(n40) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[0]  ( .D(n40), .CK(Clk), .SN(Rst), .Q(n37)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[0]  ( .D(n37), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[0] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[0]  ( .D(IRAM_DATA_OUT[0]), .CK(Clk), .RN(
        n36), .Q(IR_CU[0]), .QN(n476) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[0]  ( .D(n476), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[0] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[1]  ( .D(IRAM_DATA_OUT[1]), .CK(Clk), .RN(
        n36), .Q(IR_CU[1]), .QN(n477) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[1]  ( .D(n477), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[1] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[2]  ( .D(IRAM_DATA_OUT[2]), .CK(Clk), .RN(
        n36), .Q(n2375), .QN(n478) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[2]  ( .D(n478), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[2] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[3]  ( .D(IRAM_DATA_OUT[3]), .CK(Clk), .RN(
        n36), .Q(n2399), .QN(n479) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[3]  ( .D(n479), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[3] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[4]  ( .D(IRAM_DATA_OUT[4]), .CK(Clk), .RN(
        n36), .Q(IR_CU[4]), .QN(n480) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[4]  ( .D(n480), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[4] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[5]  ( .D(IRAM_DATA_OUT[5]), .CK(Clk), .RN(
        n36), .Q(IR_CU[5]), .QN(n482) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[5]  ( .D(n482), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[5] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[6]  ( .D(IRAM_DATA_OUT[6]), .CK(Clk), .RN(
        n36), .Q(IR_CU[6]), .QN(n35) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[6]  ( .D(n35), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[6] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[7]  ( .D(IRAM_DATA_OUT[7]), .CK(Clk), .RN(
        n36), .Q(IR_CU[7]), .QN(n34) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[7]  ( .D(n34), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[7] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[8]  ( .D(IRAM_DATA_OUT[8]), .CK(Clk), .RN(
        n36), .Q(IR_CU[8]), .QN(n33) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[8]  ( .D(n33), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[8] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[9]  ( .D(IRAM_DATA_OUT[9]), .CK(Clk), .RN(
        n36), .Q(IR_CU[9]), .QN(n32) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[9]  ( .D(n32), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[9] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[10]  ( .D(IRAM_DATA_OUT[10]), .CK(Clk), 
        .RN(n36), .QN(n484) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[10]  ( .D(n484), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[10] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[11]  ( .D(IRAM_DATA_OUT[11]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[11] ), .QN(n31) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[11]  ( .D(n31), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[11] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[12]  ( .D(IRAM_DATA_OUT[12]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[12] ), .QN(n30) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[12]  ( .D(n30), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[12] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[13]  ( .D(IRAM_DATA_OUT[13]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[13] ), .QN(n29) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[13]  ( .D(n29), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[13] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[14]  ( .D(IRAM_DATA_OUT[14]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[14] ), .QN(n28) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[14]  ( .D(n28), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[14] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[15]  ( .D(IRAM_DATA_OUT[15]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[15] ), .QN(n27) );
  DFFS_X1 \DataP/ID_EXs/IMM_OUT_reg[15]  ( .D(n27), .CK(Clk), .SN(Rst), .QN(
        \DataP/IMM_s[15] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[16]  ( .D(IRAM_DATA_OUT[16]), .CK(Clk), 
        .RN(n36), .QN(n485) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[17]  ( .D(IRAM_DATA_OUT[17]), .CK(Clk), 
        .RN(n36), .QN(n486) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[18]  ( .D(IRAM_DATA_OUT[18]), .CK(Clk), 
        .RN(n36), .QN(n487) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[19]  ( .D(IRAM_DATA_OUT[19]), .CK(Clk), 
        .RN(n36), .QN(n488) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[20]  ( .D(IRAM_DATA_OUT[20]), .CK(Clk), 
        .RN(n36), .QN(n489) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[21]  ( .D(IRAM_DATA_OUT[21]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[21] ), .QN(n26) );
  DFFS_X1 \DataP/ID_EXs/RS1_OUT_reg[0]  ( .D(n26), .CK(Clk), .SN(Rst), .Q(
        n2392) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[22]  ( .D(IRAM_DATA_OUT[22]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[22] ), .QN(n25) );
  DFFS_X1 \DataP/ID_EXs/RS1_OUT_reg[1]  ( .D(n25), .CK(Clk), .SN(Rst), .Q(
        n2429), .QN(\DataP/Rs1[1] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[23]  ( .D(IRAM_DATA_OUT[23]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[23] ), .QN(n24) );
  DFFS_X1 \DataP/ID_EXs/RS1_OUT_reg[2]  ( .D(n24), .CK(Clk), .SN(Rst), .Q(
        n2407), .QN(\DataP/Rs1[2] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[24]  ( .D(IRAM_DATA_OUT[24]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[24] ) );
  DFFR_X1 \DataP/ID_EXs/RS1_OUT_reg[3]  ( .D(\DataP/IR1[24] ), .CK(Clk), .RN(
        Rst), .QN(n523) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[25]  ( .D(IRAM_DATA_OUT[25]), .CK(Clk), 
        .RN(n36), .Q(\DataP/IR1[25] ) );
  DFFR_X1 \DataP/ID_EXs/RS1_OUT_reg[4]  ( .D(\DataP/IR1[25] ), .CK(Clk), .RN(
        Rst), .QN(n524) );
  DFFS_X1 \DataP/IF_IDs/IR_OUT_reg[26]  ( .D(IRAM_DATA_OUT[26]), .CK(Clk), 
        .SN(n36), .Q(IR_CU_26), .QN(n497) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[0]  ( .D(n497), .CK(Clk), .SN(Rst), .Q(
        n23), .QN(\DataP/opcode_E[0] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[0]  ( .D(n23), .CK(Clk), .SN(Rst), 
        .Q(n22), .QN(\DataP/opcode_M[0] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[0]  ( .D(n22), .CK(Clk), .SN(Rst), 
        .Q(n2403), .QN(\DataP/opcode_W[0] ) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[1]  ( .D(n504), .CK(Clk), .SN(Rst), .Q(
        n520), .QN(\DataP/opcode_E[1] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[1]  ( .D(n520), .CK(Clk), .SN(Rst), 
        .Q(n2249), .QN(\DataP/opcode_M[1] ) );
  DFFS_X1 \DataP/IF_IDs/IR_OUT_reg[28]  ( .D(IRAM_DATA_OUT[28]), .CK(Clk), 
        .SN(n36), .Q(IR_CU_28), .QN(n1960) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[29]  ( .D(IRAM_DATA_OUT[29]), .CK(Clk), 
        .RN(n36), .Q(n2374), .QN(n514) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[3]  ( .D(n514), .CK(Clk), .SN(Rst), .Q(
        n21), .QN(\DataP/opcode_E[3] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[3]  ( .D(n21), .CK(Clk), .SN(Rst), 
        .Q(n20), .QN(\DataP/opcode_M[3] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[3]  ( .D(n20), .CK(Clk), .SN(Rst), 
        .Q(n2401), .QN(\DataP/opcode_W[3] ) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[4]  ( .D(n515), .CK(Clk), .SN(Rst), .Q(
        n19), .QN(\DataP/opcode_E[4] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[4]  ( .D(n19), .CK(Clk), .SN(Rst), 
        .Q(n18), .QN(\DataP/opcode_M[4] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[4]  ( .D(n18), .CK(Clk), .SN(Rst), 
        .Q(n2383), .QN(\DataP/opcode_W[4] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[31]  ( .D(IRAM_DATA_OUT[31]), .CK(Clk), 
        .RN(n36), .Q(IR_CU_31), .QN(n516) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[5]  ( .D(n17), .CK(Clk), .SN(Rst), 
        .Q(n2387) );
  DLH_X1 \DataP/FORWARDING_BR/SEL_reg[1]  ( .G(\DataP/FORWARDING_BR/N12 ), .D(
        n3910), .Q(\DataP/FWD_MUX_BR_S[1] ) );
  SDFFR_X1 \CU_I/cw1_reg[8]  ( .D(n16), .SI(n607), .SE(n504), .CK(Clk), .RN(
        Rst), .Q(BR_EN_i) );
  DFFR_X1 \CU_I/cw1_reg[7]  ( .D(\CU_I/cw[7] ), .CK(Clk), .RN(Rst), .QN(n15)
         );
  DFFS_X1 \CU_I/cw2_reg[7]  ( .D(n15), .CK(Clk), .SN(Rst), .QN(DRAM_RW) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[4]  ( .D(\DataP/dest_D[4] ), .CK(Clk), .RN(
        Rst), .QN(n14) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[3]  ( .D(\DataP/dest_D[3] ), .CK(Clk), .RN(
        Rst), .QN(n13) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[2]  ( .D(\DataP/dest_D[2] ), .CK(Clk), .RN(
        Rst), .QN(n12) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[2]  ( .D(n12), .CK(Clk), .SN(Rst), .Q(
        n530), .QN(\DataP/dest_M[2] ) );
  DFFR_X1 \DataP/MEM_WB_s/RD_OUT_reg[2]  ( .D(\DataP/dest_M[2] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/add_D[2] ), .QN(n538) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[1]  ( .D(\DataP/dest_D[1] ), .CK(Clk), .RN(
        Rst), .QN(n11) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[0]  ( .D(\DataP/dest_D[0] ), .CK(Clk), .RN(
        Rst), .QN(n10) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[0]  ( .D(n10), .CK(Clk), .SN(Rst), .Q(
        n528), .QN(\DataP/dest_M[0] ) );
  DFFR_X1 \DataP/MEM_WB_s/RD_OUT_reg[0]  ( .D(\DataP/dest_M[0] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/add_D[0] ), .QN(n536) );
  DLH_X1 \DataP/FORWARDING_BR/SEL_reg[0]  ( .G(\DataP/FORWARDING_BR/N12 ), .D(
        n3909), .Q(\DataP/FWD_MUX_BR_S[0] ) );
  DFFR_X1 \CU_I/aluOpcode1_reg[2]  ( .D(\CU_I/aluOpcode_i[2] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[2]), .QN(n2391) );
  DFFS_X1 \CU_I/cw1_reg[5]  ( .D(n1358), .CK(Clk), .SN(Rst), .Q(n9) );
  DFFS_X1 \CU_I/cw2_reg[5]  ( .D(n9), .CK(Clk), .SN(Rst), .QN(DRAM_SEL[2]) );
  DFFR_X1 \CU_I/cw1_reg[0]  ( .D(\CU_I/cw[0] ), .CK(Clk), .RN(Rst), .QN(n8) );
  DFFS_X1 \CU_I/cw2_reg[0]  ( .D(n8), .CK(Clk), .SN(Rst), .Q(n7) );
  DFFS_X1 \CU_I/cw3_reg[0]  ( .D(n7), .CK(Clk), .SN(Rst), .QN(RF_WE_i) );
  DFFS_X1 \CU_I/cw1_reg[2]  ( .D(n1372), .CK(Clk), .SN(Rst), .Q(n6) );
  DFFS_X1 \CU_I/cw2_reg[2]  ( .D(n6), .CK(Clk), .SN(Rst), .Q(n5) );
  DFFS_X1 \CU_I/cw3_reg[2]  ( .D(n5), .CK(Clk), .SN(Rst), .QN(
        \WB_MUX_SEL_i[1] ) );
  DFFR_X1 \CU_I/cw1_reg[4]  ( .D(\CU_I/cw[4] ), .CK(Clk), .RN(Rst), .QN(n4) );
  DFFS_X1 \CU_I/cw2_reg[4]  ( .D(n4), .CK(Clk), .SN(Rst), .QN(DRAM_SEL[1]) );
  DFFR_X1 \CU_I/cw1_reg[3]  ( .D(\CU_I/cw[3] ), .CK(Clk), .RN(Rst), .QN(n3) );
  DFFS_X1 \CU_I/cw2_reg[3]  ( .D(n3), .CK(Clk), .SN(Rst), .QN(DRAM_SEL[0]) );
  DFFR_X1 \CU_I/cw1_reg[6]  ( .D(\CU_I/cw[6] ), .CK(Clk), .RN(Rst), .QN(n2) );
  DFFS_X1 \CU_I/cw2_reg[6]  ( .D(n2), .CK(Clk), .SN(Rst), .QN(DRAM_ENABLE) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[12]  ( .D(n337), .CK(Clk), .SN(Rst), .Q(
        n2424), .QN(\DataP/alu_out_M[12] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[13]  ( .D(n333), .CK(Clk), .SN(Rst), .Q(
        n2423), .QN(\DataP/alu_out_M[13] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[14]  ( .D(n332), .CK(Clk), .SN(Rst), .Q(
        n2418), .QN(\DataP/alu_out_M[14] ) );
  DFF_X1 \DataP/PC_reg/O_reg[14]  ( .D(\DataP/PC_reg/N16 ), .CK(Clk), .Q(
        \DataP/pc_out[14] ) );
  DFF_X1 \DataP/PC_reg/O_reg[13]  ( .D(\DataP/PC_reg/N15 ), .CK(Clk), .Q(
        \DataP/pc_out[13] ) );
  DFF_X1 \DataP/PC_reg/O_reg[12]  ( .D(\DataP/PC_reg/N14 ), .CK(Clk), .Q(
        \DataP/pc_out[12] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[4]  ( .D(n355), .CK(Clk), .SN(Rst), .Q(
        n2466), .QN(DRAM_ADDRESS[4]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[5]  ( .D(n354), .CK(Clk), .SN(Rst), .Q(
        n2450), .QN(DRAM_ADDRESS[5]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[6]  ( .D(n353), .CK(Clk), .SN(Rst), .Q(
        n2410), .QN(DRAM_ADDRESS[6]) );
  DFF_X1 \DataP/PC_reg/O_reg[6]  ( .D(\DataP/PC_reg/N8 ), .CK(Clk), .Q(
        IRAM_ADDRESS[4]) );
  DFF_X1 \DataP/PC_reg/O_reg[5]  ( .D(\DataP/PC_reg/N7 ), .CK(Clk), .Q(
        IRAM_ADDRESS[3]) );
  DFF_X1 \DataP/PC_reg/O_reg[4]  ( .D(\DataP/PC_reg/N6 ), .CK(Clk), .Q(
        IRAM_ADDRESS[2]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[1]  ( .D(n358), .CK(Clk), .SN(Rst), .Q(
        n2469), .QN(DRAM_ADDRESS[1]) );
  DFF_X1 \DataP/PC_reg/O_reg[1]  ( .D(\DataP/PC_reg/N3 ), .CK(Clk), .Q(
        \DataP/pc_out_1 ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[2]  ( .D(n357), .CK(Clk), .SN(Rst), .Q(
        n2471), .QN(DRAM_ADDRESS[2]) );
  DFF_X1 \DataP/PC_reg/O_reg[2]  ( .D(\DataP/PC_reg/N4 ), .CK(Clk), .Q(
        IRAM_ADDRESS[0]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[3]  ( .D(n356), .CK(Clk), .SN(Rst), .Q(
        n2478), .QN(DRAM_ADDRESS[3]) );
  DFF_X1 \DataP/PC_reg/O_reg[3]  ( .D(\DataP/PC_reg/N5 ), .CK(Clk), .Q(
        IRAM_ADDRESS[1]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[8]  ( .D(n345), .CK(Clk), .SN(Rst), .Q(
        n2408), .QN(DRAM_ADDRESS[8]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[9]  ( .D(n341), .CK(Clk), .SN(Rst), .Q(
        n2477), .QN(DRAM_ADDRESS[9]) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[10]  ( .D(n340), .CK(Clk), .SN(Rst), .Q(
        n2409), .QN(DRAM_ADDRESS[10]) );
  DFF_X1 \DataP/PC_reg/O_reg[10]  ( .D(\DataP/PC_reg/N12 ), .CK(Clk), .Q(
        \DataP/pc_out[10] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[11]  ( .D(n2386), .CK(Clk), .SN(Rst), 
        .Q(n2431), .QN(DRAM_ADDRESS[11]) );
  DFF_X1 \DataP/PC_reg/O_reg[9]  ( .D(\DataP/PC_reg/N11 ), .CK(Clk), .Q(
        IRAM_ADDRESS[7]) );
  DFF_X1 \DataP/PC_reg/O_reg[8]  ( .D(\DataP/PC_reg/N10 ), .CK(Clk), .Q(
        IRAM_ADDRESS[6]) );
  DFFR_X1 \CU_I/cw1_reg[1]  ( .D(\CU_I/cw[1] ), .CK(Clk), .RN(Rst), .QN(n1) );
  DFFS_X1 \CU_I/cw2_reg[1]  ( .D(n1), .CK(Clk), .SN(Rst), .QN(\CU_I/cw2[1] )
         );
  DFFR_X1 \CU_I/cw3_reg[1]  ( .D(\CU_I/cw2[1] ), .CK(Clk), .RN(Rst), .QN(n294)
         );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[28]  ( .D(n300), .CK(Clk), .SN(Rst), .Q(
        n2426), .QN(\DataP/alu_out_M[28] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[24]  ( .D(n1759), .CK(Clk), .SN(Rst), 
        .Q(n2427), .QN(\DataP/alu_out_M[24] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[25]  ( .D(n1624), .CK(Clk), .SN(Rst), 
        .Q(n2422), .QN(\DataP/alu_out_M[25] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[20]  ( .D(n317), .CK(Clk), .SN(Rst), .Q(
        n2420), .QN(\DataP/alu_out_M[20] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[21]  ( .D(n313), .CK(Clk), .SN(Rst), .Q(
        n2419), .QN(\DataP/alu_out_M[21] ) );
  DFF_X1 \DataP/PC_reg/O_reg[22]  ( .D(\DataP/PC_reg/N24 ), .CK(Clk), .Q(
        \DataP/pc_out[22] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[16]  ( .D(n326), .CK(Clk), .SN(Rst), .Q(
        n2412), .QN(\DataP/alu_out_M[16] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[18]  ( .D(n322), .CK(Clk), .SN(Rst), .Q(
        n2425), .QN(\DataP/alu_out_M[18] ) );
  DFF_X1 \DataP/PC_reg/O_reg[18]  ( .D(\DataP/PC_reg/N20 ), .CK(Clk), .Q(
        \DataP/pc_out[18] ) );
  DFF_X1 \DataP/PC_reg/O_reg[16]  ( .D(\DataP/PC_reg/N18 ), .CK(Clk), .Q(
        \DataP/pc_out[16] ) );
  DFF_X1 \DataP/PC_reg/O_reg[27]  ( .D(\DataP/PC_reg/N29 ), .CK(Clk), .Q(
        \DataP/pc_out[27] ) );
  DFF_X1 \DataP/PC_reg/O_reg[23]  ( .D(\DataP/PC_reg/N25 ), .CK(Clk), .Q(
        \DataP/pc_out[23] ) );
  DFF_X1 \DataP/PC_reg/O_reg[19]  ( .D(\DataP/PC_reg/N21 ), .CK(Clk), .Q(
        \DataP/pc_out[19] ) );
  DFF_X1 \DataP/PC_reg/O_reg[7]  ( .D(\DataP/PC_reg/N9 ), .CK(Clk), .Q(
        IRAM_ADDRESS[5]) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[4]  ( .D(n14), .CK(Clk), .SN(Rst), .Q(
        n2778), .QN(\DataP/dest_M[4] ) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[3]  ( .D(n13), .CK(Clk), .SN(Rst), .Q(
        n2777), .QN(\DataP/dest_M[3] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[5]  ( .D(n2387), .CK(Clk), .SN(Rst), 
        .Q(n3264), .QN(\DataP/opcode_W[5] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[0]  ( .D(n2768), .CK(Clk), .SN(Rst), .Q(
        n1965), .QN(\DataP/Rs2[0] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[3]  ( .D(n2767), .CK(Clk), .SN(Rst), .QN(
        \DataP/Rs2[3] ) );
  DFFS_X1 \DataP/MEM_WB_s/RD_OUT_reg[1]  ( .D(n1637), .CK(Clk), .SN(Rst), .Q(
        n2228), .QN(\DataP/add_D[1] ) );
  DFFS_X1 \DataP/MEM_WB_s/RD_OUT_reg[3]  ( .D(n2777), .CK(Clk), .SN(Rst), .Q(
        n2775), .QN(\DataP/add_D[3] ) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[1]  ( .D(n11), .CK(Clk), .SN(Rst), .Q(
        n529), .QN(\DataP/dest_M[1] ) );
  DFFS_X1 \DataP/IF_IDs/IR_OUT_reg[30]  ( .D(IRAM_DATA_OUT[30]), .CK(Clk), 
        .SN(n36), .Q(n2377), .QN(n515) );
  DFFR_X1 \CU_I/aluOpcode1_reg[0]  ( .D(\CU_I/aluOpcode_i[0] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[0]), .QN(n2395) );
  DFFR_X1 \CU_I/aluOpcode1_reg[1]  ( .D(\CU_I/aluOpcode_i[1] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[1]), .QN(n2379) );
  DFF_X2 \DataP/PC_reg/O_reg[30]  ( .D(\DataP/PC_reg/N32 ), .CK(Clk), .Q(
        \DataP/pc_out[30] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[23]  ( .D(n2217), .CK(Clk), .SN(Rst), 
        .Q(n2413), .QN(\DataP/alu_out_M[23] ) );
  DFF_X2 \DataP/PC_reg/O_reg[26]  ( .D(\DataP/PC_reg/N28 ), .CK(Clk), .Q(
        \DataP/pc_out[26] ) );
  DFF_X2 \DataP/PC_reg/O_reg[21]  ( .D(\DataP/PC_reg/N23 ), .CK(Clk), .Q(
        \DataP/pc_out[21] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[2]  ( .D(n521), .CK(Clk), .SN(Rst), 
        .Q(n2147), .QN(\DataP/opcode_M[2] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[1]  ( .D(n2249), .CK(Clk), .SN(Rst), 
        .Q(n2776), .QN(\DataP/opcode_W[1] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[2]  ( .D(n1643), .CK(Clk), .SN(Rst), 
        .Q(n2779), .QN(\DataP/opcode_W[2] ) );
  DFFR_X1 \DataP/ID_EXs/PR_OUT_reg  ( .D(\DataP/pr_D ), .CK(Clk), .RN(Rst), 
        .Q(\DataP/pr_E ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[30]  ( .D(\DataP/imm_out[31] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[30] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[24]  ( .D(\DataP/imm_out[24] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[24] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[23]  ( .D(\DataP/imm_out[23] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[23] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[22]  ( .D(\DataP/imm_out[22] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[22] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[21]  ( .D(\DataP/imm_out[21] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[21] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[20]  ( .D(\DataP/imm_out[20] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[20] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[19]  ( .D(\DataP/imm_out[19] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[19] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[18]  ( .D(\DataP/imm_out[18] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[18] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[17]  ( .D(\DataP/imm_out[17] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[17] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[16]  ( .D(\DataP/imm_out[16] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[16] ) );
  DFFR_X1 \CU_I/aluOpcode1_reg[3]  ( .D(\CU_I/aluOpcode_i[3] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[3]), .QN(n2672) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[31]  ( .D(n2414), .CK(Clk), .SN(Rst), 
        .Q(n2517), .QN(\DataP/alu_out_W[31] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[15]  ( .D(n2433), .CK(Clk), .SN(Rst), 
        .Q(n2516), .QN(\DataP/alu_out_W[15] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[28]  ( .D(n2426), .CK(Clk), .SN(Rst), 
        .Q(n2508), .QN(\DataP/alu_out_W[28] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[24]  ( .D(n2427), .CK(Clk), .SN(Rst), 
        .Q(n2513), .QN(\DataP/alu_out_W[24] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[22]  ( .D(n2428), .CK(Clk), .SN(Rst), 
        .Q(n2512), .QN(\DataP/alu_out_W[22] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[18]  ( .D(n2425), .CK(Clk), .SN(Rst), 
        .Q(n2505), .QN(\DataP/alu_out_W[18] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[12]  ( .D(n2424), .CK(Clk), .SN(Rst), 
        .Q(n2492), .QN(\DataP/alu_out_W[12] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[25]  ( .D(n2422), .CK(Clk), .SN(Rst), 
        .Q(n2507), .QN(\DataP/alu_out_W[25] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[20]  ( .D(n2420), .CK(Clk), .SN(Rst), 
        .Q(n2506), .QN(\DataP/alu_out_W[20] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[19]  ( .D(n2421), .CK(Clk), .SN(Rst), 
        .Q(n2498), .QN(\DataP/alu_out_W[19] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[13]  ( .D(n2423), .CK(Clk), .SN(Rst), 
        .Q(n2504), .QN(\DataP/alu_out_W[13] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[30]  ( .D(n2417), .CK(Clk), .SN(Rst), 
        .Q(n2496), .QN(\DataP/alu_out_W[30] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[26]  ( .D(n2415), .CK(Clk), .SN(Rst), 
        .Q(n2500), .QN(\DataP/alu_out_W[26] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[21]  ( .D(n2419), .CK(Clk), .SN(Rst), 
        .Q(n2499), .QN(\DataP/alu_out_W[21] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[17]  ( .D(n2416), .CK(Clk), .SN(Rst), 
        .Q(n2493), .QN(\DataP/alu_out_W[17] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[14]  ( .D(n2418), .CK(Clk), .SN(Rst), 
        .Q(n2497), .QN(\DataP/alu_out_W[14] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[16]  ( .D(n2412), .CK(Clk), .SN(Rst), 
        .Q(n2511), .QN(\DataP/alu_out_W[16] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[6]  ( .D(n2410), .CK(Clk), .SN(Rst), .Q(
        n2515), .QN(\DataP/alu_out_W[6] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[2]  ( .D(n2471), .CK(Clk), .SN(Rst), .Q(
        n2514), .QN(\DataP/alu_out_W[2] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[1]  ( .D(n2469), .CK(Clk), .SN(Rst), .Q(
        n2522), .QN(\DataP/alu_out_W[1] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[7]  ( .D(n2468), .CK(Clk), .SN(Rst), .Q(
        n2510), .QN(\DataP/alu_out_W[7] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[3]  ( .D(n2478), .CK(Clk), .SN(Rst), .Q(
        n2523), .QN(\DataP/alu_out_W[3] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[10]  ( .D(n2409), .CK(Clk), .SN(Rst), 
        .Q(n2503), .QN(\DataP/alu_out_W[10] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[8]  ( .D(n2408), .CK(Clk), .SN(Rst), .Q(
        n2502), .QN(\DataP/alu_out_W[8] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[4]  ( .D(n2466), .CK(Clk), .SN(Rst), .Q(
        n2509), .QN(\DataP/alu_out_W[4] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[11]  ( .D(n2431), .CK(Clk), .SN(Rst), 
        .Q(n2518), .QN(\DataP/alu_out_W[11] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[9]  ( .D(n2477), .CK(Clk), .SN(Rst), .Q(
        n2519), .QN(\DataP/alu_out_W[9] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[5]  ( .D(n2450), .CK(Clk), .SN(Rst), .Q(
        n2520), .QN(\DataP/alu_out_W[5] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[29]  ( .D(n2008), .CK(Clk), .SN(Rst), 
        .Q(n2501), .QN(\DataP/alu_out_W[29] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[27]  ( .D(n2411), .CK(Clk), .SN(Rst), 
        .Q(n2495), .QN(\DataP/alu_out_W[27] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[23]  ( .D(n2413), .CK(Clk), .SN(Rst), 
        .Q(n2494), .QN(\DataP/alu_out_W[23] ) );
  DFFS_X1 \DataP/MEM_WB_s/ALU_OUT_reg[0]  ( .D(n2472), .CK(Clk), .SN(Rst), .Q(
        n2521), .QN(\DataP/alu_out_W[0] ) );
  DFFS_X1 \CU_I/cw1_reg[10]  ( .D(n2007), .CK(Clk), .SN(Rst), .Q(n432), .QN(
        n2475) );
  DFFS_X1 \CU_I/cw1_reg[9]  ( .D(n1961), .CK(Clk), .SN(Rst), .Q(n399), .QN(
        n2481) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[31]  ( .D(n2006), .CK(Clk), .SN(Rst), .Q(
        n2436), .QN(\DataP/A_s[31] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[6]  ( .D(n2005), .CK(Clk), .SN(Rst), .Q(
        n2462), .QN(\DataP/A_s[6] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[5]  ( .D(n2004), .CK(Clk), .SN(Rst), .Q(
        n2443), .QN(\DataP/A_s[5] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[4]  ( .D(n2003), .CK(Clk), .SN(Rst), .Q(
        n2470), .QN(\DataP/A_s[4] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[3]  ( .D(n2002), .CK(Clk), .SN(Rst), .Q(
        n2458), .QN(\DataP/A_s[3] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[30]  ( .D(n2001), .CK(Clk), .SN(Rst), .Q(
        n2437), .QN(\DataP/A_s[30] ) );
  DFFS_X1 \CU_I/aluOpcode1_reg[4]  ( .D(n2000), .CK(Clk), .SN(Rst), .Q(n443), 
        .QN(n2491) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[0]  ( .D(n1999), .CK(Clk), .SN(Rst), .Q(
        n2460), .QN(\DataP/A_s[0] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[25]  ( .D(n1998), .CK(Clk), .SN(Rst), .Q(
        n2453), .QN(\DataP/A_s[25] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[24]  ( .D(n1997), .CK(Clk), .SN(Rst), .Q(
        n2463), .QN(\DataP/A_s[24] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[23]  ( .D(n1996), .CK(Clk), .SN(Rst), .Q(
        n2439), .QN(\DataP/A_s[23] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[22]  ( .D(n1995), .CK(Clk), .SN(Rst), .Q(
        n2464), .QN(\DataP/A_s[22] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[21]  ( .D(n1994), .CK(Clk), .SN(Rst), .Q(
        n2446), .QN(\DataP/A_s[21] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[20]  ( .D(n1993), .CK(Clk), .SN(Rst), .Q(
        n2454), .QN(\DataP/A_s[20] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[19]  ( .D(n1992), .CK(Clk), .SN(Rst), .Q(
        n2447), .QN(\DataP/A_s[19] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[18]  ( .D(n1991), .CK(Clk), .SN(Rst), .Q(
        n2455), .QN(\DataP/A_s[18] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[17]  ( .D(n1990), .CK(Clk), .SN(Rst), .Q(
        n2440), .QN(\DataP/A_s[17] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[16]  ( .D(n1989), .CK(Clk), .SN(Rst), .Q(
        n2465), .QN(\DataP/A_s[16] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[15]  ( .D(n1988), .CK(Clk), .SN(Rst), .Q(
        n2441), .QN(\DataP/A_s[15] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[14]  ( .D(n1987), .CK(Clk), .SN(Rst), .Q(
        n2448), .QN(\DataP/A_s[14] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[13]  ( .D(n1986), .CK(Clk), .SN(Rst), .Q(
        n2456), .QN(\DataP/A_s[13] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[12]  ( .D(n1985), .CK(Clk), .SN(Rst), .Q(
        n2442), .QN(\DataP/A_s[12] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[11]  ( .D(n1984), .CK(Clk), .SN(Rst), .Q(
        n2449), .QN(\DataP/A_s[11] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[10]  ( .D(n1983), .CK(Clk), .SN(Rst), .Q(
        n2457), .QN(\DataP/A_s[10] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[7]  ( .D(n1982), .CK(Clk), .SN(Rst), .Q(
        n2451), .QN(\DataP/A_s[7] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[1]  ( .D(n1981), .CK(Clk), .SN(Rst), .Q(
        n2461), .QN(\DataP/A_s[1] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[28]  ( .D(n1980), .CK(Clk), .SN(Rst), .Q(
        n2452), .QN(\DataP/A_s[28] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[26]  ( .D(n1979), .CK(Clk), .SN(Rst), .Q(
        n2445), .QN(\DataP/A_s[26] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[29]  ( .D(n1978), .CK(Clk), .SN(Rst), .Q(
        n2444), .QN(\DataP/A_s[29] ) );
  DFFS_X1 \DataP/ID_EXs/A_OUT_reg[27]  ( .D(n1977), .CK(Clk), .SN(Rst), .Q(
        n2438), .QN(\DataP/A_s[27] ) );
  DFFRS_X1 \DataP/PC_reg/O_reg[11]  ( .D(\DataP/PC_reg/N13 ), .CK(Clk), .RN(
        1'b1), .SN(1'b1), .Q(\DataP/pc_out[11] ) );
  DFFR_X1 \DataP/ID_EXs/NPC_L_OUT_reg[31]  ( .D(\DataP/link_addr_D[31] ), .CK(
        Clk), .RN(Rst), .QN(n292) );
  DFFRS_X1 \DataP/PC_reg/O_reg[20]  ( .D(\DataP/PC_reg/N22 ), .CK(Clk), .RN(
        1'b1), .SN(1'b1), .Q(\DataP/pc_out[20] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[1]  ( .D(n2770), .CK(Clk), .SN(Rst), .QN(
        \DataP/Rs2[1] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[29]  ( .D(n299), .CK(Clk), .SN(Rst), .Q(
        n2008), .QN(\DataP/alu_out_M[29] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[4]  ( .D(n2769), .CK(Clk), .SN(Rst), .Q(
        n2029), .QN(\DataP/Rs2[4] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[2]  ( .D(n1974), .CK(Clk), .SN(Rst), .Q(
        n1603), .QN(\DataP/Rs2[2] ) );
  DFFR_X1 \DataP/MEM_WB_s/RD_OUT_reg[4]  ( .D(n1720), .CK(Clk), .RN(Rst), .Q(
        \DataP/add_D[4] ), .QN(n540) );
  DFFR_X1 \DataP/ID_EXs/OPCODE_OUT_reg[5]  ( .D(IR_CU_31), .CK(Clk), .RN(Rst), 
        .QN(n17) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[27]  ( .D(IRAM_DATA_OUT[27]), .CK(Clk), 
        .RN(n36), .Q(IR_CU_27), .QN(n504) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[0]  ( .D(n2243), .CK(Clk), .SN(Rst), .Q(
        n2472), .QN(DRAM_ADDRESS[0]) );
  DFF_X1 \DataP/PC_reg/O_reg[28]  ( .D(\DataP/PC_reg/N30 ), .CK(Clk), .Q(
        \DataP/pc_out[28] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[27]  ( .D(n301), .CK(Clk), .SN(Rst), .Q(
        n2411), .QN(\DataP/alu_out_M[27] ) );
  DFF_X1 \DataP/PC_reg/O_reg[15]  ( .D(\DataP/PC_reg/N17 ), .CK(Clk), .Q(
        \DataP/pc_out[15] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[22]  ( .D(n1708), .CK(Clk), .SN(Rst), 
        .Q(n2428), .QN(\DataP/alu_out_M[22] ) );
  DFFR_X1 \DataP/ID_EXs/OPCODE_OUT_reg[2]  ( .D(IR_CU_28), .CK(Clk), .RN(Rst), 
        .QN(n521) );
  DFF_X2 \DataP/PC_reg/O_reg[25]  ( .D(\DataP/PC_reg/N27 ), .CK(Clk), .Q(
        \DataP/pc_out[25] ) );
  DFF_X1 \DataP/PC_reg/O_reg[24]  ( .D(\DataP/PC_reg/N26 ), .CK(Clk), .Q(
        \DataP/pc_out[24] ) );
  DFF_X1 \DataP/PC_reg/O_reg[17]  ( .D(\DataP/PC_reg/N19 ), .CK(Clk), .Q(
        \DataP/pc_out[17] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[26]  ( .D(n1598), .CK(Clk), .SN(Rst), 
        .Q(n2415), .QN(\DataP/alu_out_M[26] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[17]  ( .D(n1611), .CK(Clk), .SN(Rst), 
        .Q(n2416), .QN(\DataP/alu_out_M[17] ) );
  DFF_X1 \DataP/PC_reg/O_reg[0]  ( .D(\DataP/PC_reg/N2 ), .CK(Clk), .Q(
        \DataP/pc_out_0 ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[7]  ( .D(n1569), .CK(Clk), .SN(Rst), .Q(
        n2468), .QN(DRAM_ADDRESS[7]) );
  DFF_X1 \DataP/PC_reg/O_reg[29]  ( .D(\DataP/PC_reg/N31 ), .CK(Clk), .Q(
        \DataP/pc_out[29] ) );
  NOR2_X1 U1484 ( .A1(n3294), .A2(n3234), .ZN(n3909) );
  INV_X2 U1485 ( .A(n3880), .ZN(n2129) );
  NAND2_X1 U1486 ( .A1(n3689), .A2(\DataP/alu_a_in[23] ), .ZN(n1548) );
  NOR2_X1 U1487 ( .A1(\DataP/alu_b_in[8] ), .A2(n1577), .ZN(n1549) );
  NAND4_X1 U1488 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(n1550)
         );
  OAI211_X1 U1489 ( .C1(n3662), .C2(n3682), .A(n1566), .B(n2169), .ZN(n1551)
         );
  AND2_X2 U1490 ( .A1(n2527), .A2(n1570), .ZN(n3662) );
  NAND2_X1 U1491 ( .A1(n2667), .A2(n2665), .ZN(n1552) );
  NAND2_X1 U1492 ( .A1(n2532), .A2(n3730), .ZN(n2531) );
  NAND2_X1 U1493 ( .A1(n1553), .A2(n1554), .ZN(\DataP/alu_a_in[0] ) );
  INV_X1 U1494 ( .A(n3331), .ZN(n1553) );
  INV_X1 U1495 ( .A(n3332), .ZN(n1554) );
  AND2_X1 U1496 ( .A1(n3661), .A2(n3660), .ZN(n2219) );
  AOI21_X1 U1497 ( .B1(\DataP/alu_a_in[4] ), .B2(n2380), .A(n1922), .ZN(n2256)
         );
  NAND2_X1 U1498 ( .A1(n2727), .A2(n3797), .ZN(n2718) );
  NAND3_X1 U1499 ( .A1(n1552), .A2(n2718), .A3(n2713), .ZN(n1555) );
  AND2_X2 U1500 ( .A1(n2727), .A2(n3797), .ZN(n2382) );
  NAND2_X1 U1501 ( .A1(n2745), .A2(n2071), .ZN(n1556) );
  NOR2_X1 U1502 ( .A1(n2746), .A2(n3826), .ZN(n1557) );
  XNOR2_X1 U1503 ( .A(n1556), .B(n1557), .ZN(n1558) );
  AOI21_X1 U1504 ( .B1(n1558), .B2(n2129), .A(n3833), .ZN(n299) );
  NAND2_X1 U1505 ( .A1(n1558), .A2(n1607), .ZN(n1659) );
  NOR2_X1 U1506 ( .A1(n1559), .A2(n1838), .ZN(n3423) );
  NAND4_X1 U1507 ( .A1(n2658), .A2(n1587), .A3(n2660), .A4(n1595), .ZN(n1559)
         );
  NOR2_X1 U1508 ( .A1(\sra_131/SH[4] ), .A2(n1559), .ZN(n1704) );
  AND4_X1 U1509 ( .A1(n1560), .A2(n1561), .A3(n1562), .A4(n1563), .ZN(n4103)
         );
  AND3_X1 U1510 ( .A1(n3707), .A2(n3898), .A3(n3875), .ZN(n1560) );
  AND4_X1 U1511 ( .A1(n3741), .A2(n3731), .A3(n3872), .A4(n3613), .ZN(n1561)
         );
  AND4_X1 U1512 ( .A1(n3859), .A2(n3853), .A3(n3603), .A4(n3536), .ZN(n1562)
         );
  AND3_X1 U1513 ( .A1(n3542), .A2(n3541), .A3(n3848), .ZN(n1563) );
  OAI211_X1 U1514 ( .C1(n2728), .C2(n2382), .A(n1555), .B(n2712), .ZN(n1564)
         );
  NAND3_X1 U1515 ( .A1(n2192), .A2(n3690), .A3(n2193), .ZN(n1565) );
  BUF_X2 U1516 ( .A(n2233), .Z(n2226) );
  CLKBUF_X3 U1517 ( .A(n3401), .Z(n3213) );
  AOI211_X4 U1518 ( .C1(n2299), .C2(n2289), .A(n2287), .B(n2288), .ZN(n2290)
         );
  MUX2_X2 U1519 ( .A(n3413), .B(n3200), .S(n3886), .Z(n3414) );
  AND2_X1 U1520 ( .A1(n3685), .A2(n3649), .ZN(n1566) );
  AND2_X1 U1521 ( .A1(n3685), .A2(n3649), .ZN(n3684) );
  NAND2_X1 U1522 ( .A1(n2077), .A2(n1593), .ZN(n1567) );
  INV_X2 U1523 ( .A(n2072), .ZN(n3207) );
  NOR2_X1 U1524 ( .A1(n2659), .A2(n2090), .ZN(n1568) );
  AOI211_X1 U1525 ( .C1(n3228), .C2(n1909), .A(n1914), .B(n1918), .ZN(n1569)
         );
  AOI211_X1 U1526 ( .C1(n3228), .C2(n1909), .A(n1914), .B(n1918), .ZN(n350) );
  NAND2_X1 U1527 ( .A1(n2173), .A2(n2528), .ZN(n1570) );
  AND3_X1 U1528 ( .A1(n1636), .A2(n3681), .A3(n3686), .ZN(n1571) );
  AND3_X1 U1529 ( .A1(n1636), .A2(n3681), .A3(n3686), .ZN(n3712) );
  BUF_X1 U1530 ( .A(n3221), .Z(n1572) );
  AND4_X1 U1531 ( .A1(n3478), .A2(n3477), .A3(n3475), .A4(n3476), .ZN(n1573)
         );
  AND2_X2 U1532 ( .A1(n2723), .A2(n1599), .ZN(n1574) );
  AND2_X1 U1533 ( .A1(n2723), .A2(n1599), .ZN(n3709) );
  BUF_X2 U1534 ( .A(\DataP/alu_b_in[11] ), .Z(n2151) );
  BUF_X1 U1535 ( .A(\DataP/alu_b_in[8] ), .Z(n1575) );
  INV_X2 U1536 ( .A(n1753), .ZN(\DataP/alu_b_in[17] ) );
  BUF_X1 U1537 ( .A(n2188), .Z(n1576) );
  BUF_X1 U1538 ( .A(\DataP/alu_b_in[9] ), .Z(n1577) );
  OAI211_X1 U1539 ( .C1(n2772), .C2(n2478), .A(n2661), .B(n2662), .ZN(n1578)
         );
  BUF_X2 U1540 ( .A(\DataP/alu_b_in[10] ), .Z(n2165) );
  AND2_X1 U1541 ( .A1(n2657), .A2(n2656), .ZN(n1579) );
  AND4_X1 U1542 ( .A1(n3317), .A2(n3318), .A3(n3316), .A4(n3315), .ZN(n2380)
         );
  NAND2_X1 U1543 ( .A1(n1709), .A2(n1580), .ZN(n3694) );
  NOR2_X1 U1544 ( .A1(n3641), .A2(n3640), .ZN(n1580) );
  NAND2_X1 U1545 ( .A1(n2076), .A2(n1580), .ZN(n1760) );
  OAI211_X2 U1546 ( .C1(n2427), .C2(n2771), .A(n1841), .B(n1842), .ZN(
        \DataP/alu_b_in[24] ) );
  BUF_X2 U1547 ( .A(n3548), .Z(n1581) );
  AND2_X1 U1548 ( .A1(\DataP/alu_b_in[18] ), .A2(n1694), .ZN(n2731) );
  INV_X2 U1549 ( .A(n3201), .ZN(n3048) );
  AOI21_X1 U1550 ( .B1(n3635), .B2(n3636), .A(n2715), .ZN(n1582) );
  NAND2_X1 U1551 ( .A1(n2246), .A2(\DataP/IMM_s[1] ), .ZN(n1583) );
  NAND2_X1 U1552 ( .A1(\DataP/alu_b_in[16] ), .A2(n2535), .ZN(n2534) );
  NAND2_X1 U1553 ( .A1(n1644), .A2(n1662), .ZN(n1584) );
  AND2_X1 U1554 ( .A1(n3449), .A2(\DataP/alu_a_in[10] ), .ZN(n3489) );
  NAND4_X1 U1555 ( .A1(n1568), .A2(n1587), .A3(n1595), .A4(n1586), .ZN(n1585)
         );
  INV_X1 U1556 ( .A(n1578), .ZN(n1586) );
  AND2_X1 U1557 ( .A1(n2656), .A2(n2657), .ZN(n1587) );
  NAND2_X1 U1558 ( .A1(n3666), .A2(\DataP/alu_a_in[20] ), .ZN(n1588) );
  AND2_X1 U1559 ( .A1(n2154), .A2(n2153), .ZN(n1589) );
  OAI211_X1 U1560 ( .C1(n2604), .C2(n2607), .A(n2603), .B(n3686), .ZN(n1590)
         );
  OR2_X1 U1561 ( .A1(n3295), .A2(n1718), .ZN(n1673) );
  INV_X1 U1562 ( .A(n3429), .ZN(n1591) );
  OAI211_X1 U1563 ( .C1(n2728), .C2(n2382), .A(n2711), .B(n2712), .ZN(n1592)
         );
  AND2_X1 U1564 ( .A1(n3308), .A2(n3309), .ZN(n1593) );
  OAI21_X1 U1565 ( .B1(n2596), .B2(n2535), .A(n2701), .ZN(n1594) );
  AND4_X1 U1566 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n1595)
         );
  AND4_X1 U1567 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n2240)
         );
  CLKBUF_X3 U1568 ( .A(n2773), .Z(n1627) );
  AND2_X1 U1569 ( .A1(n3683), .A2(n1663), .ZN(n1596) );
  NAND2_X1 U1570 ( .A1(n1683), .A2(n3721), .ZN(n2583) );
  XNOR2_X1 U1571 ( .A(\DataP/Rs2[3] ), .B(\DataP/add_D[3] ), .ZN(n1962) );
  XOR2_X1 U1572 ( .A(\lt_x_135/B[12] ), .B(n1941), .Z(n1597) );
  NOR2_X2 U1573 ( .A1(n2068), .A2(n3480), .ZN(n1941) );
  BUF_X1 U1574 ( .A(n303), .Z(n1598) );
  NOR2_X1 U1575 ( .A1(n3659), .A2(n1737), .ZN(n1599) );
  BUF_X1 U1576 ( .A(\DataP/alu_b_in[19] ), .Z(n1600) );
  CLKBUF_X3 U1577 ( .A(n3401), .Z(n3214) );
  BUF_X1 U1578 ( .A(n2250), .Z(n1601) );
  INV_X1 U1579 ( .A(n2074), .ZN(\lt_x_135/B[5] ) );
  INV_X2 U1580 ( .A(n3886), .ZN(n2108) );
  OR2_X1 U1581 ( .A1(n1732), .A2(n2322), .ZN(n1602) );
  INV_X1 U1582 ( .A(n3886), .ZN(n1694) );
  AND2_X1 U1583 ( .A1(\DataP/alu_a_in[24] ), .A2(n1691), .ZN(n1604) );
  AND2_X1 U1584 ( .A1(n1904), .A2(n3717), .ZN(n1605) );
  AND2_X1 U1585 ( .A1(n2129), .A2(n1656), .ZN(n1607) );
  NAND2_X1 U1586 ( .A1(n3540), .A2(n1696), .ZN(n1608) );
  NAND2_X1 U1587 ( .A1(n1904), .A2(n2727), .ZN(n1609) );
  XOR2_X1 U1588 ( .A(n1830), .B(n2030), .Z(n1610) );
  BUF_X1 U1589 ( .A(n323), .Z(n1611) );
  XNOR2_X1 U1590 ( .A(n1612), .B(n2404), .ZN(n3796) );
  NAND2_X1 U1591 ( .A1(n1626), .A2(n1548), .ZN(n1612) );
  NAND2_X1 U1592 ( .A1(n2697), .A2(n2696), .ZN(n1613) );
  NAND2_X1 U1593 ( .A1(n2697), .A2(n2696), .ZN(n3777) );
  BUF_X1 U1594 ( .A(n1581), .Z(n1614) );
  OAI21_X1 U1595 ( .B1(n2681), .B2(n2128), .A(n2680), .ZN(n1615) );
  OR2_X4 U1596 ( .A1(n3343), .A2(n3342), .ZN(\DataP/alu_a_in[6] ) );
  NAND2_X1 U1597 ( .A1(n1615), .A2(\DataP/alu_a_in[6] ), .ZN(n1616) );
  NAND2_X1 U1598 ( .A1(n3609), .A2(n1616), .ZN(n3855) );
  INV_X1 U1599 ( .A(\DataP/alu_a_in[6] ), .ZN(n3857) );
  AND2_X1 U1600 ( .A1(n3884), .A2(n2489), .ZN(n1617) );
  AND2_X1 U1601 ( .A1(n3884), .A2(n2489), .ZN(n1618) );
  AND2_X1 U1602 ( .A1(n1571), .A2(n1582), .ZN(n1619) );
  BUF_X1 U1603 ( .A(n3221), .Z(n1620) );
  NAND2_X1 U1604 ( .A1(n1679), .A2(n3718), .ZN(n3799) );
  BUF_X1 U1605 ( .A(\DataP/dest_M[3] ), .Z(n1621) );
  BUF_X1 U1606 ( .A(n3575), .Z(n1622) );
  BUF_X1 U1607 ( .A(n1581), .Z(n1623) );
  BUF_X1 U1608 ( .A(n304), .Z(n1624) );
  BUF_X1 U1609 ( .A(\DataP/dest_M[4] ), .Z(n1625) );
  NAND3_X1 U1610 ( .A1(n2192), .A2(n3690), .A3(n2133), .ZN(n1626) );
  BUF_X2 U1611 ( .A(n2781), .Z(n2773) );
  BUF_X1 U1612 ( .A(n540), .Z(n1628) );
  INV_X1 U1613 ( .A(n1628), .ZN(n1629) );
  BUF_X1 U1614 ( .A(n536), .Z(n1630) );
  BUF_X1 U1615 ( .A(n3221), .Z(n1631) );
  BUF_X1 U1616 ( .A(n3796), .Z(n1632) );
  NAND2_X1 U1617 ( .A1(n1590), .A2(n2608), .ZN(n1633) );
  NOR2_X1 U1618 ( .A1(n3861), .A2(n3868), .ZN(n1634) );
  BUF_X1 U1619 ( .A(n2241), .Z(n1635) );
  BUF_X1 U1620 ( .A(n1551), .Z(n1636) );
  INV_X1 U1621 ( .A(\DataP/dest_M[1] ), .ZN(n1637) );
  OR2_X1 U1622 ( .A1(n2190), .A2(\DataP/alu_a_in[26] ), .ZN(n3719) );
  INV_X1 U1623 ( .A(\DataP/dest_M[2] ), .ZN(n1638) );
  NAND2_X1 U1624 ( .A1(\DataP/Rs2[4] ), .A2(\DataP/add_D[4] ), .ZN(n1641) );
  NAND2_X1 U1625 ( .A1(n1639), .A2(n1640), .ZN(n1642) );
  NAND2_X1 U1626 ( .A1(n1641), .A2(n1642), .ZN(n3245) );
  INV_X1 U1627 ( .A(\DataP/Rs2[4] ), .ZN(n1639) );
  INV_X1 U1628 ( .A(\DataP/add_D[4] ), .ZN(n1640) );
  INV_X1 U1629 ( .A(\DataP/opcode_M[2] ), .ZN(n1643) );
  BUF_X1 U1630 ( .A(n3845), .Z(n1644) );
  BUF_X1 U1631 ( .A(n3221), .Z(n1645) );
  BUF_X1 U1632 ( .A(n1571), .Z(n1646) );
  BUF_X1 U1633 ( .A(n3642), .Z(n1647) );
  BUF_X1 U1634 ( .A(n3609), .Z(n1648) );
  AND2_X1 U1635 ( .A1(n538), .A2(n540), .ZN(n1649) );
  NAND4_X1 U1636 ( .A1(n1757), .A2(n1649), .A3(n2228), .A4(n1630), .ZN(n1650)
         );
  AND2_X1 U1637 ( .A1(n3289), .A2(n1650), .ZN(n1651) );
  NAND3_X1 U1638 ( .A1(n1742), .A2(n3290), .A3(n1651), .ZN(n3293) );
  NAND2_X1 U1639 ( .A1(n3245), .A2(n1650), .ZN(n2637) );
  INV_X1 U1640 ( .A(n1650), .ZN(n1671) );
  INV_X1 U1641 ( .A(n2228), .ZN(n2229) );
  XNOR2_X1 U1642 ( .A(n2249), .B(n2147), .ZN(n1652) );
  NOR2_X1 U1643 ( .A1(n1652), .A2(n18), .ZN(n1653) );
  AND2_X1 U1644 ( .A1(n2195), .A2(n2387), .ZN(n1654) );
  OAI21_X1 U1645 ( .B1(n1653), .B2(n1654), .A(\DataP/opcode_M[3] ), .ZN(n3250)
         );
  NAND2_X1 U1646 ( .A1(n2040), .A2(n1968), .ZN(n1655) );
  NAND2_X1 U1647 ( .A1(n1659), .A2(n1658), .ZN(\DataP/PC_reg/N31 ) );
  INV_X2 U1648 ( .A(n4111), .ZN(n1656) );
  NOR2_X2 U1649 ( .A1(n4110), .A2(n4193), .ZN(n1657) );
  AOI21_X2 U1650 ( .B1(n3833), .B2(n2131), .A(n1657), .ZN(n1658) );
  NAND2_X1 U1651 ( .A1(n1661), .A2(n1660), .ZN(n3629) );
  AND2_X1 U1652 ( .A1(n2109), .A2(n2740), .ZN(n1660) );
  NAND2_X1 U1653 ( .A1(n3619), .A2(n2108), .ZN(n1661) );
  BUF_X1 U1654 ( .A(n3548), .Z(n3222) );
  AND3_X1 U1655 ( .A1(n2194), .A2(n2094), .A3(n1579), .ZN(n1755) );
  BUF_X1 U1656 ( .A(n3844), .Z(n1662) );
  NAND2_X4 U1657 ( .A1(n3908), .A2(Rst), .ZN(n4111) );
  BUF_X1 U1658 ( .A(n2239), .Z(n1663) );
  OAI21_X1 U1659 ( .B1(n313), .B2(n4111), .A(n1664), .ZN(\DataP/PC_reg/N23 )
         );
  OR2_X1 U1660 ( .A1(n4110), .A2(n4201), .ZN(n1664) );
  OAI22_X1 U1661 ( .A1(n2678), .A2(n2677), .B1(\DataP/alu_a_in[21] ), .B2(
        n2679), .ZN(n2653) );
  NAND2_X1 U1662 ( .A1(n2599), .A2(n2630), .ZN(n2678) );
  NAND2_X1 U1663 ( .A1(n2745), .A2(n2071), .ZN(n2083) );
  NAND2_X1 U1664 ( .A1(n1592), .A2(n2717), .ZN(n2745) );
  OAI211_X1 U1665 ( .C1(n3214), .C2(n37), .A(n1666), .B(n1665), .ZN(n3332) );
  NAND2_X1 U1666 ( .A1(n3209), .A2(\DataP/alu_out_W[0] ), .ZN(n1665) );
  NAND2_X1 U1667 ( .A1(n3210), .A2(DRAM_ADDRESS[0]), .ZN(n1666) );
  XNOR2_X1 U1668 ( .A(n3423), .B(n1748), .ZN(n2681) );
  NAND2_X1 U1669 ( .A1(n1668), .A2(n1667), .ZN(n2430) );
  NOR2_X1 U1670 ( .A1(n3885), .A2(n2385), .ZN(n1667) );
  INV_X1 U1671 ( .A(n3722), .ZN(n1668) );
  XNOR2_X1 U1672 ( .A(n1603), .B(n538), .ZN(n2143) );
  NAND3_X1 U1673 ( .A1(n3294), .A2(n3290), .A3(n1669), .ZN(n3279) );
  OR2_X1 U1674 ( .A1(n3279), .A2(n1743), .ZN(n2634) );
  NAND4_X1 U1675 ( .A1(n3292), .A2(n1673), .A3(n1672), .A4(n2634), .ZN(n3401)
         );
  NOR2_X2 U1676 ( .A1(n1671), .A2(n1670), .ZN(n1669) );
  INV_X2 U1677 ( .A(Rst), .ZN(n1670) );
  AOI21_X1 U1678 ( .B1(n3909), .B2(n2619), .A(n432), .ZN(n1672) );
  NAND2_X1 U1679 ( .A1(n2663), .A2(n2564), .ZN(n2590) );
  XNOR2_X1 U1680 ( .A(n1675), .B(n1674), .ZN(n2663) );
  INV_X1 U1681 ( .A(n1576), .ZN(n1674) );
  AOI21_X1 U1682 ( .B1(n1565), .B2(n1677), .A(n1676), .ZN(n1675) );
  INV_X1 U1683 ( .A(n3719), .ZN(n1676) );
  AND2_X1 U1684 ( .A1(n2705), .A2(n2584), .ZN(n1677) );
  NAND2_X1 U1685 ( .A1(n2664), .A2(n2720), .ZN(n2595) );
  AND2_X2 U1686 ( .A1(n1609), .A2(n1678), .ZN(n2664) );
  NAND3_X1 U1687 ( .A1(n1605), .A2(n1744), .A3(n2729), .ZN(n1678) );
  NAND3_X1 U1688 ( .A1(n2729), .A2(n1744), .A3(n3717), .ZN(n1679) );
  NAND2_X1 U1689 ( .A1(n2188), .A2(n1680), .ZN(n1683) );
  OR2_X1 U1690 ( .A1(n2096), .A2(n3719), .ZN(n1680) );
  AOI21_X1 U1691 ( .B1(n1681), .B2(n2582), .A(n2746), .ZN(n1682) );
  NAND2_X1 U1692 ( .A1(n1683), .A2(n3721), .ZN(n1681) );
  NAND2_X1 U1693 ( .A1(n2748), .A2(n1682), .ZN(n2021) );
  NAND2_X2 U1694 ( .A1(n2583), .A2(n2582), .ZN(n2766) );
  NAND2_X2 U1695 ( .A1(n1686), .A2(n2535), .ZN(n2585) );
  NAND2_X2 U1696 ( .A1(\DataP/alu_a_in[25] ), .A2(n1684), .ZN(n1821) );
  NOR2_X2 U1697 ( .A1(n2588), .A2(n3851), .ZN(n1684) );
  OAI21_X2 U1698 ( .B1(\DataP/alu_a_in[25] ), .B2(n1686), .A(n3894), .ZN(n1820) );
  XNOR2_X2 U1699 ( .A(\DataP/alu_a_in[25] ), .B(n1686), .ZN(n3800) );
  NOR2_X2 U1700 ( .A1(n2137), .A2(n1686), .ZN(n2282) );
  AOI21_X2 U1701 ( .B1(n2283), .B2(\DataP/alu_b_in[24] ), .A(n1685), .ZN(n2356) );
  AND2_X2 U1702 ( .A1(n2137), .A2(n1686), .ZN(n1685) );
  INV_X2 U1703 ( .A(n2588), .ZN(n1686) );
  NOR2_X2 U1704 ( .A1(n1688), .A2(n1687), .ZN(n2588) );
  NAND2_X2 U1705 ( .A1(n3504), .A2(n3505), .ZN(n1687) );
  NAND2_X2 U1706 ( .A1(n3506), .A2(n3523), .ZN(n1688) );
  OAI21_X1 U1707 ( .B1(n3695), .B2(n1692), .A(n1604), .ZN(n3718) );
  AOI21_X2 U1708 ( .B1(n3695), .B2(n1694), .A(n1689), .ZN(n3788) );
  NAND2_X2 U1709 ( .A1(n1690), .A2(n1693), .ZN(n1689) );
  INV_X2 U1710 ( .A(\DataP/alu_a_in[24] ), .ZN(n1690) );
  NAND2_X2 U1711 ( .A1(n1693), .A2(n1698), .ZN(n1691) );
  INV_X2 U1712 ( .A(n1693), .ZN(n1692) );
  NAND2_X2 U1713 ( .A1(\DataP/alu_b_in[24] ), .A2(n3886), .ZN(n1693) );
  OAI211_X1 U1714 ( .C1(n3462), .C2(n1696), .A(n1695), .B(n1608), .ZN(n3464)
         );
  OR2_X2 U1715 ( .A1(n3467), .A2(n1696), .ZN(n1695) );
  AND2_X2 U1716 ( .A1(n3464), .A2(n3491), .ZN(n3488) );
  NAND2_X1 U1717 ( .A1(n3488), .A2(n3489), .ZN(n2612) );
  INV_X2 U1718 ( .A(n2108), .ZN(n1696) );
  OAI21_X1 U1719 ( .B1(n3448), .B2(n1698), .A(n1697), .ZN(n3449) );
  NAND2_X1 U1720 ( .A1(n2165), .A2(n1698), .ZN(n1697) );
  INV_X1 U1721 ( .A(n2108), .ZN(n1698) );
  XNOR2_X1 U1722 ( .A(n3460), .B(n3459), .ZN(n3448) );
  AND2_X1 U1723 ( .A1(n2076), .A2(n1549), .ZN(n3460) );
  OAI21_X1 U1724 ( .B1(n2083), .B2(n1699), .A(n2552), .ZN(n2551) );
  NAND2_X1 U1725 ( .A1(n1701), .A2(n1700), .ZN(n1699) );
  INV_X1 U1726 ( .A(n4111), .ZN(n1700) );
  INV_X1 U1727 ( .A(n2752), .ZN(n1701) );
  NAND2_X1 U1728 ( .A1(n1703), .A2(n1702), .ZN(n2752) );
  INV_X1 U1729 ( .A(n2704), .ZN(n1702) );
  NAND2_X1 U1730 ( .A1(n1617), .A2(n3826), .ZN(n1703) );
  OAI21_X1 U1731 ( .B1(n2044), .B2(n2128), .A(n2163), .ZN(n3421) );
  XNOR2_X1 U1732 ( .A(n1704), .B(\lt_x_135/B[5] ), .ZN(n2044) );
  NAND2_X1 U1733 ( .A1(n2687), .A2(n2686), .ZN(n3836) );
  NAND2_X1 U1734 ( .A1(n1705), .A2(n2108), .ZN(n2687) );
  XNOR2_X1 U1735 ( .A(n3642), .B(n3841), .ZN(n1705) );
  INV_X1 U1736 ( .A(n3642), .ZN(n3480) );
  XNOR2_X1 U1737 ( .A(n1613), .B(n3776), .ZN(n1706) );
  BUF_X1 U1738 ( .A(n3662), .Z(n1707) );
  AOI21_X1 U1739 ( .B1(n1706), .B2(n2129), .A(n3786), .ZN(n1708) );
  AND2_X1 U1740 ( .A1(n1755), .A2(n2093), .ZN(n1709) );
  AND2_X2 U1741 ( .A1(n2075), .A2(n2027), .ZN(n2245) );
  BUF_X1 U1742 ( .A(n3864), .Z(n1710) );
  AND2_X2 U1743 ( .A1(n2093), .A2(n2092), .ZN(n2075) );
  NAND2_X1 U1744 ( .A1(n2191), .A2(n2705), .ZN(n1711) );
  AND2_X1 U1745 ( .A1(n1730), .A2(n1758), .ZN(n1712) );
  XNOR2_X1 U1746 ( .A(n3618), .B(n2106), .ZN(n1713) );
  XOR2_X1 U1747 ( .A(n3461), .B(n2151), .Z(n1714) );
  BUF_X1 U1748 ( .A(n2242), .Z(n1748) );
  AND4_X2 U1749 ( .A1(n2660), .A2(n2242), .A3(n2372), .A4(n2240), .ZN(n2093)
         );
  INV_X1 U1750 ( .A(n2232), .ZN(n1715) );
  BUF_X1 U1751 ( .A(n2240), .Z(n1716) );
  OR2_X1 U1752 ( .A1(n3669), .A2(n2631), .ZN(n2599) );
  NAND2_X1 U1753 ( .A1(n2568), .A2(n2487), .ZN(n1717) );
  OR2_X1 U1754 ( .A1(n3294), .A2(n3234), .ZN(n1718) );
  NOR2_X2 U1755 ( .A1(n3330), .A2(n3329), .ZN(n1719) );
  BUF_X2 U1756 ( .A(n3548), .Z(n3223) );
  NAND4_X4 U1757 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(
        \DataP/alu_b_in[20] ) );
  INV_X1 U1758 ( .A(n2778), .ZN(n1720) );
  CLKBUF_X3 U1759 ( .A(n3402), .Z(n3216) );
  AOI21_X1 U1760 ( .B1(n1617), .B2(n3826), .A(n2704), .ZN(n1721) );
  INV_X1 U1761 ( .A(n2732), .ZN(n1722) );
  BUF_X1 U1762 ( .A(n3763), .Z(n1723) );
  OAI211_X1 U1763 ( .C1(n2421), .C2(n2771), .A(n1928), .B(n1929), .ZN(
        \DataP/alu_b_in[19] ) );
  OAI211_X1 U1764 ( .C1(n2598), .C2(n2599), .A(n2530), .B(n2490), .ZN(n3763)
         );
  AND2_X1 U1765 ( .A1(n3601), .A2(n2082), .ZN(n1724) );
  AND2_X1 U1766 ( .A1(n3601), .A2(n2082), .ZN(n1725) );
  AND2_X1 U1767 ( .A1(n3601), .A2(n2082), .ZN(n2194) );
  BUF_X1 U1768 ( .A(n2735), .Z(n1726) );
  AND4_X2 U1769 ( .A1(n3321), .A2(n3322), .A3(n3319), .A4(n3320), .ZN(n3601)
         );
  NAND2_X1 U1770 ( .A1(n1727), .A2(n3585), .ZN(n3844) );
  NAND2_X1 U1771 ( .A1(n3588), .A2(n3586), .ZN(n1727) );
  NAND2_X1 U1772 ( .A1(n1719), .A2(n3417), .ZN(n3586) );
  NAND2_X1 U1773 ( .A1(n1729), .A2(n3575), .ZN(n3588) );
  XNOR2_X1 U1774 ( .A(n1926), .B(n1728), .ZN(n3417) );
  INV_X1 U1775 ( .A(n1716), .ZN(n1728) );
  NAND2_X1 U1776 ( .A1(n3574), .A2(n3577), .ZN(n1729) );
  NAND2_X1 U1777 ( .A1(n3415), .A2(n2232), .ZN(n3575) );
  NAND2_X1 U1778 ( .A1(n1730), .A2(n1758), .ZN(n3849) );
  NAND2_X1 U1779 ( .A1(n1731), .A2(n2108), .ZN(n1730) );
  XNOR2_X1 U1780 ( .A(n1585), .B(\sra_131/SH[4] ), .ZN(n1731) );
  AND2_X1 U1781 ( .A1(n3459), .A2(\DataP/alu_a_in[10] ), .ZN(n1732) );
  BUF_X1 U1782 ( .A(n3572), .Z(n1733) );
  OR2_X4 U1783 ( .A1(n3404), .A2(n3403), .ZN(\DataP/alu_a_in[10] ) );
  INV_X4 U1784 ( .A(n2138), .ZN(n2102) );
  BUF_X4 U1785 ( .A(\sra_131/SH[4] ), .Z(n2138) );
  NAND2_X1 U1786 ( .A1(n2549), .A2(n2547), .ZN(n1734) );
  NOR2_X1 U1787 ( .A1(n3659), .A2(n1737), .ZN(n1735) );
  INV_X1 U1788 ( .A(n2123), .ZN(n1736) );
  NOR2_X1 U1789 ( .A1(n3659), .A2(n1737), .ZN(n3691) );
  OAI211_X1 U1790 ( .C1(n2425), .C2(n1627), .A(n1901), .B(n1900), .ZN(
        \DataP/alu_b_in[18] ) );
  OR2_X1 U1791 ( .A1(\DataP/alu_b_in[19] ), .A2(\DataP/alu_b_in[18] ), .ZN(
        n1737) );
  AND2_X1 U1792 ( .A1(n2075), .A2(n2027), .ZN(n1738) );
  NAND2_X1 U1793 ( .A1(n3488), .A2(n3489), .ZN(n1739) );
  BUF_X1 U1794 ( .A(n3588), .Z(n1740) );
  INV_X1 U1795 ( .A(n3539), .ZN(n1741) );
  INV_X1 U1796 ( .A(n3288), .ZN(n1742) );
  NAND2_X1 U1797 ( .A1(n2619), .A2(n1742), .ZN(n1743) );
  AND2_X1 U1798 ( .A1(\DataP/alu_a_in[0] ), .A2(n2226), .ZN(n3577) );
  NAND2_X1 U1799 ( .A1(n1633), .A2(n2726), .ZN(n1744) );
  AND2_X1 U1800 ( .A1(n2612), .A2(n3632), .ZN(n1745) );
  AND2_X1 U1801 ( .A1(n3648), .A2(\DataP/alu_a_in[19] ), .ZN(n1746) );
  OAI21_X1 U1802 ( .B1(n2044), .B2(n2128), .A(n2163), .ZN(n1747) );
  NOR2_X1 U1803 ( .A1(n3334), .A2(n3333), .ZN(n2206) );
  BUF_X1 U1804 ( .A(n3834), .Z(n1749) );
  INV_X1 U1805 ( .A(n1595), .ZN(\DataP/alu_b_in[2] ) );
  OR2_X4 U1806 ( .A1(n3365), .A2(n3364), .ZN(\DataP/alu_a_in[25] ) );
  AND4_X2 U1807 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n2082)
         );
  INV_X1 U1808 ( .A(\DataP/alu_a_in[17] ), .ZN(n1750) );
  BUF_X2 U1809 ( .A(\DataP/alu_a_in[17] ), .Z(n1751) );
  OAI21_X1 U1810 ( .B1(n3216), .B2(n2440), .A(n1840), .ZN(\DataP/alu_a_in[17] ) );
  INV_X1 U1811 ( .A(n3841), .ZN(n1752) );
  NAND4_X1 U1812 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(
        \DataP/alu_b_in[8] ) );
  AND4_X2 U1813 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n1753)
         );
  BUF_X1 U1814 ( .A(n3574), .Z(n1754) );
  AND3_X1 U1815 ( .A1(n1724), .A2(n2094), .A3(n1579), .ZN(n2092) );
  AND4_X2 U1816 ( .A1(n2176), .A2(n2178), .A3(n2621), .A4(n2175), .ZN(n2780)
         );
  NAND2_X1 U1817 ( .A1(n2615), .A2(n1756), .ZN(n3649) );
  AND2_X1 U1818 ( .A1(n2733), .A2(n2202), .ZN(n1756) );
  INV_X1 U1819 ( .A(\DataP/add_D[3] ), .ZN(n1757) );
  NAND4_X1 U1820 ( .A1(n3457), .A2(n3456), .A3(n3454), .A4(n3455), .ZN(
        \DataP/alu_b_in[11] ) );
  NAND2_X1 U1821 ( .A1(n2380), .A2(n1698), .ZN(n1758) );
  AOI21_X1 U1822 ( .B1(n1632), .B2(n2129), .A(n3795), .ZN(n1759) );
  OR2_X1 U1823 ( .A1(n2141), .A2(n1762), .ZN(n1761) );
  INV_X1 U1824 ( .A(n1573), .ZN(n1762) );
  NOR2_X1 U1825 ( .A1(n2371), .A2(n2108), .ZN(n2390) );
  NAND4_X1 U1826 ( .A1(n3325), .A2(n3326), .A3(n3324), .A4(n3323), .ZN(
        \DataP/alu_b_in[6] ) );
  OAI21_X1 U1827 ( .B1(n3624), .B2(\DataP/alu_b_in[15] ), .A(n2145), .ZN(n2329) );
  INV_X1 U1828 ( .A(n2068), .ZN(n2043) );
  NOR2_X1 U1829 ( .A1(n1761), .A2(n2145), .ZN(n2675) );
  AOI211_X1 U1830 ( .C1(n2279), .C2(n2278), .A(n2277), .B(n2348), .ZN(n2291)
         );
  NOR2_X1 U1831 ( .A1(n2379), .A2(n2395), .ZN(n2033) );
  AND3_X2 U1832 ( .A1(n3531), .A2(n3530), .A3(n1963), .ZN(n2371) );
  NOR2_X1 U1833 ( .A1(n2068), .A2(\lt_x_135/B[12] ), .ZN(n2042) );
  XNOR2_X1 U1834 ( .A(n3620), .B(n2145), .ZN(n2685) );
  NAND2_X1 U1835 ( .A1(n1647), .A2(n2041), .ZN(n3620) );
  NOR2_X1 U1836 ( .A1(n2068), .A2(n1761), .ZN(n2041) );
  INV_X1 U1837 ( .A(n2108), .ZN(n2128) );
  INV_X1 U1838 ( .A(n2016), .ZN(n2014) );
  OR2_X2 U1839 ( .A1(n3340), .A2(n3339), .ZN(\DataP/alu_a_in[5] ) );
  OR2_X2 U1840 ( .A1(n3398), .A2(n3397), .ZN(\DataP/alu_a_in[12] ) );
  BUF_X1 U1841 ( .A(n1734), .Z(n2167) );
  NAND2_X1 U1842 ( .A1(n2040), .A2(n1968), .ZN(n3608) );
  NAND2_X1 U1843 ( .A1(n2680), .A2(n3886), .ZN(n2039) );
  INV_X1 U1844 ( .A(n2052), .ZN(n2048) );
  BUF_X1 U1845 ( .A(n3606), .Z(n2156) );
  INV_X1 U1846 ( .A(\DataP/a_out[27] ), .ZN(n1977) );
  INV_X1 U1847 ( .A(\DataP/a_out[29] ), .ZN(n1978) );
  INV_X1 U1848 ( .A(\DataP/a_out[26] ), .ZN(n1979) );
  INV_X1 U1849 ( .A(\DataP/a_out[28] ), .ZN(n1980) );
  INV_X1 U1850 ( .A(\DataP/a_out[1] ), .ZN(n1981) );
  INV_X1 U1851 ( .A(\DataP/a_out[7] ), .ZN(n1982) );
  INV_X1 U1852 ( .A(\DataP/a_out[10] ), .ZN(n1983) );
  INV_X1 U1853 ( .A(\DataP/a_out[11] ), .ZN(n1984) );
  INV_X1 U1854 ( .A(\DataP/a_out[12] ), .ZN(n1985) );
  INV_X1 U1855 ( .A(\DataP/a_out[13] ), .ZN(n1986) );
  INV_X1 U1856 ( .A(\DataP/a_out[14] ), .ZN(n1987) );
  INV_X1 U1857 ( .A(\DataP/a_out[15] ), .ZN(n1988) );
  INV_X1 U1858 ( .A(\DataP/a_out[30] ), .ZN(n2001) );
  INV_X1 U1859 ( .A(\DataP/a_out[3] ), .ZN(n2002) );
  INV_X1 U1860 ( .A(\DataP/a_out[4] ), .ZN(n2003) );
  INV_X1 U1861 ( .A(\DataP/a_out[5] ), .ZN(n2004) );
  INV_X1 U1862 ( .A(\DataP/a_out[6] ), .ZN(n2005) );
  INV_X1 U1863 ( .A(\CU_I/cw[10] ), .ZN(n2007) );
  NAND2_X1 U1864 ( .A1(n2063), .A2(n2065), .ZN(n2560) );
  NAND2_X1 U1865 ( .A1(n3777), .A2(n2066), .ZN(n2065) );
  NAND3_X1 U1866 ( .A1(n2034), .A2(n3432), .A3(n2290), .ZN(n1763) );
  OAI211_X1 U1867 ( .C1(n3562), .C2(n2391), .A(n2016), .B(n1763), .ZN(n2013)
         );
  AOI22_X1 U1868 ( .A1(n3051), .A2(n2856), .B1(n2919), .B2(n2879), .ZN(n1764)
         );
  AOI22_X1 U1869 ( .A1(n2115), .A2(n2857), .B1(n2101), .B2(n1764), .ZN(n1765)
         );
  MUX2_X1 U1870 ( .A(n1765), .B(n2901), .S(n2138), .Z(
        \DataP/ALU_C/shifter/N43 ) );
  INV_X1 U1871 ( .A(\DataP/a_out[16] ), .ZN(n1989) );
  NOR2_X1 U1872 ( .A1(n3055), .A2(n2902), .ZN(n1766) );
  OAI21_X1 U1873 ( .B1(n3897), .B2(n3495), .A(n3453), .ZN(n1767) );
  NOR2_X1 U1874 ( .A1(n3450), .A2(n3489), .ZN(n1768) );
  XNOR2_X1 U1875 ( .A(n1768), .B(n3458), .ZN(n1769) );
  OAI221_X1 U1876 ( .B1(n2102), .B2(n3132), .C1(n1866), .C2(n3071), .A(n3877), 
        .ZN(n1770) );
  INV_X1 U1877 ( .A(n3055), .ZN(n1771) );
  OAI221_X1 U1878 ( .B1(n3055), .B2(n2935), .C1(n1771), .C2(n2995), .A(n3227), 
        .ZN(n1772) );
  OAI211_X1 U1879 ( .C1(n3880), .C2(n1769), .A(n1770), .B(n1772), .ZN(n1773)
         );
  AOI211_X1 U1880 ( .C1(n3228), .C2(n1766), .A(n1767), .B(n1773), .ZN(n340) );
  AOI211_X1 U1881 ( .C1(n2301), .C2(\DataP/alu_a_in[16] ), .A(n2298), .B(n2274), .ZN(n1774) );
  AOI221_X1 U1882 ( .B1(n2320), .B2(n2257), .C1(n2256), .C2(n2257), .A(n2255), 
        .ZN(n1775) );
  AOI211_X1 U1883 ( .C1(n2266), .C2(n2267), .A(n2264), .B(n2265), .ZN(n1776)
         );
  OAI21_X1 U1884 ( .B1(n1775), .B2(n2268), .A(n1776), .ZN(n1777) );
  NAND3_X1 U1885 ( .A1(n2369), .A2(n1774), .A3(n1777), .ZN(n2292) );
  AOI22_X1 U1886 ( .A1(n3224), .A2(\DataP/alu_out_W[30] ), .B1(\DataP/B_s[30] ), .B2(n2227), .ZN(n1778) );
  OAI211_X1 U1887 ( .C1(n2417), .C2(n2772), .A(n3523), .B(n1778), .ZN(
        \DataP/alu_b_in[30] ) );
  OAI21_X1 U1888 ( .B1(n2135), .B2(n3851), .A(n3891), .ZN(n1779) );
  AOI22_X1 U1889 ( .A1(\DataP/alu_a_in[18] ), .A2(n3894), .B1(n1736), .B2(
        n1779), .ZN(n1780) );
  NAND3_X1 U1890 ( .A1(n3227), .A2(n3006), .A3(n2102), .ZN(n1781) );
  OAI211_X1 U1891 ( .C1(n3897), .C2(n3747), .A(n1780), .B(n1781), .ZN(n3748)
         );
  AOI22_X1 U1892 ( .A1(n3052), .A2(n3033), .B1(n3034), .B2(n3051), .ZN(n1782)
         );
  AOI22_X1 U1893 ( .A1(n1782), .A2(n2101), .B1(n3035), .B2(n2112), .ZN(n3037)
         );
  INV_X1 U1894 ( .A(\DataP/a_out[17] ), .ZN(n1990) );
  OAI21_X1 U1895 ( .B1(n2102), .B2(n3198), .A(n3194), .ZN(n1783) );
  AOI21_X1 U1896 ( .B1(n2221), .B2(n3837), .A(n3428), .ZN(n1784) );
  NAND2_X1 U1897 ( .A1(n3443), .A2(n3483), .ZN(n1785) );
  NOR2_X1 U1898 ( .A1(n1784), .A2(n1785), .ZN(n1786) );
  AOI211_X1 U1899 ( .C1(n1784), .C2(n1785), .A(n3880), .B(n1786), .ZN(n1787)
         );
  NOR2_X1 U1900 ( .A1(n3055), .A2(n2915), .ZN(n1788) );
  AOI22_X1 U1901 ( .A1(\DataP/ALU_C/shifter/N59 ), .A2(n3227), .B1(n3228), 
        .B2(n1788), .ZN(n1789) );
  OAI211_X1 U1902 ( .C1(n3897), .C2(n3494), .A(n3437), .B(n1789), .ZN(n1790)
         );
  AOI211_X1 U1903 ( .C1(n3877), .C2(n1783), .A(n1787), .B(n1790), .ZN(n341) );
  NAND2_X1 U1904 ( .A1(n3569), .A2(ALU_OPCODE_i[0]), .ZN(n1791) );
  AOI21_X1 U1905 ( .B1(n2034), .B2(n2290), .A(n1791), .ZN(n1792) );
  NOR3_X1 U1906 ( .A1(n1792), .A2(n1964), .A3(n2033), .ZN(n2032) );
  INV_X1 U1907 ( .A(\DataP/a_out[18] ), .ZN(n1991) );
  OAI21_X1 U1908 ( .B1(n3206), .B2(n3197), .A(n3190), .ZN(n1793) );
  OAI22_X1 U1909 ( .A1(n3841), .A2(n3842), .B1(n2110), .B2(n3840), .ZN(n1794)
         );
  INV_X1 U1910 ( .A(n3055), .ZN(n1795) );
  OAI221_X1 U1911 ( .B1(n3055), .B2(n3041), .C1(n1795), .C2(n3040), .A(n3900), 
        .ZN(n1796) );
  NOR2_X1 U1912 ( .A1(n2138), .A2(n2914), .ZN(n1797) );
  XNOR2_X1 U1913 ( .A(\DataP/alu_a_in[8] ), .B(n2204), .ZN(n1798) );
  AOI21_X1 U1914 ( .B1(n3835), .B2(n2221), .A(n3837), .ZN(n1799) );
  AOI211_X1 U1915 ( .C1(n3837), .C2(n1798), .A(n1799), .B(n3880), .ZN(n1800)
         );
  AOI21_X1 U1916 ( .B1(n3228), .B2(n1797), .A(n1800), .ZN(n1801) );
  NAND2_X1 U1917 ( .A1(n1796), .A2(n1801), .ZN(n1802) );
  AOI211_X1 U1918 ( .C1(n3877), .C2(n1793), .A(n1794), .B(n1802), .ZN(n345) );
  AOI22_X1 U1919 ( .A1(n3697), .A2(\DataP/alu_b_in[27] ), .B1(n2354), .B2(
        \DataP/alu_b_in[26] ), .ZN(n1803) );
  INV_X1 U1920 ( .A(n2355), .ZN(n1804) );
  AOI221_X1 U1921 ( .B1(n2356), .B2(n1803), .C1(n2367), .C2(n1803), .A(n1804), 
        .ZN(n2359) );
  OAI21_X1 U1922 ( .B1(\DataP/alu_a_in[16] ), .B2(\DataP/alu_b_in[16] ), .A(
        n3894), .ZN(n1805) );
  NAND3_X1 U1923 ( .A1(\DataP/alu_a_in[16] ), .A2(\DataP/alu_b_in[16] ), .A3(
        n3890), .ZN(n1806) );
  OAI211_X1 U1924 ( .C1(n3731), .C2(n3897), .A(n1805), .B(n1806), .ZN(n3732)
         );
  AOI22_X1 U1925 ( .A1(n3189), .A2(n3205), .B1(n2101), .B2(n3188), .ZN(n1807)
         );
  NAND2_X1 U1926 ( .A1(n3206), .A2(n1807), .ZN(n3190) );
  INV_X1 U1927 ( .A(\DataP/a_out[19] ), .ZN(n1992) );
  XOR2_X1 U1928 ( .A(n3854), .B(n2203), .Z(n1808) );
  INV_X1 U1929 ( .A(n3055), .ZN(n1809) );
  OAI221_X1 U1930 ( .B1(n3055), .B2(n3032), .C1(n1809), .C2(n3031), .A(n3900), 
        .ZN(n1810) );
  OAI21_X1 U1931 ( .B1(n2102), .B2(n3181), .A(n3180), .ZN(n1811) );
  NAND2_X1 U1932 ( .A1(n1811), .A2(n3877), .ZN(n1812) );
  OAI211_X1 U1933 ( .C1(n1808), .C2(n3880), .A(n1810), .B(n1812), .ZN(n1813)
         );
  AOI21_X1 U1934 ( .B1(n3894), .B2(\DataP/alu_a_in[6] ), .A(n3858), .ZN(n1814)
         );
  NAND3_X1 U1935 ( .A1(n3228), .A2(n2898), .A3(n1809), .ZN(n1815) );
  OAI211_X1 U1936 ( .C1(n3897), .C2(n3859), .A(n1814), .B(n1815), .ZN(n1816)
         );
  NOR2_X1 U1937 ( .A1(n1813), .A2(n1816), .ZN(n353) );
  NOR2_X1 U1938 ( .A1(\DataP/alu_a_in[18] ), .A2(n2341), .ZN(n1817) );
  AOI22_X1 U1939 ( .A1(n1722), .A2(n2202), .B1(n1736), .B2(n1817), .ZN(n2346)
         );
  NAND3_X1 U1940 ( .A1(n1574), .A2(n2120), .A3(n3726), .ZN(n1818) );
  NAND2_X1 U1941 ( .A1(n1818), .A2(n1694), .ZN(n1819) );
  XNOR2_X1 U1942 ( .A(n1819), .B(n2125), .ZN(n3728) );
  OAI211_X1 U1943 ( .C1(n3800), .C2(n3897), .A(n1820), .B(n1821), .ZN(n3801)
         );
  INV_X1 U1944 ( .A(\DataP/a_out[20] ), .ZN(n1993) );
  NOR2_X1 U1945 ( .A1(n3055), .A2(n2912), .ZN(n1822) );
  NAND2_X1 U1946 ( .A1(n2215), .A2(n2156), .ZN(n1823) );
  XNOR2_X1 U1947 ( .A(n1823), .B(n3607), .ZN(n1824) );
  OAI21_X1 U1948 ( .B1(n3206), .B2(n3174), .A(n3173), .ZN(n1825) );
  NAND2_X1 U1949 ( .A1(n1825), .A2(n3877), .ZN(n1826) );
  OAI21_X1 U1950 ( .B1(n3880), .B2(n1824), .A(n1826), .ZN(n1827) );
  OAI221_X1 U1951 ( .B1(n2138), .B2(n3026), .C1(n1908), .C2(n3025), .A(n3227), 
        .ZN(n1828) );
  OAI211_X1 U1952 ( .C1(n3603), .C2(n3897), .A(n3602), .B(n1828), .ZN(n1829)
         );
  AOI211_X1 U1953 ( .C1(n3228), .C2(n1822), .A(n1827), .B(n1829), .ZN(n354) );
  NAND2_X1 U1954 ( .A1(n1694), .A2(n2031), .ZN(n1830) );
  XNOR2_X1 U1955 ( .A(n1830), .B(n2030), .ZN(n3427) );
  AOI22_X1 U1956 ( .A1(\DataP/alu_out_W[27] ), .A2(n3207), .B1(
        \DataP/alu_out_M[27] ), .B2(n3211), .ZN(n1831) );
  OAI21_X1 U1957 ( .B1(n3213), .B2(n145), .A(n1831), .ZN(n1832) );
  NOR2_X1 U1958 ( .A1(n3217), .A2(n2438), .ZN(n1833) );
  NOR2_X2 U1959 ( .A1(n1832), .A2(n1833), .ZN(n3697) );
  AOI22_X1 U1960 ( .A1(n3219), .A2(\DataP/B_s[22] ), .B1(n1581), .B2(
        \DataP/IMM_s[22] ), .ZN(n1834) );
  NAND2_X1 U1961 ( .A1(n3224), .A2(\DataP/alu_out_W[22] ), .ZN(n1835) );
  OAI211_X1 U1962 ( .C1(n2428), .C2(n2772), .A(n1834), .B(n1835), .ZN(
        \DataP/alu_b_in[22] ) );
  AOI21_X1 U1963 ( .B1(n3890), .B2(n3048), .A(n3894), .ZN(n1836) );
  OAI22_X1 U1964 ( .A1(n3891), .A2(n3047), .B1(n1715), .B2(n1836), .ZN(n3578)
         );
  INV_X1 U1965 ( .A(\DataP/a_out[21] ), .ZN(n1994) );
  OAI21_X1 U1966 ( .B1(\DataP/alu_b_in[15] ), .B2(n2210), .A(n2145), .ZN(n1837) );
  OAI22_X1 U1967 ( .A1(\DataP/alu_a_in[14] ), .A2(n1837), .B1(
        \DataP/alu_a_in[15] ), .B2(n2230), .ZN(n2264) );
  INV_X1 U1968 ( .A(n1725), .ZN(n1838) );
  INV_X1 U1969 ( .A(n3214), .ZN(n1839) );
  AOI222_X1 U1970 ( .A1(n1606), .A2(n1839), .B1(\DataP/alu_out_M[17] ), .B2(
        n2209), .C1(n3207), .C2(\DataP/alu_out_W[17] ), .ZN(n1840) );
  AOI22_X1 U1971 ( .A1(n3219), .A2(\DataP/B_s[24] ), .B1(n1581), .B2(
        \DataP/IMM_s[24] ), .ZN(n1841) );
  NAND2_X1 U1972 ( .A1(n3226), .A2(\DataP/alu_out_W[24] ), .ZN(n1842) );
  NAND2_X1 U1973 ( .A1(n2026), .A2(n1694), .ZN(n1843) );
  XNOR2_X1 U1974 ( .A(n3429), .B(n1843), .ZN(n2011) );
  INV_X1 U1975 ( .A(\DataP/a_out[22] ), .ZN(n1995) );
  NOR2_X1 U1976 ( .A1(n2138), .A2(n2911), .ZN(n1844) );
  XNOR2_X1 U1977 ( .A(\DataP/alu_a_in[4] ), .B(n3849), .ZN(n1845) );
  XNOR2_X1 U1978 ( .A(n1845), .B(n3850), .ZN(n1846) );
  OAI21_X1 U1979 ( .B1(n2102), .B2(n3167), .A(n3166), .ZN(n1847) );
  NAND2_X1 U1980 ( .A1(n1847), .A2(n3877), .ZN(n1848) );
  OAI21_X1 U1981 ( .B1(n3880), .B2(n1846), .A(n1848), .ZN(n1849) );
  AOI22_X1 U1982 ( .A1(n2138), .A2(n3894), .B1(\DataP/alu_a_in[4] ), .B2(n3852), .ZN(n1850) );
  INV_X1 U1983 ( .A(n3055), .ZN(n1851) );
  OAI221_X1 U1984 ( .B1(n3055), .B2(n3020), .C1(n1851), .C2(n3019), .A(n3900), 
        .ZN(n1852) );
  OAI211_X1 U1985 ( .C1(n3853), .C2(n3897), .A(n1850), .B(n1852), .ZN(n1853)
         );
  AOI211_X1 U1986 ( .C1(n3228), .C2(n1844), .A(n1849), .B(n1853), .ZN(n355) );
  AND3_X1 U1987 ( .A1(n2123), .A2(n1722), .A3(n2108), .ZN(n2617) );
  NAND3_X1 U1988 ( .A1(n1647), .A2(n2043), .A3(n2675), .ZN(n1854) );
  XNOR2_X1 U1989 ( .A(n1854), .B(n2230), .ZN(n3616) );
  INV_X1 U1990 ( .A(n2535), .ZN(n1855) );
  NAND2_X1 U1991 ( .A1(n2213), .A2(n1855), .ZN(n1856) );
  XNOR2_X1 U1992 ( .A(\DataP/alu_b_in[20] ), .B(n1856), .ZN(n3666) );
  AOI22_X1 U1993 ( .A1(n3225), .A2(\DataP/alu_out_W[29] ), .B1(n2782), .B2(
        \DataP/alu_out_M[29] ), .ZN(n1857) );
  NAND2_X1 U1994 ( .A1(\DataP/B_s[29] ), .A2(n2227), .ZN(n1858) );
  NAND3_X1 U1995 ( .A1(n1858), .A2(n1857), .A3(n3523), .ZN(
        \DataP/alu_b_in[29] ) );
  OAI21_X1 U1996 ( .B1(n2074), .B2(n3851), .A(n3891), .ZN(n1859) );
  AOI22_X1 U1997 ( .A1(\lt_x_135/B[5] ), .A2(n3894), .B1(\DataP/alu_a_in[5] ), 
        .B2(n1859), .ZN(n3602) );
  INV_X1 U1998 ( .A(\DataP/a_out[23] ), .ZN(n1996) );
  OAI211_X1 U1999 ( .C1(n3872), .C2(n3897), .A(n3871), .B(n3870), .ZN(n1860)
         );
  NOR2_X1 U2000 ( .A1(n3055), .A2(n2905), .ZN(n1861) );
  AOI21_X1 U2001 ( .B1(n1861), .B2(n3228), .A(n1860), .ZN(n1862) );
  NOR2_X1 U2002 ( .A1(n3861), .A2(n3862), .ZN(n1863) );
  OAI211_X1 U2003 ( .C1(n3868), .C2(n3867), .A(n3866), .B(n2208), .ZN(n1864)
         );
  OAI211_X1 U2004 ( .C1(n1863), .C2(n2214), .A(n2129), .B(n1864), .ZN(n1865)
         );
  INV_X1 U2005 ( .A(n2102), .ZN(n1866) );
  OAI221_X1 U2006 ( .B1(n2102), .B2(n3138), .C1(n1866), .C2(n3088), .A(n3877), 
        .ZN(n1867) );
  OAI221_X1 U2007 ( .B1(n2138), .B2(n2953), .C1(n1888), .C2(n2998), .A(n3227), 
        .ZN(n1868) );
  AND4_X1 U2008 ( .A1(n1862), .A2(n1865), .A3(n1867), .A4(n1868), .ZN(n333) );
  AOI22_X1 U2009 ( .A1(n3211), .A2(\DataP/alu_out_M[19] ), .B1(
        \DataP/alu_out_W[19] ), .B2(n3207), .ZN(n1869) );
  OAI21_X1 U2010 ( .B1(n113), .B2(n3213), .A(n1869), .ZN(n3382) );
  AOI22_X1 U2011 ( .A1(n2103), .A2(\DataP/alu_a_in[30] ), .B1(
        \DataP/alu_a_in[31] ), .B2(n2916), .ZN(n1870) );
  AOI22_X1 U2012 ( .A1(n2105), .A2(n1870), .B1(n2891), .B2(n2917), .ZN(n1871)
         );
  AOI22_X1 U2013 ( .A1(n3202), .A2(n2892), .B1(n1871), .B2(n3053), .ZN(n1872)
         );
  AOI22_X1 U2014 ( .A1(n2115), .A2(n2893), .B1(n2101), .B2(n1872), .ZN(n1873)
         );
  MUX2_X1 U2015 ( .A(n1873), .B(n2894), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N49 ) );
  INV_X1 U2016 ( .A(n3055), .ZN(n1874) );
  NAND3_X1 U2017 ( .A1(n3904), .A2(n2810), .A3(n1874), .ZN(n3558) );
  AOI22_X1 U2018 ( .A1(n3225), .A2(\DataP/alu_out_W[28] ), .B1(\DataP/B_s[28] ), .B2(n2227), .ZN(n1875) );
  OAI211_X1 U2019 ( .C1(n2426), .C2(n1627), .A(n3523), .B(n1875), .ZN(
        \DataP/alu_b_in[28] ) );
  AOI22_X1 U2020 ( .A1(n3052), .A2(n3016), .B1(n3017), .B2(n3202), .ZN(n1876)
         );
  AOI22_X1 U2021 ( .A1(n1876), .A2(n2101), .B1(n3018), .B2(n2112), .ZN(n3020)
         );
  NAND3_X1 U2022 ( .A1(\DataP/alu_a_in[14] ), .A2(n2145), .A3(n3890), .ZN(
        n1877) );
  OAI21_X1 U2023 ( .B1(\DataP/alu_a_in[14] ), .B2(n2145), .A(n3894), .ZN(n1878) );
  OAI211_X1 U2024 ( .C1(n3875), .C2(n3897), .A(n1877), .B(n1878), .ZN(n3876)
         );
  INV_X1 U2025 ( .A(\DataP/a_out[24] ), .ZN(n1997) );
  OAI21_X1 U2026 ( .B1(n2102), .B2(n3160), .A(n3159), .ZN(n1879) );
  INV_X1 U2027 ( .A(n3228), .ZN(n1880) );
  NOR3_X1 U2028 ( .A1(n3055), .A2(n2910), .A3(n1880), .ZN(n1881) );
  AOI22_X1 U2029 ( .A1(n1973), .A2(n3846), .B1(\DataP/alu_b_in[3] ), .B2(n3894), .ZN(n1882) );
  OAI211_X1 U2030 ( .C1(n3897), .C2(n3848), .A(n3847), .B(n1882), .ZN(n1883)
         );
  AOI211_X1 U2031 ( .C1(n3877), .C2(n1879), .A(n1881), .B(n1883), .ZN(n1884)
         );
  AOI22_X1 U2032 ( .A1(n3049), .A2(n3013), .B1(n3047), .B2(n3012), .ZN(n1885)
         );
  AOI22_X1 U2033 ( .A1(n3202), .A2(n3033), .B1(n3052), .B2(n1885), .ZN(n1886)
         );
  AOI22_X1 U2034 ( .A1(n2101), .A2(n1886), .B1(n3014), .B2(n3204), .ZN(n1887)
         );
  INV_X1 U2035 ( .A(n3055), .ZN(n1888) );
  OAI221_X1 U2036 ( .B1(n3055), .B2(n1887), .C1(n1888), .C2(n3015), .A(n3227), 
        .ZN(n1889) );
  AND2_X1 U2037 ( .A1(n1884), .A2(n1889), .ZN(n356) );
  NAND2_X1 U2038 ( .A1(n2208), .A2(n3863), .ZN(n1890) );
  XOR2_X1 U2039 ( .A(n1710), .B(n1890), .Z(n1891) );
  OAI21_X1 U2040 ( .B1(n3206), .B2(n2997), .A(n2942), .ZN(n1892) );
  OAI211_X1 U2041 ( .C1(n3496), .C2(n3897), .A(n3493), .B(n3492), .ZN(n1893)
         );
  AOI21_X1 U2042 ( .B1(n3227), .B2(n1892), .A(n1893), .ZN(n1894) );
  OAI221_X1 U2043 ( .B1(n2102), .B2(n3136), .C1(n1866), .C2(n3078), .A(n3877), 
        .ZN(n1895) );
  OAI211_X1 U2044 ( .C1(n3880), .C2(n1891), .A(n1894), .B(n1895), .ZN(n1896)
         );
  NOR2_X1 U2045 ( .A1(n3055), .A2(n2904), .ZN(n1897) );
  AOI21_X1 U2046 ( .B1(n1897), .B2(n3228), .A(n1896), .ZN(n337) );
  INV_X1 U2047 ( .A(n2381), .ZN(n1898) );
  NAND2_X1 U2048 ( .A1(n2614), .A2(n1898), .ZN(n2385) );
  INV_X1 U2049 ( .A(n2209), .ZN(n1899) );
  OAI222_X1 U2050 ( .A1(n2433), .A2(n1899), .B1(n3213), .B2(n97), .C1(n2072), 
        .C2(n2516), .ZN(n2693) );
  AOI22_X1 U2051 ( .A1(n1631), .A2(\DataP/B_s[18] ), .B1(n1623), .B2(
        \DataP/IMM_s[18] ), .ZN(n1900) );
  NAND2_X1 U2052 ( .A1(n3225), .A2(\DataP/alu_out_W[18] ), .ZN(n1901) );
  OAI211_X1 U2053 ( .C1(n2772), .C2(n2478), .A(n2661), .B(n2662), .ZN(n1902)
         );
  INV_X1 U2054 ( .A(n1902), .ZN(n2660) );
  NAND2_X1 U2055 ( .A1(n1597), .A2(n2108), .ZN(n1903) );
  NAND3_X1 U2056 ( .A1(n1903), .A2(\DataP/alu_a_in[12] ), .A3(n2739), .ZN(
        n3865) );
  NOR2_X1 U2057 ( .A1(n2744), .A2(n3826), .ZN(n1904) );
  INV_X1 U2058 ( .A(n4183), .ZN(n1905) );
  AOI221_X1 U2059 ( .B1(n4184), .B2(n4183), .C1(n3907), .C2(n1905), .A(n4182), 
        .ZN(\DataP/wrong_br ) );
  OAI21_X1 U2060 ( .B1(n1613), .B2(n2067), .A(n2064), .ZN(n1906) );
  INV_X1 U2061 ( .A(n1906), .ZN(n2063) );
  AOI22_X1 U2062 ( .A1(n2101), .A2(n2857), .B1(n2858), .B2(n2115), .ZN(n1907)
         );
  INV_X1 U2063 ( .A(n3055), .ZN(n1908) );
  OAI221_X1 U2064 ( .B1(n3055), .B2(n1907), .C1(n1908), .C2(n2827), .A(n3228), 
        .ZN(n3743) );
  INV_X1 U2065 ( .A(\DataP/a_out[25] ), .ZN(n1998) );
  NOR2_X1 U2066 ( .A1(n3055), .A2(n2913), .ZN(n1909) );
  OAI21_X1 U2067 ( .B1(n3854), .B2(n3610), .A(n1648), .ZN(n1910) );
  OAI21_X1 U2068 ( .B1(n2102), .B2(n3196), .A(n3187), .ZN(n1911) );
  NAND2_X1 U2069 ( .A1(n1911), .A2(n3877), .ZN(n1912) );
  XOR2_X1 U2070 ( .A(n1910), .B(n2211), .Z(n1913) );
  OAI21_X1 U2071 ( .B1(n1913), .B2(n3880), .A(n1912), .ZN(n1914) );
  AOI22_X1 U2072 ( .A1(\DataP/alu_a_in[7] ), .A2(n3894), .B1(
        \DataP/alu_b_in[7] ), .B2(n3612), .ZN(n1915) );
  INV_X1 U2073 ( .A(n3055), .ZN(n1916) );
  OAI221_X1 U2074 ( .B1(n3055), .B2(n3037), .C1(n1916), .C2(n3036), .A(n3227), 
        .ZN(n1917) );
  OAI211_X1 U2075 ( .C1(n3897), .C2(n3613), .A(n1915), .B(n1917), .ZN(n1918)
         );
  NOR2_X1 U2076 ( .A1(n2119), .A2(n1973), .ZN(n1919) );
  NAND3_X1 U2077 ( .A1(n2254), .A2(n2080), .A3(n2081), .ZN(n1920) );
  OAI21_X1 U2078 ( .B1(\DataP/alu_a_in[2] ), .B2(n2315), .A(n1920), .ZN(n1921)
         );
  OAI22_X1 U2079 ( .A1(n1919), .A2(n1921), .B1(\lt_x_135/B[5] ), .B2(n2113), 
        .ZN(n1922) );
  NAND2_X1 U2080 ( .A1(\DataP/alu_a_in[26] ), .A2(n2127), .ZN(n1923) );
  OAI21_X1 U2081 ( .B1(n3697), .B2(\DataP/alu_b_in[27] ), .A(n1923), .ZN(n2297) );
  NAND4_X1 U2082 ( .A1(n4108), .A2(n3782), .A3(n3771), .A4(n4109), .ZN(n2743)
         );
  INV_X1 U2083 ( .A(\DataP/alu_a_in[25] ), .ZN(n1924) );
  AOI21_X1 U2084 ( .B1(n2586), .B2(n2585), .A(n1924), .ZN(n3798) );
  INV_X1 U2085 ( .A(n2108), .ZN(n1925) );
  NOR2_X1 U2086 ( .A1(n1925), .A2(n3416), .ZN(n1926) );
  AOI21_X1 U2087 ( .B1(n2128), .B2(n2739), .A(\DataP/alu_a_in[12] ), .ZN(n2735) );
  INV_X1 U2088 ( .A(n2241), .ZN(n1927) );
  NOR2_X1 U2089 ( .A1(n3725), .A2(n1927), .ZN(n2432) );
  AOI22_X1 U2090 ( .A1(n1631), .A2(\DataP/B_s[19] ), .B1(n1623), .B2(
        \DataP/IMM_s[19] ), .ZN(n1928) );
  NAND2_X1 U2091 ( .A1(n3226), .A2(\DataP/alu_out_W[19] ), .ZN(n1929) );
  INV_X1 U2092 ( .A(n3680), .ZN(n1930) );
  AOI21_X1 U2093 ( .B1(n2378), .B2(n1930), .A(n1707), .ZN(n2674) );
  INV_X1 U2094 ( .A(n3688), .ZN(n1931) );
  NOR2_X1 U2095 ( .A1(n1931), .A2(n2133), .ZN(n1932) );
  AOI22_X1 U2096 ( .A1(n1931), .A2(n2133), .B1(n3672), .B2(n1932), .ZN(n2064)
         );
  AOI21_X1 U2097 ( .B1(n2102), .B2(n3150), .A(n3195), .ZN(n1933) );
  OAI211_X1 U2098 ( .C1(n3707), .C2(n3897), .A(n3706), .B(n3705), .ZN(n1934)
         );
  AOI21_X1 U2099 ( .B1(n3227), .B2(\DataP/ALU_C/shifter/N80 ), .A(n1934), .ZN(
        n1935) );
  AOI22_X1 U2100 ( .A1(n3202), .A2(n2888), .B1(n2918), .B2(n2887), .ZN(n1936)
         );
  AOI22_X1 U2101 ( .A1(n2115), .A2(n2889), .B1(n2101), .B2(n1936), .ZN(n1937)
         );
  OAI221_X1 U2102 ( .B1(n2138), .B2(n1937), .C1(n1916), .C2(n2890), .A(n3904), 
        .ZN(n1938) );
  OAI211_X1 U2103 ( .C1(n3892), .C2(n1933), .A(n1935), .B(n1938), .ZN(n2756)
         );
  INV_X1 U2104 ( .A(\DataP/a_out[0] ), .ZN(n1999) );
  NOR2_X1 U2105 ( .A1(n3788), .A2(n2744), .ZN(n2389) );
  AOI22_X1 U2106 ( .A1(n3210), .A2(DRAM_ADDRESS[9]), .B1(n3207), .B2(
        \DataP/alu_out_W[9] ), .ZN(n1939) );
  NAND2_X1 U2107 ( .A1(n2139), .A2(\DataP/npc_E[9] ), .ZN(n1940) );
  OAI211_X1 U2108 ( .C1(n3216), .C2(n2435), .A(n1939), .B(n1940), .ZN(
        \DataP/alu_a_in[9] ) );
  XOR2_X1 U2109 ( .A(\lt_x_135/B[12] ), .B(n1941), .Z(n3481) );
  OAI211_X1 U2110 ( .C1(n2685), .C2(n2128), .A(n2651), .B(n2652), .ZN(n3631)
         );
  OAI221_X1 U2111 ( .B1(n3195), .B2(n3101), .C1(n3195), .C2(n2102), .A(n3877), 
        .ZN(n3734) );
  AOI22_X1 U2112 ( .A1(n3051), .A2(n2861), .B1(n2918), .B2(n2888), .ZN(n1942)
         );
  AOI22_X1 U2113 ( .A1(n2101), .A2(n1942), .B1(n2862), .B2(n2115), .ZN(n1943)
         );
  INV_X1 U2114 ( .A(n3055), .ZN(n1944) );
  OAI221_X1 U2115 ( .B1(n3055), .B2(n1943), .C1(n1944), .C2(n2863), .A(n3228), 
        .ZN(n3814) );
  INV_X1 U2116 ( .A(n3417), .ZN(n1945) );
  NAND2_X1 U2117 ( .A1(\DataP/alu_a_in[2] ), .A2(n1945), .ZN(n3585) );
  NOR3_X1 U2118 ( .A1(n4005), .A2(IR_CU[4]), .A3(IR_CU[5]), .ZN(n1946) );
  AOI21_X1 U2119 ( .B1(n3996), .B2(n607), .A(n1946), .ZN(n1947) );
  OAI221_X1 U2120 ( .B1(n4036), .B2(n4027), .C1(n4036), .C2(n4016), .A(n1947), 
        .ZN(n4006) );
  AOI21_X1 U2121 ( .B1(n2432), .B2(n2766), .A(n2765), .ZN(n1948) );
  NOR2_X1 U2122 ( .A1(n2746), .A2(n1948), .ZN(n2719) );
  OAI21_X1 U2123 ( .B1(n2234), .B2(n2673), .A(n2674), .ZN(n1949) );
  OAI21_X1 U2124 ( .B1(n3682), .B2(n1949), .A(n2167), .ZN(n3650) );
  INV_X1 U2125 ( .A(\DataP/a_out[31] ), .ZN(n2006) );
  NAND2_X1 U2126 ( .A1(n3964), .A2(n3965), .ZN(n1950) );
  NOR3_X1 U2127 ( .A1(n3969), .A2(n3970), .A3(n3971), .ZN(n1951) );
  NAND4_X1 U2128 ( .A1(n3972), .A2(n3973), .A3(n3968), .A4(n1951), .ZN(n1952)
         );
  NOR4_X1 U2129 ( .A1(n3966), .A2(n3967), .A3(n1950), .A4(n1952), .ZN(n1953)
         );
  INV_X1 U2130 ( .A(n3956), .ZN(n1954) );
  NAND4_X1 U2131 ( .A1(n3957), .A2(n3958), .A3(n3959), .A4(n1954), .ZN(n1955)
         );
  NOR2_X1 U2132 ( .A1(n3954), .A2(n3955), .ZN(n1956) );
  NAND3_X1 U2133 ( .A1(n3953), .A2(n3952), .A3(n1956), .ZN(n1957) );
  NOR4_X1 U2134 ( .A1(n3960), .A2(n3961), .A3(n1955), .A4(n1957), .ZN(n1958)
         );
  NAND4_X1 U2135 ( .A1(n3962), .A2(n3963), .A3(n1953), .A4(n1958), .ZN(n1959)
         );
  NAND2_X1 U2136 ( .A1(n3974), .A2(n1959), .ZN(\DataP/NPC_add/N0 ) );
  INV_X1 U2137 ( .A(n2108), .ZN(n2535) );
  INV_X2 U2138 ( .A(n3051), .ZN(n2919) );
  INV_X2 U2139 ( .A(n3051), .ZN(n2918) );
  INV_X1 U2140 ( .A(n2073), .ZN(\DataP/alu_a_in[31] ) );
  INV_X1 U2141 ( .A(n2380), .ZN(\sra_131/SH[4] ) );
  INV_X2 U2142 ( .A(n2138), .ZN(n3206) );
  AND3_X1 U2143 ( .A1(n4061), .A2(n4060), .A3(n4059), .ZN(n1961) );
  BUF_X4 U2144 ( .A(\DataP/alu_b_in[2] ), .Z(n3202) );
  CLKBUF_X3 U2145 ( .A(n3203), .Z(n3051) );
  INV_X4 U2146 ( .A(n3046), .ZN(n2103) );
  OR2_X1 U2147 ( .A1(n2578), .A2(n3327), .ZN(\DataP/alu_a_in[3] ) );
  OR2_X4 U2148 ( .A1(n3356), .A2(n3355), .ZN(\DataP/alu_a_in[29] ) );
  AND2_X1 U2149 ( .A1(n3529), .A2(n3528), .ZN(n1963) );
  OR2_X1 U2150 ( .A1(ALU_OPCODE_i[2]), .A2(n2672), .ZN(n1964) );
  OR2_X2 U2151 ( .A1(n3385), .A2(n3384), .ZN(\DataP/alu_a_in[18] ) );
  OR2_X2 U2152 ( .A1(n3377), .A2(n3376), .ZN(\DataP/alu_a_in[21] ) );
  OR2_X1 U2153 ( .A1(n4110), .A2(n4199), .ZN(n1966) );
  NAND2_X2 U2154 ( .A1(n3433), .A2(n3561), .ZN(n3886) );
  AND2_X1 U2155 ( .A1(n2355), .A2(n2306), .ZN(n1967) );
  AND2_X1 U2156 ( .A1(\DataP/alu_a_in[6] ), .A2(n2039), .ZN(n1968) );
  OR2_X1 U2157 ( .A1(n3269), .A2(n3270), .ZN(n1970) );
  AND2_X1 U2158 ( .A1(n2066), .A2(n2062), .ZN(n1971) );
  OR2_X1 U2159 ( .A1(n2067), .A2(n2708), .ZN(n1972) );
  NOR2_X4 U2160 ( .A1(n3235), .A2(n2104), .ZN(n36) );
  INV_X1 U2161 ( .A(\CU_I/aluOpcode_i[4] ), .ZN(n2000) );
  BUF_X2 U2162 ( .A(\DataP/alu_a_in[3] ), .Z(n1973) );
  INV_X1 U2163 ( .A(\DataP/add_S2[2] ), .ZN(n1974) );
  NAND2_X1 U2166 ( .A1(n2009), .A2(n3479), .ZN(n3641) );
  NOR2_X1 U2167 ( .A1(\DataP/alu_b_in[8] ), .A2(\DataP/alu_b_in[9] ), .ZN(
        n2009) );
  NAND2_X1 U2168 ( .A1(n2010), .A2(n3483), .ZN(n3485) );
  OR2_X2 U2169 ( .A1(n2011), .A2(n2099), .ZN(n3483) );
  NAND2_X1 U2170 ( .A1(n3834), .A2(n3443), .ZN(n2010) );
  NAND2_X1 U2171 ( .A1(n2011), .A2(n2099), .ZN(n3443) );
  NAND2_X1 U2172 ( .A1(n3836), .A2(n2110), .ZN(n3834) );
  NAND2_X1 U2173 ( .A1(\DataP/ALU_C/comp/N24 ), .A2(n2012), .ZN(n2016) );
  AND2_X1 U2174 ( .A1(n3561), .A2(n2391), .ZN(n2012) );
  OAI211_X1 U2175 ( .C1(n2017), .C2(n2014), .A(n2013), .B(n2015), .ZN(n3567)
         );
  NOR2_X1 U2176 ( .A1(n3571), .A2(n2379), .ZN(n2015) );
  NAND2_X1 U2177 ( .A1(\DataP/ALU_C/comp/N50 ), .A2(ALU_OPCODE_i[2]), .ZN(
        n2017) );
  NAND2_X1 U2178 ( .A1(n2018), .A2(n2361), .ZN(\DataP/ALU_C/comp/N50 ) );
  NAND2_X1 U2179 ( .A1(n2019), .A2(n1967), .ZN(n2018) );
  NAND2_X1 U2180 ( .A1(n2363), .A2(n2362), .ZN(n2019) );
  AND2_X1 U2181 ( .A1(n2594), .A2(n2593), .ZN(n2576) );
  NAND2_X1 U2182 ( .A1(n2664), .A2(n2020), .ZN(n2594) );
  AND2_X1 U2183 ( .A1(n2710), .A2(n2720), .ZN(n2020) );
  NAND2_X1 U2184 ( .A1(n2021), .A2(n2750), .ZN(n2720) );
  OAI211_X1 U2185 ( .C1(n2025), .C2(n1574), .A(n2024), .B(n2022), .ZN(n2190)
         );
  INV_X1 U2186 ( .A(n2023), .ZN(n2022) );
  OAI21_X1 U2187 ( .B1(n2485), .B2(n2025), .A(n2722), .ZN(n2023) );
  NAND4_X1 U2188 ( .A1(n3709), .A2(n2485), .A3(\DataP/alu_b_in[26] ), .A4(
        n2108), .ZN(n2024) );
  NAND2_X1 U2189 ( .A1(n2127), .A2(n2108), .ZN(n2025) );
  NAND2_X1 U2190 ( .A1(n2075), .A2(n3841), .ZN(n2026) );
  NAND2_X1 U2191 ( .A1(n2245), .A2(n1735), .ZN(n3669) );
  NOR2_X1 U2192 ( .A1(n3640), .A2(n3641), .ZN(n2027) );
  XNOR2_X1 U2193 ( .A(n1965), .B(n536), .ZN(n2144) );
  NAND2_X1 U2194 ( .A1(n2028), .A2(Rst), .ZN(n2097) );
  XNOR2_X1 U2195 ( .A(n2778), .B(n2029), .ZN(n2028) );
  INV_X1 U2196 ( .A(\DataP/alu_b_in[7] ), .ZN(n2030) );
  NAND2_X1 U2197 ( .A1(n3423), .A2(n1748), .ZN(n2031) );
  AOI21_X1 U2198 ( .B1(n2037), .B2(n2032), .A(n2671), .ZN(n2670) );
  NAND2_X1 U2199 ( .A1(n2036), .A2(n2035), .ZN(n2034) );
  INV_X1 U2200 ( .A(n2293), .ZN(n2035) );
  NAND2_X1 U2201 ( .A1(n2291), .A2(n2292), .ZN(n2036) );
  NAND2_X1 U2202 ( .A1(n2038), .A2(n2395), .ZN(n2037) );
  OAI21_X1 U2203 ( .B1(n3571), .B2(\DataP/ALU_C/comp/N24 ), .A(ALU_OPCODE_i[1]), .ZN(n2038) );
  OAI211_X1 U2204 ( .C1(n2681), .C2(n3886), .A(n2680), .B(n3857), .ZN(n3609)
         );
  NAND2_X1 U2205 ( .A1(n2681), .A2(n2680), .ZN(n2040) );
  NAND2_X1 U2206 ( .A1(n2042), .A2(n1647), .ZN(n3618) );
  NAND2_X1 U2207 ( .A1(n3421), .A2(n2113), .ZN(n3604) );
  INV_X1 U2208 ( .A(n2371), .ZN(n2145) );
  NAND2_X1 U2209 ( .A1(n2581), .A2(n2052), .ZN(n2045) );
  OAI211_X1 U2210 ( .C1(n2581), .C2(n2053), .A(n2049), .B(n2045), .ZN(n2654)
         );
  OAI211_X1 U2211 ( .C1(n2581), .C2(n2047), .A(n2046), .B(n2564), .ZN(n2055)
         );
  NAND3_X1 U2212 ( .A1(n2048), .A2(n2581), .A3(n2049), .ZN(n2046) );
  NAND2_X1 U2213 ( .A1(n2049), .A2(n2053), .ZN(n2047) );
  OAI21_X1 U2214 ( .B1(n2051), .B2(n2236), .A(n2050), .ZN(n2049) );
  NAND2_X1 U2215 ( .A1(n2236), .A2(n2400), .ZN(n2050) );
  NOR2_X1 U2216 ( .A1(n2054), .A2(n2580), .ZN(n2051) );
  NOR2_X1 U2217 ( .A1(n1635), .A2(n2400), .ZN(n2052) );
  OR2_X1 U2218 ( .A1(n2236), .A2(n2054), .ZN(n2053) );
  INV_X1 U2219 ( .A(n2400), .ZN(n2054) );
  NAND2_X1 U2220 ( .A1(n2055), .A2(n2562), .ZN(\DataP/PC_reg/N30 ) );
  NAND4_X1 U2221 ( .A1(n2060), .A2(n2058), .A3(n2057), .A4(n2056), .ZN(
        \DataP/PC_reg/N25 ) );
  NAND2_X1 U2222 ( .A1(n1613), .A2(n1971), .ZN(n2056) );
  NAND2_X1 U2223 ( .A1(n3679), .A2(n2061), .ZN(n2057) );
  INV_X1 U2224 ( .A(n2059), .ZN(n2058) );
  OAI21_X1 U2225 ( .B1(n2064), .B2(n2708), .A(n1966), .ZN(n2059) );
  OR2_X1 U2226 ( .A1(n3777), .A2(n1972), .ZN(n2060) );
  INV_X1 U2227 ( .A(n4111), .ZN(n2061) );
  NOR2_X1 U2228 ( .A1(n3880), .A2(n4111), .ZN(n2062) );
  NOR2_X1 U2229 ( .A1(n2133), .A2(n1931), .ZN(n2066) );
  NAND2_X1 U2230 ( .A1(n2133), .A2(n1717), .ZN(n2067) );
  NAND4_X1 U2231 ( .A1(n3478), .A2(n3477), .A3(n3475), .A4(n3476), .ZN(
        \DataP/alu_b_in[12] ) );
  BUF_X1 U2232 ( .A(n3641), .Z(n2068) );
  BUF_X1 U2233 ( .A(n538), .Z(n2069) );
  OR2_X1 U2234 ( .A1(n2071), .A2(n2746), .ZN(n2070) );
  AOI21_X1 U2235 ( .B1(n2766), .B2(n2432), .A(n2765), .ZN(n2071) );
  AND2_X2 U2236 ( .A1(n2634), .A2(n3292), .ZN(n2072) );
  OR4_X2 U2237 ( .A1(n2259), .A2(n2261), .A3(n2309), .A4(n1602), .ZN(n2268) );
  AND2_X2 U2238 ( .A1(n2384), .A2(n2538), .ZN(n2073) );
  AND4_X1 U2239 ( .A1(n3322), .A2(n3321), .A3(n3319), .A4(n3320), .ZN(n2074)
         );
  AND2_X1 U2240 ( .A1(n1755), .A2(n2093), .ZN(n2076) );
  AND2_X1 U2241 ( .A1(n1755), .A2(n2093), .ZN(n3642) );
  OR2_X2 U2242 ( .A1(n3399), .A2(n2690), .ZN(\DataP/alu_a_in[11] ) );
  AOI22_X1 U2243 ( .A1(n3221), .A2(\DataP/B_s[0] ), .B1(n3222), .B2(
        \DataP/IMM_s[0] ), .ZN(n2077) );
  BUF_X1 U2244 ( .A(n2783), .Z(n2078) );
  BUF_X1 U2245 ( .A(\DataP/opcode_M[1] ), .Z(n2079) );
  OR2_X1 U2246 ( .A1(n2100), .A2(n2296), .ZN(n2080) );
  OR2_X1 U2247 ( .A1(\DataP/alu_b_in[2] ), .A2(n1719), .ZN(n2081) );
  INV_X1 U2248 ( .A(n3697), .ZN(\DataP/alu_a_in[27] ) );
  BUF_X1 U2249 ( .A(n3487), .Z(n2084) );
  AND4_X1 U2250 ( .A1(n2176), .A2(n2178), .A3(n2621), .A4(n2175), .ZN(n2085)
         );
  NOR2_X1 U2251 ( .A1(n3271), .A2(n1970), .ZN(n3272) );
  CLKBUF_X3 U2252 ( .A(n3402), .Z(n3217) );
  BUF_X1 U2253 ( .A(n2282), .Z(n2086) );
  NAND4_X1 U2254 ( .A1(n2143), .A2(n1962), .A3(n2144), .A4(n3240), .ZN(n2087)
         );
  AND2_X1 U2255 ( .A1(n2620), .A2(n2398), .ZN(n2088) );
  NOR2_X1 U2256 ( .A1(n2637), .A2(n2087), .ZN(n2089) );
  NAND4_X1 U2257 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n2090)
         );
  AND3_X1 U2258 ( .A1(n3239), .A2(\DataP/opcode_W[3] ), .A3(n2625), .ZN(n2091)
         );
  OAI221_X1 U2259 ( .B1(n2100), .B2(n2296), .C1(\DataP/alu_b_in[2] ), .C2(
        n1719), .A(n2313), .ZN(n2314) );
  NOR2_X1 U2260 ( .A1(\DataP/alu_b_in[13] ), .A2(\DataP/alu_b_in[12] ), .ZN(
        n3639) );
  NOR2_X1 U2261 ( .A1(n2098), .A2(n2659), .ZN(n2094) );
  BUF_X1 U2262 ( .A(n3860), .Z(n2095) );
  AND4_X2 U2263 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n2230)
         );
  INV_X1 U2264 ( .A(\DataP/alu_b_in[1] ), .ZN(n3200) );
  BUF_X4 U2265 ( .A(n3200), .Z(n3047) );
  INV_X1 U2266 ( .A(n2781), .ZN(n2782) );
  BUF_X2 U2267 ( .A(\DataP/alu_b_in[2] ), .Z(n3203) );
  AND2_X1 U2268 ( .A1(n2190), .A2(\DataP/alu_a_in[26] ), .ZN(n2096) );
  NAND4_X1 U2269 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n2098)
         );
  NAND2_X1 U2270 ( .A1(n3717), .A2(n3797), .ZN(n2484) );
  BUF_X1 U2271 ( .A(n2219), .Z(n2155) );
  INV_X1 U2272 ( .A(\DataP/alu_a_in[9] ), .ZN(n2099) );
  INV_X1 U2273 ( .A(n2101), .ZN(n2112) );
  INV_X1 U2274 ( .A(n3054), .ZN(n2115) );
  INV_X1 U2275 ( .A(n3203), .ZN(n3053) );
  OR2_X1 U2276 ( .A1(n3380), .A2(n3379), .ZN(\DataP/alu_a_in[20] ) );
  INV_X1 U2277 ( .A(n2226), .ZN(n2118) );
  INV_X1 U2278 ( .A(n2119), .ZN(n2100) );
  BUF_X4 U2279 ( .A(n3054), .Z(n2101) );
  INV_X2 U2280 ( .A(n2226), .ZN(n3199) );
  BUF_X2 U2281 ( .A(n4190), .Z(n2104) );
  BUF_X2 U2282 ( .A(n2126), .Z(n2105) );
  INV_X1 U2283 ( .A(n2372), .ZN(\DataP/alu_b_in[7] ) );
  INV_X1 U2284 ( .A(n2141), .ZN(n2106) );
  INV_X1 U2285 ( .A(\DataP/alu_b_in[24] ), .ZN(n2107) );
  AND2_X1 U2286 ( .A1(n2389), .A2(n2133), .ZN(n2193) );
  INV_X1 U2287 ( .A(\DataP/alu_a_in[13] ), .ZN(n2109) );
  INV_X1 U2288 ( .A(\DataP/alu_a_in[8] ), .ZN(n2110) );
  INV_X1 U2289 ( .A(\DataP/alu_a_in[21] ), .ZN(n2111) );
  INV_X1 U2290 ( .A(\DataP/alu_a_in[5] ), .ZN(n2113) );
  INV_X1 U2291 ( .A(\DataP/alu_a_in[20] ), .ZN(n2114) );
  NAND2_X1 U2292 ( .A1(n2139), .A2(n1969), .ZN(n2150) );
  INV_X1 U2293 ( .A(\DataP/alu_a_in[11] ), .ZN(n2116) );
  OR2_X1 U2294 ( .A1(n3908), .A2(\DataP/wrong_br ), .ZN(n4190) );
  BUF_X2 U2295 ( .A(n3046), .Z(n2117) );
  INV_X1 U2296 ( .A(\DataP/alu_b_in[3] ), .ZN(n2119) );
  INV_X1 U2297 ( .A(\DataP/alu_b_in[28] ), .ZN(n2120) );
  NAND2_X1 U2298 ( .A1(\DataP/alu_b_in[22] ), .A2(n3886), .ZN(n2402) );
  BUF_X1 U2299 ( .A(\DataP/alu_b_in[21] ), .Z(n2152) );
  NAND4_X1 U2300 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(
        \DataP/alu_b_in[9] ) );
  NAND4_X1 U2301 ( .A1(n3442), .A2(n3441), .A3(n3439), .A4(n3440), .ZN(
        \DataP/alu_b_in[10] ) );
  INV_X1 U2302 ( .A(\DataP/alu_b_in[31] ), .ZN(n2121) );
  INV_X1 U2303 ( .A(\DataP/alu_b_in[22] ), .ZN(n2122) );
  INV_X1 U2304 ( .A(\DataP/alu_b_in[18] ), .ZN(n2123) );
  INV_X1 U2305 ( .A(\DataP/alu_b_in[23] ), .ZN(n2124) );
  INV_X1 U2306 ( .A(n3212), .ZN(n3211) );
  INV_X1 U2307 ( .A(\DataP/alu_b_in[29] ), .ZN(n2125) );
  INV_X1 U2308 ( .A(n1601), .ZN(n2126) );
  INV_X1 U2309 ( .A(\DataP/alu_b_in[26] ), .ZN(n2127) );
  INV_X1 U2310 ( .A(n3897), .ZN(n2130) );
  INV_X1 U2311 ( .A(n4111), .ZN(n2131) );
  NOR2_X1 U2312 ( .A1(n3246), .A2(n2628), .ZN(n2627) );
  AND4_X1 U2313 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n2386)
         );
  INV_X2 U2314 ( .A(n3233), .ZN(n2132) );
  AND2_X1 U2315 ( .A1(n3884), .A2(n2489), .ZN(n2755) );
  AND2_X1 U2316 ( .A1(n2764), .A2(n2760), .ZN(n2759) );
  INV_X1 U2317 ( .A(n2758), .ZN(n3635) );
  AND3_X1 U2318 ( .A1(n2168), .A2(n2155), .A3(n2167), .ZN(n2763) );
  AND2_X1 U2319 ( .A1(n3728), .A2(n2365), .ZN(n3826) );
  NAND2_X1 U2320 ( .A1(n2586), .A2(n2186), .ZN(n3797) );
  INV_X1 U2321 ( .A(n3713), .ZN(n2133) );
  NOR2_X1 U2322 ( .A1(\DataP/alu_a_in[25] ), .A2(n2187), .ZN(n2186) );
  INV_X1 U2323 ( .A(n4190), .ZN(n3231) );
  INV_X1 U2324 ( .A(n4190), .ZN(n3230) );
  AND2_X1 U2325 ( .A1(\DataP/alu_a_in[9] ), .A2(n3429), .ZN(n2259) );
  BUF_X1 U2326 ( .A(\DataP/alu_a_in[9] ), .Z(n2207) );
  AND2_X1 U2327 ( .A1(\DataP/alu_a_in[16] ), .A2(n2198), .ZN(n2197) );
  INV_X1 U2328 ( .A(n2182), .ZN(n2181) );
  INV_X1 U2329 ( .A(\DataP/alu_a_in[12] ), .ZN(n2134) );
  OAI21_X1 U2330 ( .B1(n2703), .B2(n2185), .A(n2108), .ZN(n2182) );
  INV_X1 U2331 ( .A(n2101), .ZN(n3205) );
  AND2_X1 U2332 ( .A1(n2703), .A2(n2185), .ZN(n2184) );
  BUF_X1 U2333 ( .A(\DataP/alu_a_in[11] ), .Z(n2200) );
  OR2_X1 U2334 ( .A1(n3368), .A2(n3367), .ZN(\DataP/alu_a_in[24] ) );
  OR2_X1 U2335 ( .A1(n3362), .A2(n3361), .ZN(\DataP/alu_a_in[26] ) );
  INV_X1 U2336 ( .A(\DataP/alu_a_in[18] ), .ZN(n2135) );
  OR2_X1 U2337 ( .A1(n3359), .A2(n3358), .ZN(\DataP/alu_a_in[28] ) );
  INV_X1 U2338 ( .A(\DataP/alu_a_in[23] ), .ZN(n2136) );
  OR2_X2 U2339 ( .A1(n3382), .A2(n3381), .ZN(\DataP/alu_a_in[19] ) );
  INV_X1 U2340 ( .A(\DataP/alu_a_in[25] ), .ZN(n2137) );
  INV_X1 U2341 ( .A(\DataP/alu_b_in[3] ), .ZN(n3054) );
  INV_X1 U2342 ( .A(n2226), .ZN(n2916) );
  INV_X1 U2343 ( .A(n2585), .ZN(n2187) );
  INV_X1 U2344 ( .A(n3212), .ZN(n2209) );
  INV_X1 U2345 ( .A(n2230), .ZN(\DataP/alu_b_in[15] ) );
  BUF_X1 U2346 ( .A(n1591), .Z(n2166) );
  INV_X1 U2347 ( .A(n3214), .ZN(n2139) );
  INV_X1 U2348 ( .A(\DataP/alu_b_in[6] ), .ZN(n2140) );
  BUF_X2 U2349 ( .A(n1550), .Z(n2141) );
  INV_X1 U2350 ( .A(n2782), .ZN(n2772) );
  AND3_X1 U2351 ( .A1(n3549), .A2(n3259), .A3(n399), .ZN(n3547) );
  OAI21_X1 U2352 ( .B1(n4148), .B2(n4147), .A(Rst), .ZN(n4149) );
  OR2_X1 U2353 ( .A1(n4153), .A2(\CU_I/cw[7] ), .ZN(n4147) );
  NOR2_X1 U2354 ( .A1(n4052), .A2(n4051), .ZN(\CU_I/cw[7] ) );
  AND2_X1 U2355 ( .A1(n2237), .A2(n2639), .ZN(n2398) );
  NAND2_X2 U2356 ( .A1(n3438), .A2(Rst), .ZN(n4110) );
  OR2_X2 U2357 ( .A1(n3229), .A2(n4143), .ZN(n4146) );
  NAND2_X1 U2358 ( .A1(n2626), .A2(n2627), .ZN(n3291) );
  INV_X1 U2359 ( .A(n3883), .ZN(n2626) );
  AND2_X2 U2360 ( .A1(\WB_MUX_SEL_i[1] ), .A2(n294), .ZN(n4143) );
  CLKBUF_X1 U2361 ( .A(\DataP/add_D[3] ), .Z(n2146) );
  INV_X4 U2362 ( .A(n2380), .ZN(n3055) );
  NAND2_X2 U2363 ( .A1(n3432), .A2(n3435), .ZN(n3897) );
  NOR2_X1 U2364 ( .A1(n2637), .A2(n2142), .ZN(n2636) );
  NAND4_X1 U2365 ( .A1(n2143), .A2(n1962), .A3(n2144), .A4(n3240), .ZN(n2142)
         );
  AND2_X1 U2366 ( .A1(n2174), .A2(n2636), .ZN(n2620) );
  OAI211_X1 U2367 ( .C1(n3213), .C2(n41), .A(n2149), .B(n2148), .ZN(n3334) );
  NAND2_X1 U2368 ( .A1(n3210), .A2(DRAM_ADDRESS[1]), .ZN(n2148) );
  NAND2_X1 U2369 ( .A1(n3209), .A2(\DataP/alu_out_W[1] ), .ZN(n2149) );
  NOR2_X1 U2370 ( .A1(n2090), .A2(n2659), .ZN(n2658) );
  AND4_X2 U2371 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n2242)
         );
  NAND2_X1 U2372 ( .A1(n3396), .A2(n2150), .ZN(n3398) );
  NAND4_X4 U2373 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(
        \DataP/alu_b_in[16] ) );
  AOI21_X1 U2374 ( .B1(n3843), .B2(n3420), .A(n3419), .ZN(n3426) );
  NAND2_X1 U2375 ( .A1(n3845), .A2(n3844), .ZN(n3843) );
  NAND2_X1 U2376 ( .A1(n2154), .A2(n2153), .ZN(n3412) );
  NAND2_X1 U2377 ( .A1(n3054), .A2(n3886), .ZN(n2153) );
  NAND2_X1 U2378 ( .A1(n3411), .A2(n2108), .ZN(n2154) );
  NAND2_X1 U2379 ( .A1(n3869), .A2(n3630), .ZN(n2666) );
  NAND2_X1 U2380 ( .A1(n2642), .A2(n3629), .ZN(n3869) );
  NAND2_X1 U2381 ( .A1(n2158), .A2(n2157), .ZN(n3646) );
  NAND2_X1 U2382 ( .A1(n2370), .A2(n3886), .ZN(n2157) );
  NAND2_X1 U2383 ( .A1(n3644), .A2(n2108), .ZN(n2158) );
  NOR2_X1 U2384 ( .A1(n2159), .A2(n2488), .ZN(n2557) );
  NAND2_X1 U2385 ( .A1(n2161), .A2(n2160), .ZN(n2159) );
  NAND2_X1 U2386 ( .A1(\DataP/ALU_C/shifter/N49 ), .A2(n3228), .ZN(n2160) );
  INV_X1 U2387 ( .A(n3903), .ZN(n2161) );
  OAI21_X1 U2388 ( .B1(n2533), .B2(n2531), .A(n2162), .ZN(n2602) );
  NAND2_X1 U2389 ( .A1(n3763), .A2(n1746), .ZN(n2162) );
  NAND2_X1 U2390 ( .A1(n1738), .A2(n3691), .ZN(n2213) );
  NAND2_X1 U2391 ( .A1(n2074), .A2(n3886), .ZN(n2163) );
  BUF_X1 U2392 ( .A(n1752), .Z(n2164) );
  CLKBUF_X1 U2393 ( .A(n1566), .Z(n2168) );
  OAI211_X1 U2394 ( .C1(n3662), .C2(n3682), .A(n1566), .B(n2169), .ZN(n3687)
         );
  NAND2_X1 U2395 ( .A1(n2549), .A2(n2547), .ZN(n2169) );
  NAND2_X1 U2396 ( .A1(n2546), .A2(n2108), .ZN(n2549) );
  XNOR2_X1 U2397 ( .A(n3647), .B(n1736), .ZN(n2546) );
  NOR2_X1 U2398 ( .A1(n3694), .A2(n3659), .ZN(n3647) );
  NAND2_X1 U2399 ( .A1(n3643), .A2(n2721), .ZN(n2173) );
  OAI211_X1 U2400 ( .C1(\DataP/alu_b_in[17] ), .C2(n1738), .A(n2170), .B(n2172), .ZN(n3643) );
  NAND2_X1 U2401 ( .A1(n2245), .A2(n2171), .ZN(n2170) );
  AND2_X1 U2402 ( .A1(\DataP/alu_b_in[17] ), .A2(n2370), .ZN(n2171) );
  NAND2_X1 U2403 ( .A1(\DataP/alu_b_in[16] ), .A2(n1753), .ZN(n2172) );
  NAND2_X1 U2404 ( .A1(n2173), .A2(n2528), .ZN(n3661) );
  AND2_X1 U2405 ( .A1(n3289), .A2(n2638), .ZN(n2174) );
  NAND3_X1 U2406 ( .A1(n2174), .A2(n2089), .A3(n2639), .ZN(n3258) );
  NOR2_X1 U2407 ( .A1(n2097), .A2(n2406), .ZN(n2175) );
  NAND2_X1 U2408 ( .A1(n3250), .A2(n3251), .ZN(n2176) );
  NAND2_X1 U2409 ( .A1(n2177), .A2(n3248), .ZN(n3251) );
  INV_X1 U2410 ( .A(n2179), .ZN(n2177) );
  NOR2_X1 U2411 ( .A1(n3883), .A2(n3246), .ZN(n2178) );
  NAND4_X1 U2412 ( .A1(n520), .A2(n17), .A3(n19), .A4(n21), .ZN(n3883) );
  NAND2_X1 U2413 ( .A1(n521), .A2(n23), .ZN(n3246) );
  OAI211_X1 U2414 ( .C1(n22), .C2(n2079), .A(n2180), .B(n2387), .ZN(n2179) );
  NAND2_X1 U2415 ( .A1(\DataP/opcode_M[1] ), .A2(\DataP/opcode_M[3] ), .ZN(
        n2180) );
  NAND2_X1 U2416 ( .A1(n3709), .A2(n2184), .ZN(n2183) );
  OAI211_X1 U2417 ( .C1(n2185), .C2(n1574), .A(n2183), .B(n2181), .ZN(n2189)
         );
  INV_X1 U2418 ( .A(\DataP/alu_b_in[27] ), .ZN(n2185) );
  XNOR2_X1 U2419 ( .A(n3720), .B(n3697), .ZN(n2188) );
  NAND2_X1 U2420 ( .A1(n2189), .A2(n2540), .ZN(n3720) );
  NAND3_X1 U2421 ( .A1(n2192), .A2(n3690), .A3(n2193), .ZN(n2191) );
  NAND2_X1 U2422 ( .A1(n1633), .A2(n1717), .ZN(n2192) );
  AND4_X2 U2423 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n2372)
         );
  NAND4_X1 U2424 ( .A1(n3307), .A2(n1583), .A3(n3305), .A4(n3304), .ZN(
        \DataP/alu_b_in[1] ) );
  OAI211_X1 U2425 ( .C1(\DataP/opcode_M[4] ), .C2(\DataP/opcode_M[0] ), .A(
        \DataP/opcode_M[1] ), .B(\DataP/opcode_M[2] ), .ZN(n2195) );
  NAND2_X1 U2426 ( .A1(n2196), .A2(n2197), .ZN(n3738) );
  NAND2_X1 U2427 ( .A1(n3644), .A2(n2534), .ZN(n2196) );
  XNOR2_X1 U2428 ( .A(n1760), .B(\DataP/alu_b_in[16] ), .ZN(n3644) );
  NAND2_X1 U2429 ( .A1(n2534), .A2(n2535), .ZN(n2198) );
  NAND2_X1 U2430 ( .A1(n3738), .A2(n3660), .ZN(n2527) );
  OAI21_X1 U2431 ( .B1(n3643), .B2(n2128), .A(n2397), .ZN(n3660) );
  OAI21_X1 U2432 ( .B1(n2673), .B2(n2234), .A(n2674), .ZN(n2199) );
  INV_X1 U2433 ( .A(n3537), .ZN(n2201) );
  NOR2_X1 U2434 ( .A1(n3382), .A2(n3381), .ZN(n2202) );
  BUF_X1 U2435 ( .A(n3855), .Z(n2203) );
  BUF_X1 U2436 ( .A(n3836), .Z(n2204) );
  AND2_X1 U2437 ( .A1(n3443), .A2(n1749), .ZN(n2205) );
  BUF_X2 U2438 ( .A(n3401), .Z(n3215) );
  INV_X1 U2439 ( .A(n3617), .ZN(n2208) );
  NOR2_X1 U2440 ( .A1(n3389), .A2(n2693), .ZN(n2210) );
  BUF_X1 U2441 ( .A(n3611), .Z(n2211) );
  XNOR2_X1 U2442 ( .A(n3799), .B(n2212), .ZN(n3806) );
  OR2_X1 U2443 ( .A1(n2744), .A2(n3798), .ZN(n2212) );
  BUF_X1 U2444 ( .A(n3869), .Z(n2214) );
  BUF_X1 U2445 ( .A(n3604), .Z(n2215) );
  AND2_X1 U2446 ( .A1(n2594), .A2(n2593), .ZN(n2216) );
  AOI21_X1 U2447 ( .B1(n2560), .B2(n2129), .A(n3679), .ZN(n2217) );
  BUF_X1 U2448 ( .A(n1584), .Z(n2218) );
  AND2_X1 U2449 ( .A1(n2525), .A2(n2524), .ZN(n2220) );
  OR2_X2 U2450 ( .A1(n3330), .A2(n3329), .ZN(\DataP/alu_a_in[2] ) );
  BUF_X1 U2451 ( .A(n1749), .Z(n2221) );
  AND2_X1 U2452 ( .A1(n3485), .A2(n3484), .ZN(n2222) );
  INV_X1 U2453 ( .A(n2234), .ZN(n2223) );
  INV_X1 U2454 ( .A(n1746), .ZN(n2224) );
  AND2_X1 U2455 ( .A1(n2687), .A2(n2686), .ZN(n2225) );
  BUF_X1 U2456 ( .A(n3221), .Z(n2227) );
  BUF_X2 U2457 ( .A(\DataP/alu_a_in[0] ), .Z(n2231) );
  OR2_X2 U2458 ( .A1(n3334), .A2(n3333), .ZN(n2232) );
  NAND2_X1 U2459 ( .A1(n2077), .A2(n1593), .ZN(n2233) );
  NAND2_X1 U2460 ( .A1(n2656), .A2(n2657), .ZN(\DataP/alu_b_in[0] ) );
  AND2_X1 U2461 ( .A1(n3308), .A2(n3309), .ZN(n2657) );
  AND3_X1 U2462 ( .A1(n1634), .A2(n2611), .A3(n2609), .ZN(n2234) );
  NAND2_X1 U2463 ( .A1(n3464), .A2(n3491), .ZN(n2235) );
  AND2_X1 U2464 ( .A1(n2583), .A2(n2582), .ZN(n2236) );
  AND2_X1 U2465 ( .A1(n2627), .A2(n2626), .ZN(n2237) );
  AND3_X2 U2466 ( .A1(n3549), .A2(n3259), .A3(n2481), .ZN(n3548) );
  INV_X1 U2467 ( .A(n2762), .ZN(n2238) );
  BUF_X1 U2468 ( .A(n3738), .Z(n2239) );
  BUF_X2 U2469 ( .A(n3402), .Z(n3218) );
  OAI21_X1 U2470 ( .B1(n2096), .B2(n3719), .A(n2188), .ZN(n2241) );
  AOI21_X1 U2471 ( .B1(n1733), .B2(n2491), .A(n2668), .ZN(n2243) );
  OAI221_X1 U2472 ( .B1(n2293), .B2(n2292), .C1(n2291), .C2(n2293), .A(n2290), 
        .ZN(\DataP/ALU_C/comp/N24 ) );
  NOR2_X1 U2473 ( .A1(n1760), .A2(n3659), .ZN(n2244) );
  BUF_X2 U2474 ( .A(n3548), .Z(n2246) );
  BUF_X2 U2475 ( .A(n3548), .Z(n2247) );
  AOI21_X1 U2476 ( .B1(n3251), .B2(n3250), .A(n2406), .ZN(n2248) );
  NAND4_X1 U2477 ( .A1(n3307), .A2(n1583), .A3(n3305), .A4(n3304), .ZN(n2250)
         );
  NOR2_X1 U2478 ( .A1(\DataP/alu_b_in[29] ), .A2(n2295), .ZN(n2252) );
  NAND2_X1 U2479 ( .A1(\DataP/alu_b_in[31] ), .A2(n2073), .ZN(n2251) );
  OAI21_X1 U2480 ( .B1(\DataP/alu_b_in[30] ), .B2(n2294), .A(n2251), .ZN(n2280) );
  AOI211_X1 U2481 ( .C1(\DataP/alu_a_in[28] ), .C2(n2120), .A(n2252), .B(n2280), .ZN(n2284) );
  AOI211_X1 U2482 ( .C1(\DataP/alu_a_in[24] ), .C2(n2107), .A(n2086), .B(n2297), .ZN(n2253) );
  NAND2_X1 U2483 ( .A1(n2284), .A2(n2253), .ZN(n2293) );
  AOI21_X1 U2484 ( .B1(\DataP/alu_a_in[14] ), .B2(n2371), .A(n2307), .ZN(n2267) );
  OAI211_X1 U2485 ( .C1(\lt_x_135/B[12] ), .C2(n2134), .A(n2308), .B(n2267), 
        .ZN(n2261) );
  AOI21_X1 U2486 ( .B1(\DataP/alu_a_in[6] ), .B2(n2140), .A(n2311), .ZN(n2257)
         );
  OAI22_X1 U2487 ( .A1(n2231), .A2(n2312), .B1(n2232), .B2(n2126), .ZN(n2254)
         );
  OAI22_X1 U2488 ( .A1(\DataP/alu_a_in[6] ), .A2(n2318), .B1(
        \DataP/alu_a_in[7] ), .B2(n2030), .ZN(n2255) );
  OAI22_X1 U2489 ( .A1(\DataP/alu_a_in[12] ), .A2(n2321), .B1(
        \DataP/alu_a_in[13] ), .B2(n2106), .ZN(n2266) );
  NOR2_X1 U2490 ( .A1(n2322), .A2(\DataP/alu_a_in[10] ), .ZN(n2258) );
  AOI22_X1 U2491 ( .A1(n2165), .A2(n2258), .B1(n2151), .B2(n2116), .ZN(n2263)
         );
  NOR2_X1 U2492 ( .A1(\DataP/alu_a_in[8] ), .A2(n2259), .ZN(n2260) );
  AOI22_X1 U2493 ( .A1(n2164), .A2(n2260), .B1(n2166), .B2(n2099), .ZN(n2262)
         );
  AOI221_X1 U2494 ( .B1(n1602), .B2(n2263), .C1(n2263), .C2(n2262), .A(n2261), 
        .ZN(n2265) );
  NOR2_X1 U2495 ( .A1(\DataP/alu_b_in[17] ), .A2(n1750), .ZN(n2272) );
  OAI211_X1 U2496 ( .C1(\DataP/alu_b_in[20] ), .C2(n2114), .A(n2279), .B(n2338), .ZN(n2274) );
  AOI21_X1 U2497 ( .B1(n2123), .B2(\DataP/alu_a_in[18] ), .A(n2341), .ZN(n2269) );
  OAI21_X1 U2498 ( .B1(n2152), .B2(n2111), .A(\DataP/alu_b_in[20] ), .ZN(n2270) );
  OAI22_X1 U2499 ( .A1(\DataP/alu_a_in[20] ), .A2(n2270), .B1(
        \DataP/alu_a_in[21] ), .B2(n3663), .ZN(n2278) );
  NOR2_X1 U2500 ( .A1(n2341), .A2(\DataP/alu_a_in[18] ), .ZN(n2271) );
  AOI22_X1 U2501 ( .A1(n2271), .A2(n1736), .B1(n1722), .B2(n2202), .ZN(n2276)
         );
  NOR2_X1 U2502 ( .A1(\DataP/alu_a_in[16] ), .A2(n2272), .ZN(n2273) );
  AOI22_X1 U2503 ( .A1(\DataP/alu_b_in[16] ), .A2(n2273), .B1(
        \DataP/alu_b_in[17] ), .B2(n1750), .ZN(n2275) );
  AOI221_X1 U2504 ( .B1(n2298), .B2(n2276), .C1(n2275), .C2(n2276), .A(n2274), 
        .ZN(n2277) );
  OAI21_X1 U2505 ( .B1(\DataP/alu_b_in[29] ), .B2(n2295), .A(
        \DataP/alu_b_in[28] ), .ZN(n2281) );
  OAI22_X1 U2506 ( .A1(\DataP/alu_a_in[28] ), .A2(n2281), .B1(
        \DataP/alu_a_in[29] ), .B2(n2125), .ZN(n2289) );
  AOI22_X1 U2507 ( .A1(\DataP/alu_b_in[26] ), .A2(n2354), .B1(
        \DataP/alu_b_in[27] ), .B2(n3697), .ZN(n2285) );
  NOR2_X1 U2508 ( .A1(\DataP/alu_a_in[24] ), .A2(n2282), .ZN(n2283) );
  AOI221_X1 U2509 ( .B1(n2297), .B2(n2285), .C1(n2356), .C2(n2285), .A(n2300), 
        .ZN(n2288) );
  OAI21_X1 U2510 ( .B1(\DataP/alu_a_in[31] ), .B2(n2121), .A(
        \DataP/alu_b_in[30] ), .ZN(n2286) );
  OAI22_X1 U2511 ( .A1(\DataP/alu_a_in[30] ), .A2(n2286), .B1(
        \DataP/alu_b_in[31] ), .B2(n2073), .ZN(n2287) );
  AND2_X1 U2512 ( .A1(\DataP/alu_a_in[22] ), .A2(n2122), .ZN(n2302) );
  INV_X1 U2513 ( .A(\DataP/alu_a_in[29] ), .ZN(n2295) );
  INV_X1 U2514 ( .A(\DataP/alu_a_in[30] ), .ZN(n2294) );
  INV_X1 U2515 ( .A(\DataP/alu_a_in[3] ), .ZN(n2296) );
  INV_X1 U2516 ( .A(\DataP/alu_b_in[16] ), .ZN(n2301) );
  AOI21_X1 U2517 ( .B1(\DataP/alu_a_in[23] ), .B2(n2124), .A(n2302), .ZN(n2279) );
  INV_X1 U2518 ( .A(n2269), .ZN(n2298) );
  INV_X1 U2519 ( .A(n2280), .ZN(n2299) );
  INV_X1 U2520 ( .A(n2284), .ZN(n2300) );
  NOR2_X1 U2521 ( .A1(\DataP/alu_b_in[29] ), .A2(n2365), .ZN(n2304) );
  NAND2_X1 U2522 ( .A1(\DataP/alu_a_in[31] ), .A2(n2121), .ZN(n2303) );
  OAI21_X1 U2523 ( .B1(\DataP/alu_b_in[30] ), .B2(n2364), .A(n2303), .ZN(n2351) );
  AOI211_X1 U2524 ( .C1(\DataP/alu_a_in[28] ), .C2(n2120), .A(n2304), .B(n2351), .ZN(n2355) );
  NOR2_X1 U2525 ( .A1(n3697), .A2(\DataP/alu_b_in[27] ), .ZN(n2353) );
  AOI21_X1 U2526 ( .B1(n2127), .B2(\DataP/alu_a_in[26] ), .A(n2353), .ZN(n2305) );
  AOI211_X1 U2527 ( .C1(\DataP/alu_a_in[24] ), .C2(n2107), .A(n2086), .B(n2367), .ZN(n2306) );
  NOR2_X1 U2528 ( .A1(n2166), .A2(n2099), .ZN(n2324) );
  NOR2_X1 U2529 ( .A1(\DataP/alu_b_in[15] ), .A2(n2210), .ZN(n2307) );
  AOI21_X1 U2530 ( .B1(\DataP/alu_a_in[14] ), .B2(n2371), .A(n2307), .ZN(n2333) );
  NAND2_X1 U2531 ( .A1(\DataP/alu_a_in[13] ), .A2(n2106), .ZN(n2308) );
  OAI211_X1 U2532 ( .C1(\lt_x_135/B[12] ), .C2(n2134), .A(n2333), .B(n2308), 
        .ZN(n2326) );
  NOR2_X1 U2533 ( .A1(n2164), .A2(n2110), .ZN(n2309) );
  NOR2_X1 U2534 ( .A1(n2151), .A2(n2116), .ZN(n2322) );
  OR4_X1 U2535 ( .A1(n2324), .A2(n2326), .A3(n2309), .A4(n1602), .ZN(n2336) );
  OAI21_X1 U2536 ( .B1(\lt_x_135/B[5] ), .B2(n2113), .A(n2138), .ZN(n2310) );
  OAI22_X1 U2537 ( .A1(\DataP/alu_a_in[4] ), .A2(n2310), .B1(
        \DataP/alu_a_in[5] ), .B2(n2074), .ZN(n2320) );
  NOR2_X1 U2538 ( .A1(n2366), .A2(\DataP/alu_b_in[7] ), .ZN(n2311) );
  OAI21_X1 U2539 ( .B1(n2100), .B2(n2296), .A(\DataP/alu_b_in[2] ), .ZN(n2315)
         );
  OAI21_X1 U2540 ( .B1(n2373), .B2(n2206), .A(n2226), .ZN(n2312) );
  OAI22_X1 U2541 ( .A1(n2231), .A2(n2312), .B1(n2232), .B2(n2126), .ZN(n2313)
         );
  OAI221_X1 U2542 ( .B1(n1973), .B2(n2119), .C1(\DataP/alu_a_in[2] ), .C2(
        n2315), .A(n2314), .ZN(n2316) );
  OAI21_X1 U2543 ( .B1(\lt_x_135/B[5] ), .B2(n2113), .A(n2316), .ZN(n2317) );
  AOI21_X1 U2544 ( .B1(\DataP/alu_a_in[4] ), .B2(n3206), .A(n2317), .ZN(n2319)
         );
  OAI21_X1 U2545 ( .B1(n2366), .B2(\DataP/alu_b_in[7] ), .A(
        \DataP/alu_b_in[6] ), .ZN(n2318) );
  AOI221_X1 U2546 ( .B1(n2320), .B2(n2257), .C1(n2319), .C2(n2257), .A(n2255), 
        .ZN(n2335) );
  OAI21_X1 U2547 ( .B1(n2141), .B2(n2109), .A(\lt_x_135/B[12] ), .ZN(n2321) );
  OAI22_X1 U2548 ( .A1(\DataP/alu_a_in[12] ), .A2(n2321), .B1(
        \DataP/alu_a_in[13] ), .B2(n2106), .ZN(n2332) );
  NOR2_X1 U2549 ( .A1(\DataP/alu_a_in[10] ), .A2(n2322), .ZN(n2323) );
  AOI22_X1 U2550 ( .A1(n2165), .A2(n2323), .B1(n2151), .B2(n2116), .ZN(n2328)
         );
  NOR2_X1 U2551 ( .A1(\DataP/alu_a_in[8] ), .A2(n2324), .ZN(n2325) );
  AOI22_X1 U2552 ( .A1(n2164), .A2(n2325), .B1(n2166), .B2(n2099), .ZN(n2327)
         );
  AOI221_X1 U2553 ( .B1(n1602), .B2(n2328), .C1(n2327), .C2(n2328), .A(n2326), 
        .ZN(n2331) );
  OAI22_X1 U2554 ( .A1(\DataP/alu_a_in[14] ), .A2(n2329), .B1(
        \DataP/alu_a_in[15] ), .B2(n2230), .ZN(n2330) );
  AOI211_X1 U2555 ( .C1(n2333), .C2(n2332), .A(n2331), .B(n2330), .ZN(n2334)
         );
  OAI21_X1 U2556 ( .B1(n2336), .B2(n2335), .A(n2334), .ZN(n2340) );
  NOR2_X1 U2557 ( .A1(\DataP/alu_b_in[17] ), .A2(n1750), .ZN(n2342) );
  NOR2_X1 U2558 ( .A1(\DataP/alu_b_in[23] ), .A2(n2136), .ZN(n2337) );
  AOI21_X1 U2559 ( .B1(\DataP/alu_a_in[22] ), .B2(n2122), .A(n2337), .ZN(n2350) );
  NAND2_X1 U2560 ( .A1(\DataP/alu_a_in[21] ), .A2(n3663), .ZN(n2338) );
  OAI211_X1 U2561 ( .C1(\DataP/alu_b_in[20] ), .C2(n2114), .A(n2350), .B(n2338), .ZN(n2344) );
  NOR2_X1 U2562 ( .A1(n1722), .A2(n2202), .ZN(n2341) );
  AOI211_X1 U2563 ( .C1(\DataP/alu_a_in[16] ), .C2(n2370), .A(n2344), .B(n2298), .ZN(n2339) );
  NAND3_X1 U2564 ( .A1(n2340), .A2(n2369), .A3(n2339), .ZN(n2363) );
  NOR2_X1 U2565 ( .A1(\DataP/alu_a_in[16] ), .A2(n2342), .ZN(n2343) );
  AOI22_X1 U2566 ( .A1(\DataP/alu_b_in[16] ), .A2(n2343), .B1(
        \DataP/alu_b_in[17] ), .B2(n1750), .ZN(n2345) );
  AOI221_X1 U2567 ( .B1(n2298), .B2(n2346), .C1(n2345), .C2(n2346), .A(n2344), 
        .ZN(n2349) );
  OAI21_X1 U2568 ( .B1(\DataP/alu_b_in[23] ), .B2(n2136), .A(
        \DataP/alu_b_in[22] ), .ZN(n2347) );
  OAI22_X1 U2569 ( .A1(\DataP/alu_a_in[22] ), .A2(n2347), .B1(
        \DataP/alu_a_in[23] ), .B2(n2124), .ZN(n2348) );
  AOI211_X1 U2570 ( .C1(n2350), .C2(n2278), .A(n2349), .B(n2348), .ZN(n2362)
         );
  OAI21_X1 U2571 ( .B1(\DataP/alu_b_in[29] ), .B2(n2365), .A(
        \DataP/alu_b_in[28] ), .ZN(n2352) );
  OAI22_X1 U2572 ( .A1(\DataP/alu_a_in[28] ), .A2(n2352), .B1(
        \DataP/alu_a_in[29] ), .B2(n2125), .ZN(n2360) );
  NOR2_X1 U2573 ( .A1(\DataP/alu_a_in[26] ), .A2(n2353), .ZN(n2354) );
  OAI21_X1 U2574 ( .B1(\DataP/alu_b_in[31] ), .B2(n2073), .A(
        \DataP/alu_b_in[30] ), .ZN(n2357) );
  OAI22_X1 U2575 ( .A1(\DataP/alu_a_in[30] ), .A2(n2357), .B1(
        \DataP/alu_a_in[31] ), .B2(n2121), .ZN(n2358) );
  AOI211_X1 U2576 ( .C1(n2368), .C2(n2360), .A(n2359), .B(n2358), .ZN(n2361)
         );
  INV_X1 U2577 ( .A(n2126), .ZN(n2373) );
  INV_X1 U2578 ( .A(\DataP/alu_a_in[29] ), .ZN(n2365) );
  INV_X1 U2579 ( .A(\DataP/alu_a_in[30] ), .ZN(n2364) );
  INV_X1 U2580 ( .A(n2305), .ZN(n2367) );
  INV_X1 U2581 ( .A(\DataP/alu_a_in[7] ), .ZN(n2366) );
  INV_X1 U2582 ( .A(n2342), .ZN(n2369) );
  INV_X1 U2583 ( .A(\DataP/alu_b_in[16] ), .ZN(n2370) );
  INV_X1 U2584 ( .A(n2351), .ZN(n2368) );
  NAND2_X1 U2585 ( .A1(n2620), .A2(n2398), .ZN(n3259) );
  INV_X1 U2586 ( .A(\DataP/alu_b_in[20] ), .ZN(n3664) );
  INV_X1 U2587 ( .A(\DataP/alu_b_in[21] ), .ZN(n3663) );
  BUF_X2 U2588 ( .A(n3547), .Z(n3219) );
  NOR2_X1 U2589 ( .A1(n516), .A2(n4044), .ZN(n4049) );
  AND2_X1 U2590 ( .A1(n2776), .A2(n2403), .ZN(n2480) );
  INV_X1 U2591 ( .A(n4055), .ZN(n4036) );
  NOR2_X1 U2592 ( .A1(IR_CU_27), .A2(IR_CU_26), .ZN(n4055) );
  INV_X1 U2593 ( .A(n3131), .ZN(n3195) );
  AND3_X1 U2594 ( .A1(\DataP/opcode_W[2] ), .A2(\DataP/opcode_W[4] ), .A3(
        n2401), .ZN(n2483) );
  INV_X1 U2595 ( .A(n4188), .ZN(n491) );
  INV_X1 U2596 ( .A(n4187), .ZN(n492) );
  INV_X1 U2597 ( .A(n4156), .ZN(n4148) );
  NAND2_X1 U2598 ( .A1(n516), .A2(n1960), .ZN(n3994) );
  BUF_X1 U2599 ( .A(n3900), .Z(n3227) );
  AND3_X1 U2600 ( .A1(n3409), .A2(n3886), .A3(n3408), .ZN(n3880) );
  INV_X1 U2601 ( .A(n3892), .ZN(n3877) );
  INV_X1 U2602 ( .A(n4186), .ZN(n493) );
  INV_X1 U2603 ( .A(n4185), .ZN(n494) );
  INV_X1 U2604 ( .A(n4189), .ZN(n490) );
  NOR2_X1 U2605 ( .A1(n486), .A2(n4149), .ZN(\DataP/add_S2[1] ) );
  NOR2_X1 U2606 ( .A1(n487), .A2(n4149), .ZN(\DataP/add_S2[2] ) );
  NOR2_X1 U2607 ( .A1(n488), .A2(n4149), .ZN(\DataP/add_S2[3] ) );
  NOR2_X1 U2608 ( .A1(n489), .A2(n4149), .ZN(\DataP/add_S2[4] ) );
  NOR2_X1 U2609 ( .A1(n485), .A2(n4149), .ZN(\DataP/add_S2[0] ) );
  INV_X1 U2610 ( .A(n4151), .ZN(n4052) );
  NOR3_X1 U2611 ( .A1(n3994), .A2(n4155), .A3(n4036), .ZN(n4153) );
  NOR2_X1 U2612 ( .A1(n3994), .A2(n2374), .ZN(n16) );
  BUF_X1 U2613 ( .A(n3904), .Z(n3228) );
  OR2_X1 U2614 ( .A1(n2773), .A2(n2471), .ZN(n3312) );
  AND4_X1 U2615 ( .A1(n3249), .A2(n1638), .A3(n528), .A4(n1637), .ZN(n2406) );
  NOR2_X1 U2616 ( .A1(n504), .A2(n497), .ZN(n4166) );
  OR2_X1 U2617 ( .A1(n4101), .A2(ALU_OPCODE_i[0]), .ZN(n4184) );
  AND2_X2 U2618 ( .A1(n3638), .A2(n3637), .ZN(n3680) );
  AND2_X1 U2619 ( .A1(BR_EN_i), .A2(n4102), .ZN(n3908) );
  NOR2_X1 U2620 ( .A1(ALU_OPCODE_i[3]), .A2(ALU_OPCODE_i[0]), .ZN(n3561) );
  BUF_X1 U2621 ( .A(n4222), .Z(n3232) );
  NOR2_X1 U2622 ( .A1(n3231), .A2(n3235), .ZN(n4222) );
  INV_X1 U2623 ( .A(Rst), .ZN(n3236) );
  INV_X1 U2624 ( .A(Rst), .ZN(n3235) );
  INV_X1 U2625 ( .A(\DataP/npc_mux_sel ), .ZN(n3233) );
  BUF_X1 U2626 ( .A(n4144), .Z(n3229) );
  NOR2_X1 U2627 ( .A1(\WB_MUX_SEL_i[1] ), .A2(n294), .ZN(n4144) );
  INV_X1 U2628 ( .A(n4165), .ZN(n4181) );
  NAND2_X2 U2629 ( .A1(n1586), .A2(n3310), .ZN(\DataP/alu_b_in[3] ) );
  OR2_X2 U2630 ( .A1(n3392), .A2(n3391), .ZN(\DataP/alu_a_in[14] ) );
  INV_X2 U2631 ( .A(n3212), .ZN(n3210) );
  BUF_X2 U2632 ( .A(n3547), .Z(n3221) );
  NOR4_X1 U2633 ( .A1(n443), .A2(ALU_OPCODE_i[3]), .A3(ALU_OPCODE_i[2]), .A4(
        ALU_OPCODE_i[1]), .ZN(n4102) );
  INV_X2 U2634 ( .A(n3891), .ZN(n3894) );
  INV_X2 U2635 ( .A(\DataP/alu_b_in[2] ), .ZN(n3052) );
  OR2_X2 U2636 ( .A1(n3371), .A2(n3370), .ZN(\DataP/alu_a_in[23] ) );
  OR2_X2 U2637 ( .A1(n3374), .A2(n3373), .ZN(\DataP/alu_a_in[22] ) );
  OR2_X2 U2638 ( .A1(n3388), .A2(n3387), .ZN(\DataP/alu_a_in[16] ) );
  OR2_X2 U2639 ( .A1(n3299), .A2(n3298), .ZN(\DataP/alu_a_in[7] ) );
  OR2_X2 U2640 ( .A1(n3337), .A2(n3336), .ZN(\DataP/alu_a_in[4] ) );
  OR2_X2 U2641 ( .A1(n3346), .A2(n3345), .ZN(\DataP/alu_a_in[8] ) );
  OR2_X2 U2642 ( .A1(n3395), .A2(n3394), .ZN(\DataP/alu_a_in[13] ) );
  OR2_X2 U2643 ( .A1(n3389), .A2(n2693), .ZN(\DataP/alu_a_in[15] ) );
  BUF_X2 U2644 ( .A(n2088), .Z(n3226) );
  OR2_X2 U2645 ( .A1(n3353), .A2(n3352), .ZN(\DataP/alu_a_in[30] ) );
  BUF_X2 U2646 ( .A(n2088), .Z(n3224) );
  BUF_X2 U2647 ( .A(n2088), .Z(n3225) );
  BUF_X2 U2648 ( .A(n3547), .Z(n3220) );
  INV_X2 U2649 ( .A(n2072), .ZN(n3208) );
  AOI211_X1 U2650 ( .C1(n4183), .C2(n3907), .A(n4182), .B(n3906), .ZN(
        \DataP/right_br ) );
  AND2_X1 U2651 ( .A1(n4184), .A2(n1905), .ZN(n3906) );
  NAND2_X1 U2652 ( .A1(n3435), .A2(ALU_OPCODE_i[0]), .ZN(n3907) );
  INV_X1 U2653 ( .A(\DataP/add_S2[3] ), .ZN(n2767) );
  INV_X1 U2654 ( .A(\DataP/add_S2[1] ), .ZN(n2770) );
  AOI211_X1 U2655 ( .C1(n3877), .C2(\DataP/ALU_C/shifter/N83 ), .A(n3584), .B(
        n3583), .ZN(n358) );
  AND2_X1 U2656 ( .A1(\DataP/ALU_C/shifter/N51 ), .A2(n3227), .ZN(n3583) );
  OAI211_X1 U2657 ( .C1(n3880), .C2(n3582), .A(n3581), .B(n3580), .ZN(n3584)
         );
  AOI21_X1 U2658 ( .B1(n2130), .B2(n3579), .A(n3578), .ZN(n3580) );
  NAND2_X1 U2659 ( .A1(\DataP/ALU_C/shifter/N19 ), .A2(n3904), .ZN(n3581) );
  INV_X1 U2660 ( .A(n2827), .ZN(n2908) );
  NAND2_X1 U2661 ( .A1(n1622), .A2(n1754), .ZN(n3576) );
  AOI211_X1 U2662 ( .C1(n3877), .C2(\DataP/ALU_C/shifter/N84 ), .A(n3596), .B(
        n3595), .ZN(n357) );
  OAI211_X1 U2663 ( .C1(n3880), .C2(n3594), .A(n3593), .B(n3592), .ZN(n3595)
         );
  AOI21_X1 U2664 ( .B1(n2130), .B2(n3591), .A(n3590), .ZN(n3592) );
  OAI22_X1 U2665 ( .A1(n1719), .A2(n3589), .B1(n3052), .B2(n3891), .ZN(n3590)
         );
  AOI21_X1 U2666 ( .B1(\DataP/alu_b_in[2] ), .B2(n3890), .A(n3894), .ZN(n3589)
         );
  NAND2_X1 U2667 ( .A1(\DataP/ALU_C/shifter/N20 ), .A2(n3228), .ZN(n3593) );
  INV_X1 U2668 ( .A(n2884), .ZN(n2909) );
  NAND2_X1 U2669 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  AND2_X1 U2670 ( .A1(\DataP/ALU_C/shifter/N52 ), .A2(n3227), .ZN(n3596) );
  INV_X1 U2671 ( .A(\DataP/add_S2[0] ), .ZN(n2768) );
  INV_X1 U2672 ( .A(\DataP/add_S2[4] ), .ZN(n2769) );
  OAI22_X1 U2673 ( .A1(n356), .A2(n4111), .B1(n4219), .B2(n4110), .ZN(
        \DataP/PC_reg/N5 ) );
  AOI21_X1 U2674 ( .B1(n2101), .B2(n3891), .A(n3856), .ZN(n3846) );
  OAI211_X1 U2675 ( .C1(n1644), .C2(n1662), .A(n2218), .B(n2129), .ZN(n3847)
         );
  INV_X1 U2676 ( .A(n2895), .ZN(n2910) );
  INV_X1 U2677 ( .A(n2897), .ZN(n2912) );
  OAI22_X1 U2678 ( .A1(n355), .A2(n4111), .B1(n4218), .B2(n4110), .ZN(
        \DataP/PC_reg/N6 ) );
  OAI21_X1 U2679 ( .B1(n3851), .B2(n2102), .A(n3891), .ZN(n3852) );
  INV_X1 U2680 ( .A(n2896), .ZN(n2911) );
  OAI22_X1 U2681 ( .A1(n353), .A2(n4111), .B1(n4216), .B2(n4110), .ZN(
        \DataP/PC_reg/N8 ) );
  AOI211_X1 U2682 ( .C1(n3857), .C2(n3891), .A(n1748), .B(n3856), .ZN(n3858)
         );
  OAI22_X1 U2683 ( .A1(n345), .A2(n4111), .B1(n4214), .B2(n4110), .ZN(
        \DataP/PC_reg/N10 ) );
  AOI21_X1 U2684 ( .B1(n3841), .B2(n2130), .A(n3894), .ZN(n3840) );
  INV_X1 U2685 ( .A(n3838), .ZN(n3856) );
  NOR2_X1 U2686 ( .A1(n2130), .A2(n3894), .ZN(n3839) );
  INV_X1 U2687 ( .A(n2900), .ZN(n2914) );
  AOI22_X1 U2688 ( .A1(n3436), .A2(n2166), .B1(n3894), .B2(n2207), .ZN(n3437)
         );
  OAI21_X1 U2689 ( .B1(n2099), .B2(n3851), .A(n3891), .ZN(n3436) );
  INV_X1 U2690 ( .A(n2901), .ZN(n2915) );
  INV_X1 U2691 ( .A(n3835), .ZN(n3428) );
  OAI21_X1 U2692 ( .B1(n2366), .B2(n3851), .A(n3891), .ZN(n3612) );
  INV_X1 U2693 ( .A(n2899), .ZN(n2913) );
  INV_X1 U2694 ( .A(n1655), .ZN(n3610) );
  AOI21_X1 U2695 ( .B1(n3607), .B2(n2156), .A(n3605), .ZN(n3854) );
  INV_X1 U2696 ( .A(n2215), .ZN(n3605) );
  OAI21_X1 U2697 ( .B1(n3850), .B2(n3600), .A(n3599), .ZN(n3607) );
  INV_X1 U2698 ( .A(n3598), .ZN(n3600) );
  NAND2_X1 U2699 ( .A1(n2218), .A2(n3597), .ZN(n3850) );
  AOI22_X1 U2700 ( .A1(n3452), .A2(n2165), .B1(n3894), .B2(
        \DataP/alu_a_in[10] ), .ZN(n3453) );
  OAI21_X1 U2701 ( .B1(n3451), .B2(n3851), .A(n3891), .ZN(n3452) );
  INV_X1 U2702 ( .A(n2863), .ZN(n2902) );
  INV_X1 U2703 ( .A(n3484), .ZN(n3450) );
  INV_X1 U2704 ( .A(n2875), .ZN(n2904) );
  NAND2_X1 U2705 ( .A1(\DataP/alu_a_in[12] ), .A2(n2655), .ZN(n3492) );
  NOR2_X1 U2706 ( .A1(n1573), .A2(n3851), .ZN(n2655) );
  OAI21_X1 U2707 ( .B1(\DataP/alu_a_in[12] ), .B2(\lt_x_135/B[12] ), .A(n3894), 
        .ZN(n3493) );
  NAND2_X1 U2708 ( .A1(\DataP/ALU_C/shifter/N29 ), .A2(n3228), .ZN(n3471) );
  INV_X1 U2709 ( .A(n2868), .ZN(n2903) );
  AOI21_X1 U2710 ( .B1(n3540), .B2(n2130), .A(n3470), .ZN(n3472) );
  OAI22_X1 U2711 ( .A1(n3469), .A2(n3468), .B1(n3467), .B2(n3891), .ZN(n3470)
         );
  AOI21_X1 U2712 ( .B1(n2200), .B2(n3890), .A(n3894), .ZN(n3469) );
  AOI22_X1 U2713 ( .A1(n3227), .A2(\DataP/ALU_C/shifter/N61 ), .B1(
        \DataP/ALU_C/shifter/N93 ), .B2(n3877), .ZN(n3473) );
  NAND2_X1 U2714 ( .A1(n3466), .A2(n2129), .ZN(n3474) );
  XNOR2_X1 U2715 ( .A(n3465), .B(n3488), .ZN(n3466) );
  OAI21_X1 U2716 ( .B1(n3458), .B2(n3489), .A(n3484), .ZN(n3465) );
  NAND2_X1 U2717 ( .A1(n3446), .A2(n3445), .ZN(n3458) );
  NAND2_X1 U2718 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  NAND2_X1 U2719 ( .A1(n3483), .A2(n3835), .ZN(n3444) );
  NAND2_X1 U2720 ( .A1(n3837), .A2(n2205), .ZN(n3446) );
  NAND2_X1 U2721 ( .A1(n2084), .A2(n3482), .ZN(n3837) );
  OAI22_X1 U2722 ( .A1(n333), .A2(n4111), .B1(n4110), .B2(n4209), .ZN(
        \DataP/PC_reg/N15 ) );
  INV_X1 U2723 ( .A(\DataP/npc[13] ), .ZN(n4209) );
  OAI21_X1 U2724 ( .B1(\DataP/alu_a_in[13] ), .B2(n2141), .A(n3894), .ZN(n3871) );
  INV_X1 U2725 ( .A(n2882), .ZN(n2905) );
  NAND2_X1 U2726 ( .A1(n1710), .A2(n3863), .ZN(n3866) );
  OAI22_X1 U2727 ( .A1(n326), .A2(n4111), .B1(n4110), .B2(n4206), .ZN(
        \DataP/PC_reg/N18 ) );
  INV_X1 U2728 ( .A(\DataP/npc[16] ), .ZN(n4206) );
  AOI21_X1 U2729 ( .B1(n3737), .B2(n2129), .A(n3736), .ZN(n326) );
  NAND2_X1 U2730 ( .A1(\DataP/ALU_C/shifter/N34 ), .A2(n3228), .ZN(n3733) );
  AOI21_X1 U2731 ( .B1(\DataP/ALU_C/shifter/N66 ), .B2(n3227), .A(n3732), .ZN(
        n3735) );
  OAI22_X1 U2732 ( .A1(n319), .A2(n4111), .B1(n4110), .B2(n4203), .ZN(
        \DataP/PC_reg/N21 ) );
  INV_X1 U2733 ( .A(\DataP/npc[19] ), .ZN(n4203) );
  AOI21_X1 U2734 ( .B1(n3658), .B2(n2129), .A(n3657), .ZN(n319) );
  NAND2_X1 U2735 ( .A1(\DataP/ALU_C/shifter/N37 ), .A2(n3904), .ZN(n3654) );
  AOI21_X1 U2736 ( .B1(\DataP/ALU_C/shifter/N69 ), .B2(n3900), .A(n3653), .ZN(
        n3655) );
  OAI211_X1 U2737 ( .C1(n4106), .C2(n3897), .A(n3652), .B(n3651), .ZN(n3653)
         );
  NAND2_X1 U2738 ( .A1(\DataP/alu_a_in[19] ), .A2(n3894), .ZN(n3651) );
  OAI211_X1 U2739 ( .C1(\DataP/alu_a_in[19] ), .C2(n3894), .A(n1722), .B(n3838), .ZN(n3652) );
  NAND2_X1 U2740 ( .A1(\DataP/ALU_C/shifter/N101 ), .A2(n3877), .ZN(n3656) );
  OAI22_X1 U2741 ( .A1(n322), .A2(n4111), .B1(n4110), .B2(n4204), .ZN(
        \DataP/PC_reg/N20 ) );
  INV_X1 U2742 ( .A(\DataP/npc[18] ), .ZN(n4204) );
  INV_X1 U2743 ( .A(n3752), .ZN(n322) );
  OAI211_X1 U2744 ( .C1(n3751), .C2(n3880), .A(n3750), .B(n3749), .ZN(n3752)
         );
  NAND2_X1 U2745 ( .A1(\DataP/ALU_C/shifter/N100 ), .A2(n3877), .ZN(n3749) );
  AOI21_X1 U2746 ( .B1(n3904), .B2(\DataP/ALU_C/shifter/N36 ), .A(n3748), .ZN(
        n3750) );
  NAND3_X1 U2747 ( .A1(n2724), .A2(n3635), .A3(n2378), .ZN(n2673) );
  OAI22_X1 U2748 ( .A1(n323), .A2(n4111), .B1(n4110), .B2(n4205), .ZN(
        \DataP/PC_reg/N19 ) );
  INV_X1 U2749 ( .A(\DataP/npc[17] ), .ZN(n4205) );
  AOI21_X1 U2750 ( .B1(\DataP/ALU_C/shifter/N67 ), .B2(n3227), .A(n3742), .ZN(
        n3744) );
  OAI211_X1 U2751 ( .C1(n3741), .C2(n3897), .A(n3740), .B(n3739), .ZN(n3742)
         );
  OAI211_X1 U2752 ( .C1(n1751), .C2(n3894), .A(\DataP/alu_b_in[17] ), .B(n3838), .ZN(n3739) );
  NAND2_X1 U2753 ( .A1(n1751), .A2(n3894), .ZN(n3740) );
  NAND2_X1 U2754 ( .A1(\DataP/ALU_C/shifter/N99 ), .A2(n3877), .ZN(n3745) );
  NAND2_X1 U2755 ( .A1(n2078), .A2(n3680), .ZN(n3729) );
  OAI22_X1 U2756 ( .A1(n311), .A2(n4111), .B1(n4110), .B2(n4200), .ZN(
        \DataP/PC_reg/N24 ) );
  INV_X1 U2757 ( .A(\DataP/npc[22] ), .ZN(n4200) );
  AOI21_X1 U2758 ( .B1(n3787), .B2(n2129), .A(n3786), .ZN(n311) );
  OAI21_X1 U2759 ( .B1(n3892), .B2(n3785), .A(n3784), .ZN(n3786) );
  AOI21_X1 U2760 ( .B1(n3904), .B2(\DataP/ALU_C/shifter/N40 ), .A(n3783), .ZN(
        n3784) );
  OAI211_X1 U2761 ( .C1(n3897), .C2(n3782), .A(n3781), .B(n3780), .ZN(n3783)
         );
  AOI22_X1 U2762 ( .A1(n3779), .A2(\DataP/alu_b_in[22] ), .B1(n3894), .B2(
        \DataP/alu_a_in[22] ), .ZN(n3780) );
  OAI21_X1 U2763 ( .B1(n3778), .B2(n3851), .A(n3891), .ZN(n3779) );
  NAND2_X1 U2764 ( .A1(\DataP/ALU_C/shifter/N72 ), .A2(n3227), .ZN(n3781) );
  INV_X1 U2765 ( .A(\DataP/ALU_C/shifter/N104 ), .ZN(n3785) );
  XNOR2_X1 U2766 ( .A(n3777), .B(n3776), .ZN(n3787) );
  INV_X1 U2767 ( .A(\DataP/npc[21] ), .ZN(n4201) );
  OAI21_X1 U2768 ( .B1(n3892), .B2(n3774), .A(n3773), .ZN(n3775) );
  AOI21_X1 U2769 ( .B1(n3904), .B2(\DataP/ALU_C/shifter/N39 ), .A(n3772), .ZN(
        n3773) );
  OAI211_X1 U2770 ( .C1(n3897), .C2(n3771), .A(n3770), .B(n3769), .ZN(n3772)
         );
  AOI22_X1 U2771 ( .A1(n3768), .A2(n2152), .B1(n3894), .B2(
        \DataP/alu_a_in[21] ), .ZN(n3769) );
  OAI21_X1 U2772 ( .B1(n2111), .B2(n3851), .A(n3891), .ZN(n3768) );
  NAND2_X1 U2773 ( .A1(\DataP/ALU_C/shifter/N71 ), .A2(n3227), .ZN(n3770) );
  INV_X1 U2774 ( .A(\DataP/ALU_C/shifter/N103 ), .ZN(n3774) );
  INV_X1 U2775 ( .A(n1588), .ZN(n3765) );
  OAI22_X1 U2776 ( .A1(n317), .A2(n4111), .B1(n4110), .B2(n4202), .ZN(
        \DataP/PC_reg/N22 ) );
  INV_X1 U2777 ( .A(\DataP/npc[20] ), .ZN(n4202) );
  AOI21_X1 U2778 ( .B1(n3761), .B2(n2129), .A(n3760), .ZN(n317) );
  NAND2_X1 U2779 ( .A1(\DataP/ALU_C/shifter/N38 ), .A2(n3228), .ZN(n3757) );
  AOI21_X1 U2780 ( .B1(\DataP/ALU_C/shifter/N70 ), .B2(n3227), .A(n3756), .ZN(
        n3758) );
  OAI211_X1 U2781 ( .C1(n4107), .C2(n3897), .A(n3755), .B(n3754), .ZN(n3756)
         );
  NAND2_X1 U2782 ( .A1(\DataP/alu_a_in[20] ), .A2(n3894), .ZN(n3754) );
  OAI211_X1 U2783 ( .C1(\DataP/alu_a_in[20] ), .C2(n3894), .A(
        \DataP/alu_b_in[20] ), .B(n3838), .ZN(n3755) );
  NAND2_X1 U2784 ( .A1(\DataP/ALU_C/shifter/N102 ), .A2(n3877), .ZN(n3759) );
  OAI22_X1 U2785 ( .A1(n308), .A2(n4111), .B1(n4110), .B2(n4198), .ZN(
        \DataP/PC_reg/N26 ) );
  INV_X1 U2786 ( .A(\DataP/npc[24] ), .ZN(n4198) );
  AOI21_X1 U2787 ( .B1(n3796), .B2(n2129), .A(n3795), .ZN(n308) );
  NAND2_X1 U2788 ( .A1(\DataP/ALU_C/shifter/N42 ), .A2(n3228), .ZN(n3792) );
  AOI21_X1 U2789 ( .B1(\DataP/ALU_C/shifter/N74 ), .B2(n3227), .A(n3791), .ZN(
        n3793) );
  OAI211_X1 U2790 ( .C1(n4109), .C2(n3897), .A(n3790), .B(n3789), .ZN(n3791)
         );
  NAND2_X1 U2791 ( .A1(\DataP/alu_a_in[24] ), .A2(n3894), .ZN(n3789) );
  OAI211_X1 U2792 ( .C1(\DataP/alu_a_in[24] ), .C2(n3894), .A(
        \DataP/alu_b_in[24] ), .B(n3838), .ZN(n3790) );
  NAND2_X1 U2793 ( .A1(\DataP/ALU_C/shifter/N106 ), .A2(n3877), .ZN(n3794) );
  INV_X1 U2794 ( .A(n3127), .ZN(n3197) );
  AND3_X1 U2795 ( .A1(n2555), .A2(n2556), .A3(n2558), .ZN(n297) );
  OR2_X1 U2796 ( .A1(n2752), .A2(n2083), .ZN(n2555) );
  AOI21_X1 U2797 ( .B1(n2654), .B2(n2129), .A(n3824), .ZN(n300) );
  INV_X1 U2798 ( .A(\DataP/npc[26] ), .ZN(n4196) );
  NAND2_X1 U2799 ( .A1(\DataP/ALU_C/shifter/N108 ), .A2(n3877), .ZN(n3812) );
  INV_X1 U2800 ( .A(n3133), .ZN(\DataP/ALU_C/shifter/N108 ) );
  AOI21_X1 U2801 ( .B1(\DataP/ALU_C/shifter/N76 ), .B2(n3227), .A(n3811), .ZN(
        n3813) );
  OAI211_X1 U2802 ( .C1(n3810), .C2(n3897), .A(n3809), .B(n3808), .ZN(n3811)
         );
  NAND2_X1 U2803 ( .A1(\DataP/alu_a_in[26] ), .A2(n3894), .ZN(n3808) );
  OAI211_X1 U2804 ( .C1(\DataP/alu_a_in[26] ), .C2(n3894), .A(
        \DataP/alu_b_in[26] ), .B(n3838), .ZN(n3809) );
  NAND2_X1 U2805 ( .A1(n3719), .A2(n2584), .ZN(n3807) );
  OAI211_X1 U2806 ( .C1(n2216), .C2(n2756), .A(n2574), .B(n2482), .ZN(n2774)
         );
  INV_X1 U2807 ( .A(n2756), .ZN(n2575) );
  INV_X1 U2808 ( .A(\DataP/npc[31] ), .ZN(n4191) );
  NAND2_X1 U2809 ( .A1(n1721), .A2(n2754), .ZN(n2753) );
  OAI21_X1 U2810 ( .B1(n3905), .B2(n3902), .A(n3901), .ZN(n3903) );
  AOI21_X1 U2811 ( .B1(\DataP/ALU_C/shifter/N81 ), .B2(n3227), .A(n3899), .ZN(
        n3901) );
  OAI21_X1 U2812 ( .B1(n3898), .B2(n3897), .A(n3896), .ZN(n3899) );
  AOI22_X1 U2813 ( .A1(\DataP/alu_a_in[31] ), .A2(n3895), .B1(n3894), .B2(
        \DataP/alu_b_in[31] ), .ZN(n3896) );
  NAND2_X1 U2814 ( .A1(\DataP/alu_b_in[31] ), .A2(n3890), .ZN(n3893) );
  NOR2_X1 U2815 ( .A1(n3905), .A2(n2750), .ZN(n2749) );
  NOR2_X1 U2816 ( .A1(n2754), .A2(n3905), .ZN(n2751) );
  NAND2_X1 U2817 ( .A1(n3888), .A2(n2129), .ZN(n3905) );
  INV_X1 U2818 ( .A(n3889), .ZN(n3888) );
  AOI21_X1 U2819 ( .B1(n2663), .B2(n2129), .A(n3704), .ZN(n301) );
  INV_X1 U2820 ( .A(\DataP/npc[23] ), .ZN(n4199) );
  OAI211_X1 U2821 ( .C1(n3678), .C2(n3892), .A(n3677), .B(n3676), .ZN(n3679)
         );
  NAND2_X1 U2822 ( .A1(\DataP/ALU_C/shifter/N41 ), .A2(n3228), .ZN(n3676) );
  AOI21_X1 U2823 ( .B1(\DataP/ALU_C/shifter/N73 ), .B2(n3227), .A(n3675), .ZN(
        n3677) );
  OAI211_X1 U2824 ( .C1(n4108), .C2(n3897), .A(n3674), .B(n3673), .ZN(n3675)
         );
  NAND2_X1 U2825 ( .A1(\DataP/alu_a_in[23] ), .A2(n3894), .ZN(n3673) );
  OAI211_X1 U2826 ( .C1(\DataP/alu_a_in[23] ), .C2(n3894), .A(
        \DataP/alu_b_in[23] ), .B(n3838), .ZN(n3674) );
  INV_X1 U2827 ( .A(\DataP/ALU_C/shifter/N105 ), .ZN(n3678) );
  INV_X1 U2828 ( .A(n3125), .ZN(n3196) );
  INV_X1 U2829 ( .A(n1717), .ZN(n3672) );
  NAND2_X1 U2830 ( .A1(n2763), .A2(n2761), .ZN(n2760) );
  NOR2_X1 U2831 ( .A1(n3680), .A2(n2762), .ZN(n2761) );
  INV_X1 U2832 ( .A(n3683), .ZN(n2762) );
  INV_X1 U2833 ( .A(\DataP/npc[28] ), .ZN(n4194) );
  OAI211_X1 U2834 ( .C1(n3892), .C2(n3137), .A(n3823), .B(n3822), .ZN(n3824)
         );
  AOI21_X1 U2835 ( .B1(\DataP/ALU_C/shifter/N78 ), .B2(n3227), .A(n3821), .ZN(
        n3822) );
  OAI21_X1 U2836 ( .B1(n3897), .B2(n3820), .A(n3819), .ZN(n3821) );
  AOI22_X1 U2837 ( .A1(n3818), .A2(\DataP/alu_b_in[28] ), .B1(n3894), .B2(
        \DataP/alu_a_in[28] ), .ZN(n3819) );
  OAI21_X1 U2838 ( .B1(n3817), .B2(n3851), .A(n3891), .ZN(n3818) );
  NAND2_X1 U2839 ( .A1(\DataP/ALU_C/shifter/N46 ), .A2(n3228), .ZN(n3823) );
  INV_X1 U2840 ( .A(n3798), .ZN(n2747) );
  OAI22_X1 U2841 ( .A1(n304), .A2(n4111), .B1(n4110), .B2(n4197), .ZN(
        \DataP/PC_reg/N27 ) );
  INV_X1 U2842 ( .A(\DataP/npc[25] ), .ZN(n4197) );
  AOI21_X1 U2843 ( .B1(n3806), .B2(n2129), .A(n3805), .ZN(n304) );
  AOI21_X1 U2844 ( .B1(\DataP/ALU_C/shifter/N75 ), .B2(n3227), .A(n3801), .ZN(
        n3802) );
  NAND2_X1 U2845 ( .A1(\DataP/ALU_C/shifter/N43 ), .A2(n3228), .ZN(n3803) );
  NAND2_X1 U2846 ( .A1(\DataP/ALU_C/shifter/N107 ), .A2(n3877), .ZN(n3804) );
  INV_X1 U2847 ( .A(n3130), .ZN(n3198) );
  OAI22_X1 U2848 ( .A1(n330), .A2(n4111), .B1(n4110), .B2(n4207), .ZN(
        \DataP/PC_reg/N17 ) );
  INV_X1 U2849 ( .A(\DataP/npc[15] ), .ZN(n4207) );
  AOI21_X1 U2850 ( .B1(n2689), .B2(n2129), .A(n2688), .ZN(n330) );
  NAND2_X1 U2851 ( .A1(n3626), .A2(n3627), .ZN(n2688) );
  AOI21_X1 U2852 ( .B1(\DataP/ALU_C/shifter/N65 ), .B2(n3900), .A(n3625), .ZN(
        n3627) );
  OAI211_X1 U2853 ( .C1(n3624), .C2(n3891), .A(n3623), .B(n3622), .ZN(n3625)
         );
  OAI211_X1 U2854 ( .C1(\DataP/alu_a_in[15] ), .C2(n3894), .A(
        \DataP/alu_b_in[15] ), .B(n3838), .ZN(n3622) );
  NAND2_X1 U2855 ( .A1(n3621), .A2(n2130), .ZN(n3623) );
  AOI22_X1 U2856 ( .A1(\DataP/ALU_C/shifter/N33 ), .A2(n3228), .B1(n3877), 
        .B2(\DataP/ALU_C/shifter/N97 ), .ZN(n3626) );
  INV_X1 U2857 ( .A(n2894), .ZN(n2907) );
  INV_X1 U2858 ( .A(\DataP/npc[29] ), .ZN(n4193) );
  OAI211_X1 U2859 ( .C1(n3892), .C2(n3139), .A(n3832), .B(n3831), .ZN(n3833)
         );
  AOI21_X1 U2860 ( .B1(\DataP/ALU_C/shifter/N79 ), .B2(n3227), .A(n3830), .ZN(
        n3831) );
  OAI21_X1 U2861 ( .B1(n3897), .B2(n3829), .A(n3828), .ZN(n3830) );
  AOI22_X1 U2862 ( .A1(n3827), .A2(\DataP/alu_b_in[29] ), .B1(n3894), .B2(
        \DataP/alu_a_in[29] ), .ZN(n3828) );
  OAI21_X1 U2863 ( .B1(n2365), .B2(n3851), .A(n3891), .ZN(n3827) );
  NAND2_X1 U2864 ( .A1(\DataP/ALU_C/shifter/N47 ), .A2(n3904), .ZN(n3832) );
  AND2_X1 U2865 ( .A1(n2766), .A2(n2748), .ZN(n2717) );
  AOI21_X1 U2866 ( .B1(n2756), .B2(n2131), .A(n2474), .ZN(n2707) );
  INV_X1 U2867 ( .A(\DataP/npc[30] ), .ZN(n4192) );
  NAND2_X1 U2868 ( .A1(\DataP/alu_a_in[30] ), .A2(n3894), .ZN(n3705) );
  OAI211_X1 U2869 ( .C1(\DataP/alu_a_in[30] ), .C2(n3894), .A(
        \DataP/alu_b_in[30] ), .B(n3838), .ZN(n3706) );
  NAND2_X1 U2870 ( .A1(n3891), .A2(n3851), .ZN(n3838) );
  OR2_X1 U2871 ( .A1(n3880), .A2(n4111), .ZN(n2708) );
  AOI21_X1 U2872 ( .B1(n3713), .B2(n1548), .A(n3788), .ZN(n3717) );
  AND2_X1 U2873 ( .A1(n3715), .A2(n1717), .ZN(n2726) );
  NOR2_X1 U2874 ( .A1(n3725), .A2(n3798), .ZN(n2748) );
  NAND2_X1 U2875 ( .A1(n3711), .A2(\DataP/alu_a_in[30] ), .ZN(n3884) );
  INV_X1 U2876 ( .A(n3710), .ZN(n3711) );
  NAND2_X1 U2877 ( .A1(n3710), .A2(n2364), .ZN(n3902) );
  OAI21_X1 U2878 ( .B1(n2566), .B2(n2535), .A(n2565), .ZN(n3710) );
  NAND2_X1 U2879 ( .A1(n2614), .A2(n2535), .ZN(n2565) );
  XNOR2_X1 U2880 ( .A(n2567), .B(\DataP/alu_b_in[30] ), .ZN(n2566) );
  NOR2_X1 U2881 ( .A1(n3722), .A2(n2381), .ZN(n2567) );
  INV_X1 U2882 ( .A(n3728), .ZN(n3727) );
  NOR2_X1 U2883 ( .A1(n3724), .A2(\DataP/alu_a_in[28] ), .ZN(n2765) );
  INV_X1 U2884 ( .A(n3816), .ZN(n3724) );
  NOR2_X1 U2885 ( .A1(n3816), .A2(n3817), .ZN(n3725) );
  INV_X1 U2886 ( .A(\DataP/alu_a_in[28] ), .ZN(n3817) );
  XNOR2_X1 U2887 ( .A(n3722), .B(\DataP/alu_b_in[28] ), .ZN(n3723) );
  NAND2_X1 U2888 ( .A1(n3709), .A2(n3726), .ZN(n3722) );
  NOR2_X1 U2889 ( .A1(n3708), .A2(\DataP/alu_b_in[27] ), .ZN(n3726) );
  AOI21_X1 U2890 ( .B1(n3704), .B2(n2131), .A(n2592), .ZN(n2591) );
  NOR2_X1 U2891 ( .A1(n4110), .A2(n4195), .ZN(n2592) );
  INV_X1 U2892 ( .A(\DataP/npc[27] ), .ZN(n4195) );
  OAI211_X1 U2893 ( .C1(n3892), .C2(n3135), .A(n3703), .B(n3702), .ZN(n3704)
         );
  AOI21_X1 U2894 ( .B1(\DataP/ALU_C/shifter/N77 ), .B2(n3227), .A(n3701), .ZN(
        n3702) );
  OAI21_X1 U2895 ( .B1(n3897), .B2(n3700), .A(n3699), .ZN(n3701) );
  AOI22_X1 U2896 ( .A1(n3698), .A2(\DataP/alu_b_in[27] ), .B1(n3894), .B2(
        \DataP/alu_a_in[27] ), .ZN(n3699) );
  OAI21_X1 U2897 ( .B1(n3697), .B2(n3851), .A(n3891), .ZN(n3698) );
  NAND2_X1 U2898 ( .A1(\DataP/ALU_C/shifter/N45 ), .A2(n3228), .ZN(n3703) );
  INV_X1 U2899 ( .A(n3708), .ZN(n2703) );
  NAND2_X1 U2900 ( .A1(n2485), .A2(n2127), .ZN(n3708) );
  AND2_X1 U2901 ( .A1(n2588), .A2(n2107), .ZN(n2485) );
  AOI21_X1 U2902 ( .B1(n2389), .B2(n2715), .A(n2706), .ZN(n2705) );
  INV_X1 U2903 ( .A(n3696), .ZN(n2706) );
  OAI21_X1 U2904 ( .B1(n3798), .B2(n2727), .A(n3797), .ZN(n3696) );
  NAND2_X1 U2905 ( .A1(\DataP/alu_b_in[23] ), .A2(n2535), .ZN(n2701) );
  NAND2_X1 U2906 ( .A1(n3692), .A2(n2122), .ZN(n2702) );
  INV_X1 U2907 ( .A(\DataP/alu_a_in[22] ), .ZN(n3778) );
  AND2_X1 U2908 ( .A1(n3683), .A2(n2239), .ZN(n3730) );
  NAND2_X1 U2909 ( .A1(n3646), .A2(n3645), .ZN(n3683) );
  INV_X1 U2910 ( .A(\DataP/alu_a_in[16] ), .ZN(n3645) );
  NAND2_X1 U2911 ( .A1(n3763), .A2(n1588), .ZN(n2606) );
  XNOR2_X1 U2912 ( .A(n1574), .B(\DataP/alu_b_in[24] ), .ZN(n3695) );
  INV_X1 U2913 ( .A(n3668), .ZN(n3692) );
  NAND2_X1 U2914 ( .A1(n2679), .A2(n3886), .ZN(n2676) );
  INV_X1 U2915 ( .A(n2679), .ZN(n2598) );
  AND3_X1 U2916 ( .A1(n2224), .A2(n3714), .A3(n3680), .ZN(n3681) );
  NAND2_X1 U2917 ( .A1(n2402), .A2(n3886), .ZN(n2569) );
  NAND2_X1 U2918 ( .A1(n3663), .A2(n3664), .ZN(n3668) );
  NOR2_X1 U2919 ( .A1(\DataP/alu_a_in[18] ), .A2(n2548), .ZN(n2547) );
  INV_X1 U2920 ( .A(n2757), .ZN(n2548) );
  NAND2_X1 U2921 ( .A1(n2732), .A2(n2731), .ZN(n2730) );
  INV_X1 U2922 ( .A(\DataP/alu_b_in[19] ), .ZN(n2732) );
  OR2_X1 U2923 ( .A1(n2244), .A2(n2486), .ZN(n2733) );
  OR2_X1 U2924 ( .A1(n2135), .A2(n2757), .ZN(n2524) );
  NAND2_X1 U2925 ( .A1(n2546), .A2(n2526), .ZN(n2525) );
  NOR2_X1 U2926 ( .A1(n2135), .A2(n2535), .ZN(n2526) );
  NAND2_X1 U2927 ( .A1(n2301), .A2(n1753), .ZN(n3659) );
  NAND2_X1 U2928 ( .A1(n3616), .A2(n3615), .ZN(n3638) );
  AND2_X1 U2929 ( .A1(\DataP/alu_a_in[15] ), .A2(n2108), .ZN(n3615) );
  NAND2_X1 U2930 ( .A1(n3614), .A2(n2479), .ZN(n2577) );
  INV_X1 U2931 ( .A(\DataP/alu_a_in[15] ), .ZN(n3624) );
  INV_X1 U2932 ( .A(n3616), .ZN(n3614) );
  NAND2_X1 U2933 ( .A1(n3633), .A2(n3632), .ZN(n2724) );
  AND2_X1 U2934 ( .A1(n2647), .A2(n2643), .ZN(n2642) );
  AND2_X1 U2935 ( .A1(n3632), .A2(n1739), .ZN(n2611) );
  INV_X1 U2936 ( .A(n3632), .ZN(n3636) );
  INV_X1 U2937 ( .A(n3630), .ZN(n3868) );
  NAND2_X1 U2938 ( .A1(n3628), .A2(n3865), .ZN(n3861) );
  OAI22_X1 U2939 ( .A1(n332), .A2(n4111), .B1(n4110), .B2(n4208), .ZN(
        \DataP/PC_reg/N16 ) );
  INV_X1 U2940 ( .A(\DataP/npc[14] ), .ZN(n4208) );
  INV_X1 U2941 ( .A(n3882), .ZN(n332) );
  OAI211_X1 U2942 ( .C1(n3881), .C2(n3880), .A(n3879), .B(n3878), .ZN(n3882)
         );
  AOI22_X1 U2943 ( .A1(\DataP/ALU_C/shifter/N32 ), .A2(n3228), .B1(n3877), 
        .B2(\DataP/ALU_C/shifter/N96 ), .ZN(n3878) );
  INV_X1 U2944 ( .A(n2890), .ZN(n2906) );
  AOI21_X1 U2945 ( .B1(\DataP/ALU_C/shifter/N64 ), .B2(n3227), .A(n3876), .ZN(
        n3879) );
  XNOR2_X1 U2946 ( .A(n3874), .B(n3873), .ZN(n3881) );
  AND2_X1 U2947 ( .A1(n3631), .A2(n3632), .ZN(n3873) );
  NOR2_X1 U2948 ( .A1(n2652), .A2(n2650), .ZN(n2649) );
  NOR2_X1 U2949 ( .A1(n2390), .A2(n2108), .ZN(n2650) );
  INV_X1 U2950 ( .A(n2390), .ZN(n2651) );
  INV_X1 U2951 ( .A(n3629), .ZN(n3867) );
  OAI21_X1 U2952 ( .B1(n1713), .B2(n2738), .A(n2393), .ZN(n3630) );
  NAND2_X1 U2953 ( .A1(n2740), .A2(n2128), .ZN(n2737) );
  XNOR2_X1 U2954 ( .A(n3618), .B(n2106), .ZN(n3619) );
  OAI21_X1 U2955 ( .B1(n1597), .B2(n2736), .A(n1726), .ZN(n3863) );
  INV_X1 U2956 ( .A(n2739), .ZN(n2736) );
  INV_X1 U2957 ( .A(n3865), .ZN(n3617) );
  NOR2_X1 U2958 ( .A1(\DataP/alu_b_in[11] ), .A2(\DataP/alu_b_in[10] ), .ZN(
        n3479) );
  AND2_X1 U2959 ( .A1(n3491), .A2(n3490), .ZN(n3628) );
  NAND2_X1 U2960 ( .A1(n1714), .A2(n3463), .ZN(n3491) );
  AND2_X1 U2961 ( .A1(n2200), .A2(n2108), .ZN(n3463) );
  INV_X1 U2962 ( .A(n2200), .ZN(n3467) );
  XNOR2_X1 U2963 ( .A(n3461), .B(n2151), .ZN(n3462) );
  NAND2_X1 U2964 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  NAND2_X1 U2965 ( .A1(n3485), .A2(n3484), .ZN(n3486) );
  NAND2_X1 U2966 ( .A1(n3447), .A2(n3451), .ZN(n3484) );
  INV_X1 U2967 ( .A(\DataP/alu_a_in[10] ), .ZN(n3451) );
  OAI211_X1 U2968 ( .C1(n3426), .C2(n3425), .A(n3424), .B(n3611), .ZN(n3487)
         );
  NAND2_X1 U2969 ( .A1(n3855), .A2(n1655), .ZN(n3424) );
  XNOR2_X1 U2970 ( .A(n3427), .B(\DataP/alu_a_in[7] ), .ZN(n3611) );
  NAND2_X1 U2971 ( .A1(n3608), .A2(n3606), .ZN(n3425) );
  NAND2_X1 U2972 ( .A1(n3422), .A2(\DataP/alu_a_in[5] ), .ZN(n3606) );
  INV_X1 U2973 ( .A(n1747), .ZN(n3422) );
  NAND2_X1 U2974 ( .A1(n3604), .A2(n3599), .ZN(n3419) );
  NAND2_X1 U2975 ( .A1(n3849), .A2(n3418), .ZN(n3599) );
  INV_X1 U2976 ( .A(\DataP/alu_a_in[4] ), .ZN(n3418) );
  INV_X1 U2977 ( .A(n3414), .ZN(n3415) );
  XNOR2_X1 U2978 ( .A(n3412), .B(n1973), .ZN(n3845) );
  AND2_X1 U2979 ( .A1(n3598), .A2(n3597), .ZN(n3420) );
  NAND2_X1 U2980 ( .A1(n1589), .A2(n1973), .ZN(n3597) );
  XNOR2_X1 U2981 ( .A(n3410), .B(\DataP/alu_b_in[3] ), .ZN(n3411) );
  NOR2_X1 U2982 ( .A1(\DataP/alu_b_in[0] ), .A2(\DataP/alu_b_in[1] ), .ZN(
        n3416) );
  NAND2_X1 U2983 ( .A1(n1712), .A2(\DataP/alu_a_in[4] ), .ZN(n3598) );
  NAND2_X1 U2984 ( .A1(n2225), .A2(\DataP/alu_a_in[8] ), .ZN(n3835) );
  NAND2_X1 U2985 ( .A1(n1610), .A2(\DataP/alu_a_in[7] ), .ZN(n3482) );
  INV_X1 U2986 ( .A(n1577), .ZN(n3429) );
  INV_X1 U2987 ( .A(n3310), .ZN(n2659) );
  INV_X1 U2988 ( .A(n3908), .ZN(n3438) );
  AOI21_X1 U2989 ( .B1(n3572), .B2(n2491), .A(n2668), .ZN(n296) );
  OAI21_X1 U2990 ( .B1(n2670), .B2(n2491), .A(n2669), .ZN(n2668) );
  AOI21_X1 U2991 ( .B1(\DataP/ALU_C/shifter/N82 ), .B2(n3877), .A(n3573), .ZN(
        n2669) );
  NAND4_X1 U2992 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3573)
         );
  OAI21_X1 U2993 ( .B1(n3555), .B2(n3894), .A(n3554), .ZN(n3556) );
  NAND2_X1 U2994 ( .A1(n3435), .A2(n3561), .ZN(n3891) );
  AOI21_X1 U2995 ( .B1(n3880), .B2(n3897), .A(n3577), .ZN(n3555) );
  NOR2_X1 U2996 ( .A1(n3237), .A2(ALU_OPCODE_i[1]), .ZN(n3435) );
  NAND2_X1 U2997 ( .A1(ALU_OPCODE_i[2]), .A2(n443), .ZN(n3237) );
  INV_X1 U2998 ( .A(n3562), .ZN(n3432) );
  XNOR2_X1 U2999 ( .A(ALU_OPCODE_i[2]), .B(n4100), .ZN(n3407) );
  NAND2_X1 U3000 ( .A1(n3405), .A2(n3563), .ZN(n3409) );
  OAI21_X1 U3001 ( .B1(n443), .B2(ALU_OPCODE_i[3]), .A(n3562), .ZN(n3405) );
  NAND2_X1 U3002 ( .A1(n1741), .A2(n3890), .ZN(n3557) );
  OR2_X1 U3003 ( .A1(n3434), .A2(n3562), .ZN(n3851) );
  INV_X1 U3004 ( .A(n3433), .ZN(n3434) );
  AND2_X1 U3005 ( .A1(n3406), .A2(ALU_OPCODE_i[1]), .ZN(n3433) );
  NOR2_X1 U3006 ( .A1(ALU_OPCODE_i[2]), .A2(n2491), .ZN(n3406) );
  INV_X1 U3007 ( .A(n3561), .ZN(n3430) );
  NAND2_X1 U3008 ( .A1(\DataP/ALU_C/shifter/N50 ), .A2(n3900), .ZN(n3559) );
  NOR2_X1 U3009 ( .A1(n3562), .A2(n4101), .ZN(n3900) );
  INV_X1 U3010 ( .A(n4101), .ZN(n3431) );
  NOR2_X1 U3011 ( .A1(n3571), .A2(n3570), .ZN(n2671) );
  OAI211_X1 U3012 ( .C1(n3568), .C2(n2391), .A(n3567), .B(n3566), .ZN(n3572)
         );
  OAI21_X1 U3013 ( .B1(n3565), .B2(n3571), .A(n3564), .ZN(n3566) );
  INV_X1 U3014 ( .A(n3570), .ZN(n3564) );
  NOR2_X1 U3015 ( .A1(ALU_OPCODE_i[2]), .A2(ALU_OPCODE_i[1]), .ZN(n3563) );
  INV_X1 U3016 ( .A(\DataP/ALU_C/comp/N50 ), .ZN(n3565) );
  AOI22_X1 U3017 ( .A1(\DataP/ALU_C/comp/N50 ), .A2(n3560), .B1(n3561), .B2(
        n3571), .ZN(n3568) );
  INV_X1 U3018 ( .A(n3569), .ZN(n3571) );
  NAND2_X1 U3019 ( .A1(n2683), .A2(n2682), .ZN(n3560) );
  NAND2_X1 U3020 ( .A1(n3561), .A2(ALU_OPCODE_i[1]), .ZN(n2682) );
  NAND2_X1 U3021 ( .A1(n3569), .A2(n2684), .ZN(n2683) );
  NOR2_X1 U3022 ( .A1(n3562), .A2(ALU_OPCODE_i[1]), .ZN(n2684) );
  NAND2_X1 U3023 ( .A1(n2672), .A2(ALU_OPCODE_i[0]), .ZN(n3562) );
  NAND2_X1 U3024 ( .A1(n4103), .A2(n2741), .ZN(n3569) );
  AND2_X1 U3025 ( .A1(n2742), .A2(n4104), .ZN(n2741) );
  NOR3_X1 U3026 ( .A1(n3511), .A2(n3579), .A3(n3510), .ZN(n4104) );
  NAND4_X1 U3027 ( .A1(n3829), .A2(n3820), .A3(n3700), .A4(n3810), .ZN(n3510)
         );
  XNOR2_X1 U3028 ( .A(\DataP/alu_a_in[26] ), .B(\DataP/alu_b_in[26] ), .ZN(
        n3810) );
  XNOR2_X1 U3029 ( .A(\DataP/alu_a_in[27] ), .B(\DataP/alu_b_in[27] ), .ZN(
        n3700) );
  XNOR2_X1 U3030 ( .A(\DataP/alu_a_in[28] ), .B(\DataP/alu_b_in[28] ), .ZN(
        n3820) );
  XNOR2_X1 U3031 ( .A(\DataP/alu_a_in[29] ), .B(\DataP/alu_b_in[29] ), .ZN(
        n3829) );
  BUF_X1 U3032 ( .A(n3200), .Z(n3201) );
  INV_X1 U3033 ( .A(n3800), .ZN(n3511) );
  NOR2_X1 U3034 ( .A1(n4105), .A2(n2743), .ZN(n2742) );
  XNOR2_X1 U3035 ( .A(\DataP/alu_a_in[22] ), .B(\DataP/alu_b_in[22] ), .ZN(
        n3782) );
  XNOR2_X1 U3036 ( .A(\DataP/alu_a_in[21] ), .B(n2152), .ZN(n3771) );
  XNOR2_X1 U3037 ( .A(\DataP/alu_a_in[24] ), .B(\DataP/alu_b_in[24] ), .ZN(
        n4109) );
  XNOR2_X1 U3038 ( .A(\DataP/alu_a_in[23] ), .B(\DataP/alu_b_in[23] ), .ZN(
        n4108) );
  XNOR2_X1 U3039 ( .A(\DataP/alu_a_in[19] ), .B(n1722), .ZN(n4106) );
  XNOR2_X1 U3040 ( .A(\DataP/alu_a_in[20] ), .B(\DataP/alu_b_in[20] ), .ZN(
        n4107) );
  AND4_X1 U3041 ( .A1(n3747), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n2434)
         );
  XNOR2_X1 U3042 ( .A(\DataP/alu_a_in[9] ), .B(n2166), .ZN(n3494) );
  XNOR2_X1 U3043 ( .A(\DataP/alu_a_in[10] ), .B(n2165), .ZN(n3495) );
  XNOR2_X1 U3044 ( .A(\DataP/alu_a_in[12] ), .B(\lt_x_135/B[12] ), .ZN(n3496)
         );
  XNOR2_X1 U3045 ( .A(\DataP/alu_a_in[18] ), .B(n1736), .ZN(n3747) );
  XNOR2_X1 U3046 ( .A(\DataP/alu_b_in[3] ), .B(n1973), .ZN(n3848) );
  INV_X1 U3047 ( .A(n3540), .ZN(n3541) );
  XNOR2_X1 U3048 ( .A(\DataP/alu_a_in[11] ), .B(n3468), .ZN(n3540) );
  INV_X1 U3049 ( .A(n2151), .ZN(n3468) );
  AOI211_X1 U3050 ( .C1(n3539), .C2(n3554), .A(n3538), .B(n3621), .ZN(n3542)
         );
  XNOR2_X1 U3051 ( .A(\DataP/alu_a_in[15] ), .B(n2230), .ZN(n3621) );
  XNOR2_X1 U3052 ( .A(n3841), .B(\DataP/alu_a_in[8] ), .ZN(n3538) );
  INV_X1 U3053 ( .A(n1575), .ZN(n3841) );
  INV_X1 U3054 ( .A(n2231), .ZN(n3537) );
  INV_X1 U3055 ( .A(n3577), .ZN(n3539) );
  INV_X1 U3056 ( .A(n3591), .ZN(n3536) );
  XNOR2_X1 U3057 ( .A(\DataP/alu_a_in[2] ), .B(n3052), .ZN(n3591) );
  XNOR2_X1 U3058 ( .A(\DataP/alu_a_in[4] ), .B(n3055), .ZN(n3853) );
  XNOR2_X1 U3059 ( .A(\DataP/alu_a_in[6] ), .B(\DataP/alu_b_in[6] ), .ZN(n3859) );
  XNOR2_X1 U3060 ( .A(\DataP/alu_a_in[7] ), .B(\DataP/alu_b_in[7] ), .ZN(n3613) );
  XNOR2_X1 U3061 ( .A(\DataP/alu_a_in[13] ), .B(n2141), .ZN(n3872) );
  XNOR2_X1 U3062 ( .A(\DataP/alu_a_in[16] ), .B(\DataP/alu_b_in[16] ), .ZN(
        n3731) );
  XNOR2_X1 U3063 ( .A(n1751), .B(\DataP/alu_b_in[17] ), .ZN(n3741) );
  XNOR2_X1 U3064 ( .A(\DataP/alu_a_in[14] ), .B(n2145), .ZN(n3875) );
  INV_X1 U3065 ( .A(n3885), .ZN(n3898) );
  XNOR2_X1 U3066 ( .A(\DataP/alu_a_in[31] ), .B(n2121), .ZN(n3885) );
  XNOR2_X1 U3067 ( .A(\DataP/alu_a_in[30] ), .B(\DataP/alu_b_in[30] ), .ZN(
        n3707) );
  NOR2_X1 U3068 ( .A1(n3216), .A2(n2447), .ZN(n3381) );
  NOR2_X1 U3069 ( .A1(n3216), .A2(n2455), .ZN(n3384) );
  OAI21_X1 U3070 ( .B1(n3214), .B2(n109), .A(n3383), .ZN(n3385) );
  AOI22_X1 U3071 ( .A1(n3211), .A2(\DataP/alu_out_M[18] ), .B1(n3208), .B2(
        \DataP/alu_out_W[18] ), .ZN(n3383) );
  NAND4_X1 U3072 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(
        \DataP/alu_b_in[21] ) );
  NAND2_X1 U3073 ( .A1(n3224), .A2(\DataP/alu_out_W[21] ), .ZN(n3550) );
  OR2_X1 U3074 ( .A1(n2771), .A2(n2419), .ZN(n3551) );
  NAND2_X1 U3075 ( .A1(n3223), .A2(\DataP/IMM_s[21] ), .ZN(n3552) );
  NAND2_X1 U3076 ( .A1(n1572), .A2(\DataP/B_s[21] ), .ZN(n3553) );
  NOR2_X1 U3077 ( .A1(n3216), .A2(n2446), .ZN(n3376) );
  OAI21_X1 U3078 ( .B1(n3215), .B2(n121), .A(n3375), .ZN(n3377) );
  AOI22_X1 U3079 ( .A1(n3211), .A2(\DataP/alu_out_M[21] ), .B1(n3207), .B2(
        \DataP/alu_out_W[21] ), .ZN(n3375) );
  NOR2_X1 U3080 ( .A1(n3217), .A2(n2439), .ZN(n3370) );
  OAI21_X1 U3081 ( .B1(n3215), .B2(n129), .A(n3369), .ZN(n3371) );
  AOI22_X1 U3082 ( .A1(n3211), .A2(\DataP/alu_out_M[23] ), .B1(n3207), .B2(
        \DataP/alu_out_W[23] ), .ZN(n3369) );
  NAND4_X1 U3083 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(
        \DataP/alu_b_in[23] ) );
  NAND2_X1 U3084 ( .A1(n3224), .A2(\DataP/alu_out_W[23] ), .ZN(n3543) );
  OR2_X1 U3085 ( .A1(n1627), .A2(n2413), .ZN(n3544) );
  NAND2_X1 U3086 ( .A1(n1614), .A2(\DataP/IMM_s[23] ), .ZN(n3545) );
  NAND2_X1 U3087 ( .A1(n1620), .A2(\DataP/B_s[23] ), .ZN(n3546) );
  NOR2_X1 U3088 ( .A1(n3217), .A2(n2464), .ZN(n3373) );
  OAI21_X1 U3089 ( .B1(n3213), .B2(n125), .A(n3372), .ZN(n3374) );
  AOI22_X1 U3090 ( .A1(n3211), .A2(\DataP/alu_out_M[22] ), .B1(n3207), .B2(
        \DataP/alu_out_W[22] ), .ZN(n3372) );
  NOR2_X1 U3091 ( .A1(n3216), .A2(n2454), .ZN(n3379) );
  OAI21_X1 U3092 ( .B1(n3215), .B2(n117), .A(n3378), .ZN(n3380) );
  AOI22_X1 U3093 ( .A1(n3211), .A2(\DataP/alu_out_M[20] ), .B1(n3207), .B2(
        \DataP/alu_out_W[20] ), .ZN(n3378) );
  NAND2_X1 U3094 ( .A1(n3225), .A2(\DataP/alu_out_W[20] ), .ZN(n3497) );
  OR2_X1 U3095 ( .A1(n2772), .A2(n2420), .ZN(n3498) );
  NAND2_X1 U3096 ( .A1(n2247), .A2(\DataP/IMM_s[20] ), .ZN(n3499) );
  NAND2_X1 U3097 ( .A1(n3221), .A2(\DataP/B_s[20] ), .ZN(n3500) );
  NAND2_X1 U3098 ( .A1(n3224), .A2(\DataP/alu_out_W[16] ), .ZN(n3532) );
  OR2_X1 U3099 ( .A1(n2773), .A2(n2412), .ZN(n3533) );
  NAND2_X1 U3100 ( .A1(n3223), .A2(\DataP/IMM_s[16] ), .ZN(n3534) );
  NAND2_X1 U3101 ( .A1(n3219), .A2(\DataP/B_s[16] ), .ZN(n3535) );
  NOR2_X1 U3102 ( .A1(n3216), .A2(n2465), .ZN(n3387) );
  OAI21_X1 U3103 ( .B1(n3215), .B2(n101), .A(n3386), .ZN(n3388) );
  AOI22_X1 U3104 ( .A1(n2209), .A2(\DataP/alu_out_M[16] ), .B1(n3207), .B2(
        \DataP/alu_out_W[16] ), .ZN(n3386) );
  NAND2_X1 U3105 ( .A1(n3224), .A2(\DataP/alu_out_W[17] ), .ZN(n3519) );
  OR2_X1 U3106 ( .A1(n1627), .A2(n2416), .ZN(n3520) );
  NAND2_X1 U3107 ( .A1(n1623), .A2(\DataP/IMM_s[17] ), .ZN(n3521) );
  NAND2_X1 U3108 ( .A1(n1645), .A2(\DataP/B_s[17] ), .ZN(n3522) );
  AOI22_X1 U3109 ( .A1(n3221), .A2(\DataP/B_s[0] ), .B1(n3222), .B2(
        \DataP/IMM_s[0] ), .ZN(n2656) );
  NOR2_X1 U3110 ( .A1(n3218), .A2(n2461), .ZN(n3333) );
  NOR2_X1 U3111 ( .A1(n3218), .A2(n2460), .ZN(n3331) );
  NAND2_X1 U3112 ( .A1(n3226), .A2(\DataP/alu_out_W[2] ), .ZN(n3311) );
  NOR2_X1 U3113 ( .A1(n3218), .A2(n2459), .ZN(n3329) );
  OAI21_X1 U3114 ( .B1(n3215), .B2(n45), .A(n3328), .ZN(n3330) );
  AOI22_X1 U3115 ( .A1(n3210), .A2(DRAM_ADDRESS[2]), .B1(n3208), .B2(
        \DataP/alu_out_W[2] ), .ZN(n3328) );
  NAND2_X1 U3116 ( .A1(n2246), .A2(\DataP/IMM_s[3] ), .ZN(n2661) );
  NAND2_X1 U3117 ( .A1(n3220), .A2(\DataP/B_s[3] ), .ZN(n2662) );
  NOR2_X1 U3118 ( .A1(n3218), .A2(n2458), .ZN(n3327) );
  NOR2_X1 U3119 ( .A1(n3218), .A2(n2451), .ZN(n3298) );
  OAI21_X1 U3120 ( .B1(n3213), .B2(n65), .A(n3297), .ZN(n3299) );
  AOI22_X1 U3121 ( .A1(n3210), .A2(DRAM_ADDRESS[7]), .B1(n3208), .B2(
        \DataP/alu_out_W[7] ), .ZN(n3297) );
  NAND2_X1 U3122 ( .A1(n3226), .A2(\DataP/alu_out_W[7] ), .ZN(n3300) );
  NAND2_X1 U3123 ( .A1(n3223), .A2(\DataP/IMM_s[7] ), .ZN(n3302) );
  NAND2_X1 U3124 ( .A1(n3225), .A2(\DataP/alu_out_W[6] ), .ZN(n3323) );
  OR2_X1 U3125 ( .A1(n2773), .A2(n2410), .ZN(n3324) );
  NOR2_X1 U3126 ( .A1(n3218), .A2(n2462), .ZN(n3342) );
  OAI21_X1 U3127 ( .B1(n3213), .B2(n61), .A(n3341), .ZN(n3343) );
  AOI22_X1 U3128 ( .A1(n3210), .A2(DRAM_ADDRESS[6]), .B1(n3207), .B2(
        \DataP/alu_out_W[6] ), .ZN(n3341) );
  NAND2_X1 U3129 ( .A1(n3226), .A2(\DataP/alu_out_W[4] ), .ZN(n3315) );
  NOR2_X1 U3130 ( .A1(n3217), .A2(n2443), .ZN(n3339) );
  OAI21_X1 U3131 ( .B1(n3215), .B2(n57), .A(n3338), .ZN(n3340) );
  AOI22_X1 U3132 ( .A1(n3210), .A2(DRAM_ADDRESS[5]), .B1(n3208), .B2(
        \DataP/alu_out_W[5] ), .ZN(n3338) );
  NOR2_X1 U3133 ( .A1(n3214), .A2(n53), .ZN(n3336) );
  OAI21_X1 U3134 ( .B1(n3218), .B2(n2470), .A(n3335), .ZN(n3337) );
  AOI22_X1 U3135 ( .A1(n3210), .A2(DRAM_ADDRESS[4]), .B1(n3208), .B2(
        \DataP/alu_out_W[4] ), .ZN(n3335) );
  OR2_X1 U3136 ( .A1(n2072), .A2(n2518), .ZN(n2692) );
  NOR2_X1 U3137 ( .A1(n3216), .A2(n2449), .ZN(n3399) );
  NAND2_X1 U3138 ( .A1(n3225), .A2(\DataP/alu_out_W[11] ), .ZN(n3454) );
  OR2_X1 U3139 ( .A1(n2773), .A2(n2431), .ZN(n3455) );
  NOR2_X1 U3140 ( .A1(n3217), .A2(n2457), .ZN(n3403) );
  OAI21_X1 U3141 ( .B1(n3215), .B2(n77), .A(n3400), .ZN(n3404) );
  AOI22_X1 U3142 ( .A1(n2209), .A2(DRAM_ADDRESS[10]), .B1(n3209), .B2(
        \DataP/alu_out_W[10] ), .ZN(n3400) );
  NAND2_X1 U3143 ( .A1(n3225), .A2(\DataP/alu_out_W[10] ), .ZN(n3439) );
  OR2_X1 U3144 ( .A1(n2773), .A2(n2409), .ZN(n3440) );
  NOR2_X1 U3145 ( .A1(n3213), .A2(n69), .ZN(n3345) );
  OAI21_X1 U3146 ( .B1(n3218), .B2(n2467), .A(n3344), .ZN(n3346) );
  AOI22_X1 U3147 ( .A1(n3210), .A2(DRAM_ADDRESS[8]), .B1(n3208), .B2(
        \DataP/alu_out_W[8] ), .ZN(n3344) );
  NAND2_X1 U3148 ( .A1(n3225), .A2(\DataP/alu_out_W[8] ), .ZN(n3347) );
  OR2_X1 U3149 ( .A1(n2773), .A2(n2408), .ZN(n3348) );
  NAND4_X1 U3150 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(
        \DataP/alu_b_in[13] ) );
  NAND2_X1 U3151 ( .A1(n3224), .A2(\DataP/alu_out_W[13] ), .ZN(n3524) );
  OR2_X1 U3152 ( .A1(n2772), .A2(n2423), .ZN(n3525) );
  NAND2_X1 U3153 ( .A1(n2247), .A2(\DataP/IMM_s[13] ), .ZN(n3526) );
  NAND2_X1 U3154 ( .A1(n3219), .A2(\DataP/B_s[13] ), .ZN(n3527) );
  NOR2_X1 U3155 ( .A1(n3216), .A2(n2456), .ZN(n3394) );
  OAI21_X1 U3156 ( .B1(n3214), .B2(n89), .A(n3393), .ZN(n3395) );
  AOI22_X1 U3157 ( .A1(n2209), .A2(\DataP/alu_out_M[13] ), .B1(n3208), .B2(
        \DataP/alu_out_W[13] ), .ZN(n3393) );
  NOR2_X1 U3158 ( .A1(n3216), .A2(n2441), .ZN(n3389) );
  NAND2_X1 U3159 ( .A1(n3224), .A2(\DataP/alu_out_W[15] ), .ZN(n3512) );
  OR2_X1 U3160 ( .A1(n2771), .A2(n2433), .ZN(n3513) );
  NAND2_X1 U3161 ( .A1(n2246), .A2(\DataP/IMM_s[15] ), .ZN(n3514) );
  NAND2_X1 U3162 ( .A1(n3219), .A2(\DataP/B_s[15] ), .ZN(n3515) );
  NAND2_X1 U3163 ( .A1(n3224), .A2(\DataP/alu_out_W[14] ), .ZN(n3528) );
  OR2_X1 U3164 ( .A1(n2773), .A2(n2418), .ZN(n3529) );
  NAND2_X1 U3165 ( .A1(n2246), .A2(\DataP/IMM_s[14] ), .ZN(n3530) );
  NAND2_X1 U3166 ( .A1(n3219), .A2(\DataP/B_s[14] ), .ZN(n3531) );
  NOR2_X1 U3167 ( .A1(n3216), .A2(n2448), .ZN(n3391) );
  OAI21_X1 U3168 ( .B1(n3214), .B2(n93), .A(n3390), .ZN(n3392) );
  AOI22_X1 U3169 ( .A1(n2209), .A2(\DataP/alu_out_M[14] ), .B1(n3209), .B2(
        \DataP/alu_out_W[14] ), .ZN(n3390) );
  NOR2_X1 U3170 ( .A1(n3216), .A2(n2442), .ZN(n3397) );
  AOI22_X1 U3171 ( .A1(n2209), .A2(\DataP/alu_out_M[12] ), .B1(n3208), .B2(
        \DataP/alu_out_W[12] ), .ZN(n3396) );
  BUF_X1 U3172 ( .A(n1762), .Z(\lt_x_135/B[12] ) );
  NAND2_X1 U3173 ( .A1(n3219), .A2(\DataP/B_s[12] ), .ZN(n3478) );
  OR2_X1 U3174 ( .A1(n2773), .A2(n2424), .ZN(n3476) );
  NAND2_X1 U3175 ( .A1(n3225), .A2(\DataP/alu_out_W[12] ), .ZN(n3475) );
  NAND2_X1 U3176 ( .A1(n3226), .A2(\DataP/alu_out_W[9] ), .ZN(n3260) );
  NAND2_X1 U3177 ( .A1(n2247), .A2(\DataP/IMM_s[9] ), .ZN(n3262) );
  NAND4_X1 U3178 ( .A1(n3523), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(
        \DataP/alu_b_in[27] ) );
  NAND2_X1 U3179 ( .A1(n3224), .A2(\DataP/alu_out_W[27] ), .ZN(n3507) );
  OR2_X1 U3180 ( .A1(n1627), .A2(n2411), .ZN(n3508) );
  NAND2_X1 U3181 ( .A1(n2227), .A2(\DataP/B_s[27] ), .ZN(n3509) );
  NOR2_X1 U3182 ( .A1(n3217), .A2(n2445), .ZN(n3361) );
  OAI21_X1 U3183 ( .B1(n3214), .B2(n141), .A(n3360), .ZN(n3362) );
  AOI22_X1 U3184 ( .A1(n3211), .A2(\DataP/alu_out_M[26] ), .B1(n3208), .B2(
        \DataP/alu_out_W[26] ), .ZN(n3360) );
  NAND4_X1 U3185 ( .A1(n3523), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(
        \DataP/alu_b_in[26] ) );
  NAND2_X1 U3186 ( .A1(n3225), .A2(\DataP/alu_out_W[26] ), .ZN(n3501) );
  OR2_X1 U3187 ( .A1(n1627), .A2(n2415), .ZN(n3502) );
  NAND2_X1 U3188 ( .A1(n2227), .A2(\DataP/B_s[26] ), .ZN(n3503) );
  NOR2_X1 U3189 ( .A1(n3217), .A2(n2453), .ZN(n3364) );
  OAI21_X1 U3190 ( .B1(n3214), .B2(n137), .A(n3363), .ZN(n3365) );
  AOI22_X1 U3191 ( .A1(n3211), .A2(\DataP/alu_out_M[25] ), .B1(n3208), .B2(
        \DataP/alu_out_W[25] ), .ZN(n3363) );
  OR2_X1 U3192 ( .A1(n2772), .A2(n2422), .ZN(n3504) );
  NAND2_X1 U3193 ( .A1(n3225), .A2(\DataP/alu_out_W[25] ), .ZN(n3505) );
  NAND2_X1 U3194 ( .A1(n1645), .A2(\DataP/B_s[25] ), .ZN(n3506) );
  NOR2_X1 U3195 ( .A1(n3217), .A2(n2463), .ZN(n3367) );
  OAI21_X1 U3196 ( .B1(n3213), .B2(n133), .A(n3366), .ZN(n3368) );
  AOI22_X1 U3197 ( .A1(n3211), .A2(\DataP/alu_out_M[24] ), .B1(n3208), .B2(
        \DataP/alu_out_W[24] ), .ZN(n3366) );
  NAND4_X1 U3198 ( .A1(n3523), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(
        \DataP/alu_b_in[31] ) );
  NAND2_X1 U3199 ( .A1(n3224), .A2(\DataP/alu_out_W[31] ), .ZN(n3516) );
  OR2_X1 U3200 ( .A1(n1627), .A2(n2414), .ZN(n3517) );
  NAND2_X1 U3201 ( .A1(n2227), .A2(\DataP/B_s[31] ), .ZN(n3518) );
  NOR2_X1 U3202 ( .A1(n2539), .A2(n2405), .ZN(n2538) );
  NOR2_X1 U3203 ( .A1(n3217), .A2(n2437), .ZN(n3352) );
  OAI21_X1 U3204 ( .B1(n3215), .B2(n157), .A(n3351), .ZN(n3353) );
  AOI22_X1 U3205 ( .A1(n3210), .A2(\DataP/alu_out_M[30] ), .B1(n3208), .B2(
        \DataP/alu_out_W[30] ), .ZN(n3351) );
  NOR2_X1 U3206 ( .A1(n3217), .A2(n2444), .ZN(n3355) );
  OAI21_X1 U3207 ( .B1(n3213), .B2(n153), .A(n3354), .ZN(n3356) );
  AOI22_X1 U3208 ( .A1(n3211), .A2(\DataP/alu_out_M[29] ), .B1(n3207), .B2(
        \DataP/alu_out_W[29] ), .ZN(n3354) );
  NAND2_X1 U3209 ( .A1(n2246), .A2(\DataP/IMM_s[30] ), .ZN(n3523) );
  NOR2_X1 U3210 ( .A1(n3253), .A2(n3252), .ZN(n3257) );
  XNOR2_X1 U3211 ( .A(\DataP/Rs2[0] ), .B(n528), .ZN(n3253) );
  NOR2_X1 U3212 ( .A1(n3255), .A2(n3254), .ZN(n3256) );
  XNOR2_X1 U3213 ( .A(\DataP/Rs2[2] ), .B(n530), .ZN(n3254) );
  XNOR2_X1 U3214 ( .A(\DataP/Rs2[3] ), .B(n2777), .ZN(n3255) );
  NOR2_X1 U3215 ( .A1(n3217), .A2(n2452), .ZN(n3358) );
  OAI21_X1 U3216 ( .B1(n3214), .B2(n149), .A(n3357), .ZN(n3359) );
  AOI22_X1 U3217 ( .A1(n3211), .A2(\DataP/alu_out_M[28] ), .B1(n3207), .B2(
        \DataP/alu_out_W[28] ), .ZN(n3357) );
  NOR2_X1 U3218 ( .A1(n3246), .A2(n3883), .ZN(n2629) );
  INV_X1 U3219 ( .A(Rst), .ZN(n2628) );
  AOI21_X1 U3220 ( .B1(n3287), .B2(n17), .A(n3286), .ZN(n3296) );
  NOR2_X1 U3221 ( .A1(n3285), .A2(n3284), .ZN(n3286) );
  NOR2_X1 U3222 ( .A1(n3280), .A2(n521), .ZN(n3281) );
  NOR2_X1 U3223 ( .A1(n3279), .A2(n3288), .ZN(n3910) );
  NOR2_X1 U3224 ( .A1(n3278), .A2(n3277), .ZN(n3290) );
  NAND4_X1 U3225 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3278)
         );
  XNOR2_X1 U3226 ( .A(n530), .B(\DataP/Rs1[2] ), .ZN(n3270) );
  XNOR2_X1 U3227 ( .A(n528), .B(n2392), .ZN(n3268) );
  AOI21_X1 U3228 ( .B1(n3265), .B2(n3264), .A(n2091), .ZN(n3288) );
  NAND3_X1 U3229 ( .A1(n3239), .A2(\DataP/opcode_W[3] ), .A3(n2625), .ZN(n2635) );
  NAND2_X1 U3230 ( .A1(n2622), .A2(n2624), .ZN(n3265) );
  AND2_X1 U3231 ( .A1(n3902), .A2(n3884), .ZN(n2376) );
  AND2_X1 U3232 ( .A1(n1570), .A2(n2238), .ZN(n2378) );
  OR2_X1 U3233 ( .A1(\DataP/alu_b_in[29] ), .A2(\DataP/alu_b_in[28] ), .ZN(
        n2381) );
  OAI211_X1 U3234 ( .C1(n3621), .C2(n2108), .A(n3638), .B(n2577), .ZN(n2758)
         );
  OR2_X1 U3235 ( .A1(n3217), .A2(n2436), .ZN(n2384) );
  INV_X1 U3236 ( .A(n2740), .ZN(n2738) );
  AND2_X1 U3237 ( .A1(\DataP/alu_a_in[21] ), .A2(n2679), .ZN(n2388) );
  INV_X1 U3238 ( .A(n1618), .ZN(n2754) );
  NOR2_X1 U3239 ( .A1(n3430), .A2(n4101), .ZN(n3904) );
  INV_X1 U3240 ( .A(n2165), .ZN(n3459) );
  INV_X1 U3241 ( .A(n2233), .ZN(n3046) );
  AND2_X1 U3242 ( .A1(\DataP/alu_a_in[13] ), .A2(n2737), .ZN(n2393) );
  AND2_X1 U3243 ( .A1(n2763), .A2(n2238), .ZN(n2394) );
  AND2_X1 U3244 ( .A1(n1723), .A2(n3762), .ZN(n2396) );
  INV_X1 U3245 ( .A(n3851), .ZN(n3890) );
  AND2_X1 U3246 ( .A1(\DataP/alu_a_in[17] ), .A2(n2721), .ZN(n2397) );
  XOR2_X1 U3247 ( .A(n3816), .B(n3817), .Z(n2400) );
  INV_X1 U3248 ( .A(n3797), .ZN(n2744) );
  INV_X1 U3249 ( .A(n3296), .ZN(n2619) );
  NAND2_X1 U3250 ( .A1(n3689), .A2(\DataP/alu_a_in[23] ), .ZN(n3715) );
  OR2_X1 U3251 ( .A1(n2727), .A2(n3788), .ZN(n2404) );
  NAND2_X1 U3252 ( .A1(n3727), .A2(\DataP/alu_a_in[29] ), .ZN(n3825) );
  INV_X1 U3253 ( .A(n3825), .ZN(n2746) );
  AND2_X1 U3254 ( .A1(n3210), .A2(\DataP/alu_out_M[31] ), .ZN(n2405) );
  INV_X1 U3255 ( .A(n3826), .ZN(n2750) );
  AND3_X1 U3256 ( .A1(n3835), .A2(n3482), .A3(n3483), .ZN(n2473) );
  NOR2_X1 U3257 ( .A1(n4110), .A2(n4192), .ZN(n2474) );
  AND2_X1 U3258 ( .A1(n2725), .A2(n2394), .ZN(n2476) );
  AND2_X1 U3259 ( .A1(n3624), .A2(n2108), .ZN(n2479) );
  OR2_X1 U3260 ( .A1(n2756), .A2(n2129), .ZN(n2482) );
  NAND2_X1 U3261 ( .A1(n2525), .A2(n2524), .ZN(n3682) );
  NAND2_X1 U3262 ( .A1(n3665), .A2(n2114), .ZN(n3766) );
  INV_X1 U3263 ( .A(n3766), .ZN(n2607) );
  INV_X1 U3264 ( .A(\DataP/alu_b_in[30] ), .ZN(n2614) );
  OR2_X1 U3265 ( .A1(n1600), .A2(n2535), .ZN(n2486) );
  AND2_X1 U3266 ( .A1(\DataP/alu_a_in[22] ), .A2(n2569), .ZN(n2487) );
  AND2_X1 U3267 ( .A1(n2755), .A2(n2749), .ZN(n2488) );
  NAND2_X1 U3268 ( .A1(n3720), .A2(\DataP/alu_a_in[27] ), .ZN(n3721) );
  OR2_X1 U3269 ( .A1(n3825), .A2(n3826), .ZN(n2489) );
  AND2_X1 U3270 ( .A1(n2111), .A2(n2676), .ZN(n2490) );
  INV_X1 U3271 ( .A(Rst), .ZN(n3234) );
  NAND2_X1 U3272 ( .A1(n3648), .A2(\DataP/alu_a_in[19] ), .ZN(n3685) );
  NAND2_X1 U3273 ( .A1(n2615), .A2(n2733), .ZN(n3648) );
  AND2_X1 U3274 ( .A1(n1750), .A2(n2529), .ZN(n2528) );
  NAND2_X1 U3275 ( .A1(n2721), .A2(n2128), .ZN(n2529) );
  INV_X1 U3276 ( .A(n3666), .ZN(n3665) );
  OR2_X1 U3277 ( .A1(n2630), .A2(n2598), .ZN(n2530) );
  INV_X1 U3278 ( .A(n2653), .ZN(n2532) );
  NAND4_X1 U3279 ( .A1(n1734), .A2(n2219), .A3(n2220), .A4(n3684), .ZN(n2533)
         );
  AOI21_X1 U3280 ( .B1(n2536), .B2(n2129), .A(n3775), .ZN(n313) );
  XNOR2_X1 U3281 ( .A(n2537), .B(n2396), .ZN(n2536) );
  AOI21_X1 U3282 ( .B1(n3767), .B2(n3766), .A(n3765), .ZN(n2537) );
  OAI22_X1 U3283 ( .A1(n3213), .A2(n161), .B1(n2072), .B2(n2517), .ZN(n2539)
         );
  NAND2_X1 U3284 ( .A1(\DataP/alu_b_in[27] ), .A2(n2535), .ZN(n2540) );
  XNOR2_X1 U3285 ( .A(n2541), .B(n3635), .ZN(n2689) );
  OAI21_X1 U3286 ( .B1(n3874), .B2(n3636), .A(n3631), .ZN(n2541) );
  AOI21_X1 U3287 ( .B1(n2542), .B2(n3630), .A(n3867), .ZN(n3874) );
  OAI21_X1 U3288 ( .B1(n3864), .B2(n3617), .A(n3863), .ZN(n2542) );
  AOI21_X1 U3289 ( .B1(n2543), .B2(n2129), .A(n3746), .ZN(n323) );
  XNOR2_X1 U3290 ( .A(n2544), .B(n2155), .ZN(n2543) );
  AOI21_X1 U3291 ( .B1(n3729), .B2(n2238), .A(n2545), .ZN(n2544) );
  INV_X1 U3292 ( .A(n1663), .ZN(n2545) );
  OAI211_X1 U3293 ( .C1(n4111), .C2(n2558), .A(n2550), .B(n2553), .ZN(
        \DataP/PC_reg/N33 ) );
  INV_X1 U3294 ( .A(n2551), .ZN(n2550) );
  OR2_X1 U3295 ( .A1(n4110), .A2(n4191), .ZN(n2552) );
  NAND2_X1 U3296 ( .A1(n2554), .A2(n2131), .ZN(n2553) );
  INV_X1 U3297 ( .A(n2556), .ZN(n2554) );
  AND2_X1 U3298 ( .A1(n2557), .A2(n2753), .ZN(n2556) );
  NAND2_X1 U3299 ( .A1(n2083), .A2(n2751), .ZN(n2558) );
  NAND2_X1 U3300 ( .A1(n2783), .A2(n1646), .ZN(n3690) );
  NAND2_X1 U3301 ( .A1(n2559), .A2(n2759), .ZN(n3767) );
  NAND2_X1 U3302 ( .A1(n2476), .A2(n2700), .ZN(n2559) );
  AND2_X1 U3303 ( .A1(n2724), .A2(n3635), .ZN(n2700) );
  OAI22_X1 U3304 ( .A1(n303), .A2(n4111), .B1(n4110), .B2(n4196), .ZN(
        \DataP/PC_reg/N28 ) );
  AOI21_X1 U3305 ( .B1(n2561), .B2(n2129), .A(n3815), .ZN(n303) );
  XNOR2_X1 U3306 ( .A(n1711), .B(n3807), .ZN(n2561) );
  AOI21_X1 U3307 ( .B1(n3824), .B2(n2131), .A(n2563), .ZN(n2562) );
  NOR2_X1 U3308 ( .A1(n4110), .A2(n4194), .ZN(n2563) );
  NOR2_X1 U3309 ( .A1(n3880), .A2(n4111), .ZN(n2564) );
  NAND2_X1 U3310 ( .A1(n3762), .A2(n3764), .ZN(n3667) );
  NAND2_X1 U3311 ( .A1(n3666), .A2(\DataP/alu_a_in[20] ), .ZN(n3764) );
  OAI21_X1 U3312 ( .B1(n3886), .B2(n2678), .A(n2388), .ZN(n3762) );
  NAND2_X1 U3313 ( .A1(n2568), .A2(n2487), .ZN(n3714) );
  NAND2_X1 U3314 ( .A1(n3670), .A2(n2402), .ZN(n2568) );
  XNOR2_X1 U3315 ( .A(n2570), .B(n2122), .ZN(n3670) );
  NOR2_X1 U3316 ( .A1(n3668), .A2(n3669), .ZN(n2570) );
  NAND2_X1 U3317 ( .A1(n2576), .A2(n2571), .ZN(n2709) );
  NAND3_X1 U3318 ( .A1(n2595), .A2(n2376), .A3(n2070), .ZN(n2571) );
  NAND2_X1 U3319 ( .A1(n2595), .A2(n2572), .ZN(n2574) );
  NOR2_X1 U3320 ( .A1(n2719), .A2(n2573), .ZN(n2572) );
  NAND2_X1 U3321 ( .A1(n2376), .A2(n2575), .ZN(n2573) );
  OAI21_X1 U3322 ( .B1(n3215), .B2(n49), .A(n2579), .ZN(n2578) );
  AOI22_X1 U3323 ( .A1(n3210), .A2(DRAM_ADDRESS[3]), .B1(n3209), .B2(
        \DataP/alu_out_W[3] ), .ZN(n2579) );
  INV_X1 U3324 ( .A(n1635), .ZN(n2580) );
  NAND2_X1 U3325 ( .A1(n1564), .A2(n2747), .ZN(n2581) );
  NAND2_X1 U3326 ( .A1(n2584), .A2(n3721), .ZN(n2582) );
  INV_X1 U3327 ( .A(n2096), .ZN(n2584) );
  NAND2_X1 U3328 ( .A1(n2587), .A2(n2108), .ZN(n2586) );
  XNOR2_X1 U3329 ( .A(n2589), .B(n2588), .ZN(n2587) );
  NAND2_X1 U3330 ( .A1(n1574), .A2(n2107), .ZN(n2589) );
  NAND2_X1 U3331 ( .A1(n2590), .A2(n2591), .ZN(\DataP/PC_reg/N29 ) );
  NAND2_X1 U3332 ( .A1(n2719), .A2(n2710), .ZN(n2593) );
  XNOR2_X1 U3333 ( .A(n1594), .B(\DataP/alu_a_in[23] ), .ZN(n3713) );
  OAI21_X1 U3334 ( .B1(n2596), .B2(n2535), .A(n2701), .ZN(n3689) );
  XNOR2_X1 U3335 ( .A(n2597), .B(n2124), .ZN(n2596) );
  NOR2_X1 U3336 ( .A1(n3669), .A2(n2702), .ZN(n2597) );
  OAI21_X1 U3337 ( .B1(n2610), .B2(n3489), .A(n2600), .ZN(n3860) );
  AOI21_X1 U3338 ( .B1(n3486), .B2(n2601), .A(n2235), .ZN(n2600) );
  NAND2_X1 U3339 ( .A1(n3487), .A2(n2473), .ZN(n2610) );
  NAND2_X1 U3340 ( .A1(n3860), .A2(n3628), .ZN(n3864) );
  INV_X1 U3341 ( .A(n3489), .ZN(n2601) );
  NAND2_X1 U3342 ( .A1(n2602), .A2(n3753), .ZN(n2603) );
  AND2_X1 U3343 ( .A1(n3766), .A2(n1588), .ZN(n3753) );
  OAI211_X1 U3344 ( .C1(n2604), .C2(n2607), .A(n2603), .B(n3686), .ZN(n2605)
         );
  OR2_X1 U3345 ( .A1(n2606), .A2(n3687), .ZN(n2604) );
  NAND2_X1 U3346 ( .A1(n2605), .A2(n2608), .ZN(n3716) );
  INV_X1 U3347 ( .A(n3776), .ZN(n2608) );
  NAND2_X1 U3348 ( .A1(n3688), .A2(n1717), .ZN(n3776) );
  NAND2_X1 U3349 ( .A1(n3671), .A2(n3778), .ZN(n3688) );
  NAND3_X1 U3350 ( .A1(n1745), .A2(n2609), .A3(n3634), .ZN(n2725) );
  NAND3_X1 U3351 ( .A1(n2610), .A2(n3488), .A3(n2222), .ZN(n2609) );
  NAND2_X1 U3352 ( .A1(n2430), .A2(n2613), .ZN(n3887) );
  OAI21_X1 U3353 ( .B1(n2385), .B2(n3722), .A(n3885), .ZN(n2613) );
  AOI21_X1 U3354 ( .B1(n3647), .B2(n2617), .A(n2616), .ZN(n2615) );
  NAND2_X1 U3355 ( .A1(n2730), .A2(n2734), .ZN(n2616) );
  NAND2_X1 U3356 ( .A1(n2618), .A2(n3909), .ZN(n3212) );
  NAND2_X1 U3357 ( .A1(n3295), .A2(n3296), .ZN(n2618) );
  NAND2_X1 U3358 ( .A1(n3293), .A2(n2629), .ZN(n3295) );
  NAND2_X1 U3359 ( .A1(n2085), .A2(n3258), .ZN(n2781) );
  AND2_X1 U3360 ( .A1(n3256), .A2(n3257), .ZN(n2621) );
  NAND3_X1 U3361 ( .A1(n2635), .A2(n2622), .A3(n2624), .ZN(n2639) );
  NAND2_X1 U3362 ( .A1(n2480), .A2(n2623), .ZN(n2622) );
  XNOR2_X1 U3363 ( .A(n2779), .B(n2383), .ZN(n2623) );
  NAND2_X1 U3364 ( .A1(n2483), .A2(\DataP/opcode_W[1] ), .ZN(n2624) );
  OAI211_X1 U3365 ( .C1(\DataP/opcode_W[0] ), .C2(\DataP/opcode_W[4] ), .A(
        \DataP/opcode_W[2] ), .B(\DataP/opcode_W[1] ), .ZN(n2625) );
  OAI21_X1 U3366 ( .B1(n2213), .B2(\DataP/alu_b_in[20] ), .A(n3663), .ZN(n2630) );
  NAND2_X1 U3367 ( .A1(n2152), .A2(n3664), .ZN(n2631) );
  NAND4_X1 U3368 ( .A1(n2634), .A2(n3292), .A3(n2633), .A4(n2632), .ZN(n3402)
         );
  OR2_X1 U3369 ( .A1(n3295), .A2(n1718), .ZN(n2632) );
  AOI21_X1 U3370 ( .B1(n3909), .B2(n2619), .A(n2475), .ZN(n2633) );
  NAND2_X1 U3371 ( .A1(n2635), .A2(\DataP/opcode_W[5] ), .ZN(n2638) );
  NAND4_X1 U3372 ( .A1(n2640), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3289)
         );
  NOR2_X1 U3373 ( .A1(n3241), .A2(n2641), .ZN(n2640) );
  XNOR2_X1 U3374 ( .A(n2775), .B(\DataP/dest_M[3] ), .ZN(n2641) );
  AOI21_X1 U3375 ( .B1(n3481), .B2(n1726), .A(n2644), .ZN(n2643) );
  NAND2_X1 U3376 ( .A1(n2646), .A2(n2645), .ZN(n2644) );
  NAND2_X1 U3377 ( .A1(n2393), .A2(n2738), .ZN(n2645) );
  NAND2_X1 U3378 ( .A1(n2735), .A2(n2736), .ZN(n2646) );
  NAND2_X1 U3379 ( .A1(n1713), .A2(n2393), .ZN(n2647) );
  NAND2_X1 U3380 ( .A1(n2648), .A2(n2649), .ZN(n3632) );
  NAND2_X1 U3381 ( .A1(n2685), .A2(n2651), .ZN(n2648) );
  INV_X1 U3382 ( .A(\DataP/alu_a_in[14] ), .ZN(n2652) );
  NAND2_X1 U3383 ( .A1(n2667), .A2(n2665), .ZN(n2716) );
  NOR2_X1 U3384 ( .A1(n3633), .A2(n2758), .ZN(n2665) );
  NAND2_X1 U3385 ( .A1(n2666), .A2(n3873), .ZN(n3633) );
  NAND2_X1 U3386 ( .A1(n3860), .A2(n1634), .ZN(n2667) );
  NOR2_X1 U3387 ( .A1(n3861), .A2(n3868), .ZN(n3634) );
  NAND2_X1 U3388 ( .A1(n3414), .A2(n2206), .ZN(n3574) );
  NAND3_X1 U3389 ( .A1(n2725), .A2(n2724), .A3(n3635), .ZN(n2783) );
  NAND2_X1 U3390 ( .A1(n2111), .A2(n2108), .ZN(n2677) );
  NAND2_X1 U3391 ( .A1(n3663), .A2(n3886), .ZN(n2679) );
  NAND2_X1 U3392 ( .A1(\DataP/alu_b_in[6] ), .A2(n3886), .ZN(n2680) );
  NAND2_X1 U3393 ( .A1(n3841), .A2(n3886), .ZN(n2686) );
  OAI211_X1 U3394 ( .C1(n3215), .C2(n81), .A(n2692), .B(n2691), .ZN(n2690) );
  NAND2_X1 U3395 ( .A1(n2209), .A2(DRAM_ADDRESS[11]), .ZN(n2691) );
  AOI21_X1 U3396 ( .B1(n2695), .B2(n2698), .A(n2694), .ZN(n2696) );
  INV_X1 U3397 ( .A(n3686), .ZN(n2694) );
  INV_X1 U3398 ( .A(n2759), .ZN(n2695) );
  NAND4_X1 U3399 ( .A1(n2700), .A2(n2223), .A3(n2394), .A4(n2698), .ZN(n2697)
         );
  NOR2_X1 U3400 ( .A1(n2699), .A2(n2607), .ZN(n2698) );
  INV_X1 U3401 ( .A(n1723), .ZN(n2699) );
  NAND3_X1 U3402 ( .A1(n3889), .A2(n2129), .A3(n3902), .ZN(n2704) );
  OAI21_X1 U3403 ( .B1(n2709), .B2(n2708), .A(n2707), .ZN(\DataP/PC_reg/N32 )
         );
  INV_X1 U3404 ( .A(n2376), .ZN(n2710) );
  NAND2_X1 U3405 ( .A1(n1552), .A2(n1619), .ZN(n2729) );
  NAND3_X1 U3406 ( .A1(n2716), .A2(n2718), .A3(n2713), .ZN(n2711) );
  NAND2_X1 U3407 ( .A1(n2484), .A2(n2718), .ZN(n2712) );
  AND2_X1 U3408 ( .A1(n3712), .A2(n2714), .ZN(n2713) );
  AOI21_X1 U3409 ( .B1(n3635), .B2(n3636), .A(n2715), .ZN(n2714) );
  INV_X1 U3410 ( .A(n3715), .ZN(n2715) );
  OR2_X1 U3411 ( .A1(\DataP/alu_b_in[17] ), .A2(n2108), .ZN(n2721) );
  NAND2_X1 U3412 ( .A1(\DataP/alu_b_in[26] ), .A2(n2535), .ZN(n2722) );
  NOR2_X1 U3413 ( .A1(n3693), .A2(n3694), .ZN(n2723) );
  NAND2_X1 U3414 ( .A1(n3716), .A2(n2726), .ZN(n2728) );
  INV_X1 U3415 ( .A(n3718), .ZN(n2727) );
  NAND2_X1 U3416 ( .A1(n1600), .A2(n2535), .ZN(n2734) );
  NAND2_X1 U3417 ( .A1(n1573), .A2(n2128), .ZN(n2739) );
  NAND2_X1 U3418 ( .A1(n2141), .A2(n2128), .ZN(n2740) );
  NAND2_X1 U3419 ( .A1(n1736), .A2(n2535), .ZN(n2757) );
  AND2_X1 U3420 ( .A1(n1636), .A2(n2224), .ZN(n2764) );
  AOI21_X1 U3421 ( .B1(n3283), .B2(\DataP/opcode_E[4] ), .A(n17), .ZN(n3285)
         );
  NAND2_X1 U3422 ( .A1(n3226), .A2(\DataP/alu_out_W[0] ), .ZN(n3308) );
  NAND2_X1 U3423 ( .A1(n3226), .A2(\DataP/alu_out_W[3] ), .ZN(n3310) );
  INV_X1 U3424 ( .A(n2782), .ZN(n2771) );
  NAND2_X1 U3425 ( .A1(n3221), .A2(\DataP/B_s[8] ), .ZN(n3350) );
  NAND2_X1 U3426 ( .A1(n3219), .A2(\DataP/B_s[11] ), .ZN(n3457) );
  NAND2_X1 U3427 ( .A1(n3219), .A2(\DataP/B_s[2] ), .ZN(n3314) );
  NAND2_X1 U3428 ( .A1(n3221), .A2(\DataP/B_s[6] ), .ZN(n3326) );
  NAND2_X1 U3429 ( .A1(n3221), .A2(\DataP/B_s[9] ), .ZN(n3263) );
  NAND2_X1 U3430 ( .A1(n3219), .A2(\DataP/B_s[10] ), .ZN(n3442) );
  NAND2_X1 U3431 ( .A1(n3220), .A2(\DataP/B_s[4] ), .ZN(n3318) );
  NAND2_X1 U3432 ( .A1(n3219), .A2(\DataP/B_s[7] ), .ZN(n3303) );
  NAND2_X1 U3433 ( .A1(n3220), .A2(\DataP/B_s[5] ), .ZN(n3322) );
  OR2_X1 U3434 ( .A1(n2773), .A2(n2450), .ZN(n3320) );
  NAND2_X1 U3435 ( .A1(n3226), .A2(\DataP/alu_out_W[5] ), .ZN(n3319) );
  NAND2_X1 U3436 ( .A1(n3763), .A2(n3667), .ZN(n3686) );
  XNOR2_X1 U3437 ( .A(n2069), .B(n2407), .ZN(n3275) );
  XNOR2_X1 U3438 ( .A(n1638), .B(n538), .ZN(n3243) );
  NOR2_X1 U3439 ( .A1(\DataP/dest_M[4] ), .A2(n1621), .ZN(n3249) );
  XNOR2_X1 U3440 ( .A(n2392), .B(n1630), .ZN(n3276) );
  XNOR2_X1 U3441 ( .A(n528), .B(n536), .ZN(n3242) );
  NAND2_X1 U3442 ( .A1(n3238), .A2(\DataP/opcode_W[5] ), .ZN(n3239) );
  NAND2_X1 U3443 ( .A1(n3226), .A2(\DataP/alu_out_W[1] ), .ZN(n3304) );
  XNOR2_X1 U3444 ( .A(n529), .B(\DataP/Rs1[1] ), .ZN(n3269) );
  XNOR2_X1 U3445 ( .A(\DataP/Rs2[1] ), .B(n529), .ZN(n3252) );
  XNOR2_X1 U3446 ( .A(n1628), .B(n524), .ZN(n3273) );
  XNOR2_X1 U3447 ( .A(\DataP/dest_M[4] ), .B(n540), .ZN(n3241) );
  AND2_X1 U3448 ( .A1(n2220), .A2(n2167), .ZN(n2784) );
  XNOR2_X1 U3449 ( .A(n2199), .B(n2784), .ZN(n3751) );
  XNOR2_X1 U3450 ( .A(\DataP/add_D[1] ), .B(n2429), .ZN(n3277) );
  XNOR2_X1 U3451 ( .A(\DataP/add_D[1] ), .B(\DataP/Rs2[1] ), .ZN(n3240) );
  XNOR2_X1 U3452 ( .A(\DataP/dest_M[1] ), .B(\DataP/add_D[1] ), .ZN(n3244) );
  OAI21_X1 U3453 ( .B1(\DataP/opcode_W[1] ), .B2(\DataP/opcode_W[2] ), .A(
        \DataP/opcode_W[4] ), .ZN(n3238) );
  XNOR2_X1 U3454 ( .A(n3650), .B(n2168), .ZN(n3658) );
  NOR2_X1 U3455 ( .A1(n21), .A2(\DataP/opcode_E[0] ), .ZN(n3282) );
  NAND2_X1 U3456 ( .A1(n3537), .A2(n3199), .ZN(n3554) );
  NAND2_X1 U3457 ( .A1(n521), .A2(n520), .ZN(n3283) );
  XNOR2_X1 U3458 ( .A(\DataP/alu_a_in[5] ), .B(\lt_x_135/B[5] ), .ZN(n3603) );
  INV_X1 U3459 ( .A(n2095), .ZN(n3862) );
  NAND2_X1 U3460 ( .A1(n3220), .A2(\DataP/B_s[1] ), .ZN(n3307) );
  XNOR2_X1 U3461 ( .A(n1757), .B(n523), .ZN(n3274) );
  NAND2_X1 U3462 ( .A1(n2780), .A2(n3258), .ZN(n3549) );
  OAI21_X1 U3463 ( .B1(n521), .B2(n3883), .A(Rst), .ZN(
        \DataP/FORWARDING_BR/N12 ) );
  NAND2_X1 U3464 ( .A1(n2248), .A2(n3272), .ZN(n3294) );
  NOR2_X1 U3465 ( .A1(\DataP/opcode_M[2] ), .A2(\DataP/opcode_M[1] ), .ZN(
        n3247) );
  XNOR2_X1 U3466 ( .A(n2232), .B(n3047), .ZN(n3579) );
  OAI21_X1 U3467 ( .B1(n521), .B2(n520), .A(\DataP/opcode_E[3] ), .ZN(n3284)
         );
  OR2_X1 U3468 ( .A1(n3293), .A2(n3291), .ZN(n3292) );
  NAND2_X1 U3469 ( .A1(n3416), .A2(n1716), .ZN(n3410) );
  XNOR2_X1 U3470 ( .A(n2250), .B(n1567), .ZN(n3413) );
  NAND2_X1 U3471 ( .A1(n2246), .A2(\DataP/IMM_s[11] ), .ZN(n3456) );
  NAND2_X1 U3472 ( .A1(n1581), .A2(\DataP/IMM_s[8] ), .ZN(n3349) );
  NAND2_X1 U3473 ( .A1(n3223), .A2(\DataP/IMM_s[10] ), .ZN(n3441) );
  NAND2_X1 U3474 ( .A1(n3223), .A2(\DataP/IMM_s[6] ), .ZN(n3325) );
  NAND2_X1 U3475 ( .A1(n2247), .A2(\DataP/IMM_s[12] ), .ZN(n3477) );
  OR2_X1 U3476 ( .A1(n2773), .A2(n2477), .ZN(n3261) );
  NAND2_X1 U3477 ( .A1(n3222), .A2(\DataP/IMM_s[4] ), .ZN(n3317) );
  OR2_X1 U3478 ( .A1(n2773), .A2(n2468), .ZN(n3301) );
  OR2_X1 U3479 ( .A1(n2771), .A2(n2466), .ZN(n3316) );
  NAND2_X1 U3480 ( .A1(n1581), .A2(\DataP/IMM_s[2] ), .ZN(n3313) );
  NAND2_X1 U3481 ( .A1(n2247), .A2(\DataP/IMM_s[5] ), .ZN(n3321) );
  OR2_X1 U3482 ( .A1(n2773), .A2(n2472), .ZN(n3309) );
  NAND2_X1 U3483 ( .A1(n3223), .A2(\DataP/IMM_s[1] ), .ZN(n3306) );
  OR2_X1 U3484 ( .A1(n2773), .A2(n2469), .ZN(n3305) );
  NAND4_X1 U3485 ( .A1(n2201), .A2(n2918), .A3(n2126), .A4(n2916), .ZN(n2853)
         );
  NOR2_X1 U3486 ( .A1(n3204), .A2(n2853), .ZN(n2810) );
  NAND2_X1 U3487 ( .A1(n2231), .A2(n2916), .ZN(n2785) );
  AOI22_X1 U3488 ( .A1(n2103), .A2(n2232), .B1(\DataP/alu_a_in[2] ), .B2(n2916), .ZN(n2787) );
  AOI22_X1 U3489 ( .A1(n2917), .A2(n2785), .B1(n2787), .B2(n2105), .ZN(n2799)
         );
  NAND2_X1 U3490 ( .A1(n2918), .A2(n2799), .ZN(n2820) );
  AOI22_X1 U3491 ( .A1(n2103), .A2(n1973), .B1(\DataP/alu_a_in[4] ), .B2(n2916), .ZN(n2786) );
  AOI22_X1 U3492 ( .A1(n2103), .A2(\DataP/alu_a_in[5] ), .B1(
        \DataP/alu_a_in[6] ), .B2(n2916), .ZN(n2790) );
  AOI22_X1 U3493 ( .A1(n2917), .A2(n2786), .B1(n2790), .B2(n2105), .ZN(n2798)
         );
  AOI22_X1 U3494 ( .A1(n2103), .A2(\DataP/alu_a_in[7] ), .B1(
        \DataP/alu_a_in[8] ), .B2(n2916), .ZN(n2789) );
  AOI22_X1 U3495 ( .A1(n2103), .A2(n2207), .B1(\DataP/alu_a_in[10] ), .B2(
        n2916), .ZN(n2791) );
  AOI22_X1 U3496 ( .A1(n2917), .A2(n2789), .B1(n2791), .B2(n2105), .ZN(n2801)
         );
  AOI22_X1 U3497 ( .A1(n3202), .A2(n2798), .B1(n2801), .B2(n3052), .ZN(n2819)
         );
  AOI22_X1 U3498 ( .A1(n3204), .A2(n2820), .B1(n2819), .B2(n2101), .ZN(n2863)
         );
  AOI22_X1 U3499 ( .A1(n2103), .A2(n2231), .B1(n2232), .B2(n2916), .ZN(n2792)
         );
  AOI22_X1 U3500 ( .A1(n2103), .A2(\DataP/alu_a_in[2] ), .B1(n1973), .B2(n2118), .ZN(n2794) );
  AOI22_X1 U3501 ( .A1(n2917), .A2(n2792), .B1(n2794), .B2(n2105), .ZN(n2803)
         );
  NAND2_X1 U3502 ( .A1(n2918), .A2(n2803), .ZN(n2825) );
  AOI22_X1 U3503 ( .A1(n2103), .A2(\DataP/alu_a_in[4] ), .B1(
        \DataP/alu_a_in[5] ), .B2(n2916), .ZN(n2793) );
  AOI22_X1 U3504 ( .A1(n2103), .A2(\DataP/alu_a_in[6] ), .B1(
        \DataP/alu_a_in[7] ), .B2(n2916), .ZN(n2796) );
  AOI22_X1 U3505 ( .A1(n2917), .A2(n2793), .B1(n2796), .B2(n2105), .ZN(n2802)
         );
  AOI22_X1 U3506 ( .A1(n2103), .A2(\DataP/alu_a_in[8] ), .B1(n2207), .B2(n2916), .ZN(n2795) );
  AOI22_X1 U3507 ( .A1(n2103), .A2(\DataP/alu_a_in[10] ), .B1(n2200), .B2(
        n2118), .ZN(n2797) );
  AOI22_X1 U3508 ( .A1(n2917), .A2(n2795), .B1(n2797), .B2(n2105), .ZN(n2805)
         );
  AOI22_X1 U3509 ( .A1(n3202), .A2(n2802), .B1(n2805), .B2(n3053), .ZN(n2824)
         );
  AOI22_X1 U3510 ( .A1(n2115), .A2(n2825), .B1(n2824), .B2(n2101), .ZN(n2868)
         );
  NOR2_X1 U3511 ( .A1(n3055), .A2(n2903), .ZN(\DataP/ALU_C/shifter/N29 ) );
  NOR2_X1 U3512 ( .A1(n3050), .A2(n2785), .ZN(n2788) );
  AOI22_X1 U3513 ( .A1(n2917), .A2(n2787), .B1(n2786), .B2(n2105), .ZN(n2807)
         );
  AOI22_X1 U3514 ( .A1(n3202), .A2(n2788), .B1(n2807), .B2(n3052), .ZN(n2831)
         );
  AOI22_X1 U3515 ( .A1(n2917), .A2(n2790), .B1(n2789), .B2(n2105), .ZN(n2806)
         );
  AOI22_X1 U3516 ( .A1(n2103), .A2(n2200), .B1(\DataP/alu_a_in[12] ), .B2(
        n2118), .ZN(n2800) );
  AOI22_X1 U3517 ( .A1(n3049), .A2(n2791), .B1(n2800), .B2(n2105), .ZN(n2809)
         );
  AOI22_X1 U3518 ( .A1(n3051), .A2(n2806), .B1(n2809), .B2(n3052), .ZN(n2830)
         );
  AOI22_X1 U3519 ( .A1(n2115), .A2(n2831), .B1(n2830), .B2(n2101), .ZN(n2875)
         );
  NOR2_X1 U3520 ( .A1(n2917), .A2(n2792), .ZN(n2816) );
  AOI22_X1 U3521 ( .A1(n2917), .A2(n2794), .B1(n2793), .B2(n2105), .ZN(n2813)
         );
  AOI22_X1 U3522 ( .A1(n3051), .A2(n2816), .B1(n2813), .B2(n3052), .ZN(n2836)
         );
  AOI22_X1 U3523 ( .A1(n2917), .A2(n2796), .B1(n2795), .B2(n2105), .ZN(n2812)
         );
  AOI22_X1 U3524 ( .A1(n2103), .A2(\DataP/alu_a_in[12] ), .B1(
        \DataP/alu_a_in[13] ), .B2(n2118), .ZN(n2804) );
  AOI22_X1 U3525 ( .A1(n3050), .A2(n2797), .B1(n2804), .B2(n2105), .ZN(n2815)
         );
  AOI22_X1 U3526 ( .A1(n3202), .A2(n2812), .B1(n2815), .B2(n2919), .ZN(n2835)
         );
  AOI22_X1 U3527 ( .A1(n3204), .A2(n2836), .B1(n2835), .B2(n2101), .ZN(n2882)
         );
  AOI22_X1 U3528 ( .A1(n3202), .A2(n2799), .B1(n2798), .B2(n3053), .ZN(n2841)
         );
  AOI22_X1 U3529 ( .A1(n2103), .A2(\DataP/alu_a_in[13] ), .B1(
        \DataP/alu_a_in[14] ), .B2(n2118), .ZN(n2808) );
  AOI22_X1 U3530 ( .A1(n2917), .A2(n2800), .B1(n2808), .B2(n2105), .ZN(n2818)
         );
  AOI22_X1 U3531 ( .A1(n3202), .A2(n2801), .B1(n2818), .B2(n3053), .ZN(n2840)
         );
  AOI22_X1 U3532 ( .A1(n2115), .A2(n2841), .B1(n2840), .B2(n2101), .ZN(n2890)
         );
  NOR2_X1 U3533 ( .A1(n3055), .A2(n2906), .ZN(\DataP/ALU_C/shifter/N32 ) );
  AOI22_X1 U3534 ( .A1(n3202), .A2(n2803), .B1(n2802), .B2(n2919), .ZN(n2846)
         );
  AOI22_X1 U3535 ( .A1(n2103), .A2(\DataP/alu_a_in[14] ), .B1(
        \DataP/alu_a_in[15] ), .B2(n2118), .ZN(n2814) );
  AOI22_X1 U3536 ( .A1(n2917), .A2(n2804), .B1(n2814), .B2(n2105), .ZN(n2823)
         );
  AOI22_X1 U3537 ( .A1(n3202), .A2(n2805), .B1(n2823), .B2(n3053), .ZN(n2845)
         );
  AOI22_X1 U3538 ( .A1(n2115), .A2(n2846), .B1(n2845), .B2(n2101), .ZN(n2894)
         );
  NOR2_X1 U3539 ( .A1(n3055), .A2(n2907), .ZN(\DataP/ALU_C/shifter/N33 ) );
  AOI22_X1 U3540 ( .A1(n3202), .A2(n2807), .B1(n2806), .B2(n3053), .ZN(n2852)
         );
  AOI22_X1 U3541 ( .A1(n2103), .A2(\DataP/alu_a_in[15] ), .B1(
        \DataP/alu_a_in[16] ), .B2(n2118), .ZN(n2817) );
  AOI22_X1 U3542 ( .A1(n3049), .A2(n2808), .B1(n2817), .B2(n2105), .ZN(n2829)
         );
  AOI22_X1 U3543 ( .A1(n3202), .A2(n2809), .B1(n2829), .B2(n3053), .ZN(n2851)
         );
  AOI22_X1 U3544 ( .A1(n2115), .A2(n2852), .B1(n2851), .B2(n2101), .ZN(n2811)
         );
  MUX2_X1 U3545 ( .A(n2811), .B(n2810), .S(n2138), .Z(
        \DataP/ALU_C/shifter/N34 ) );
  AOI22_X1 U3546 ( .A1(n3202), .A2(n2813), .B1(n2812), .B2(n2919), .ZN(n2858)
         );
  AOI22_X1 U3547 ( .A1(n2103), .A2(\DataP/alu_a_in[16] ), .B1(n1751), .B2(
        n2118), .ZN(n2822) );
  AOI22_X1 U3548 ( .A1(n3049), .A2(n2814), .B1(n2822), .B2(n2105), .ZN(n2834)
         );
  AOI22_X1 U3549 ( .A1(n3202), .A2(n2815), .B1(n2834), .B2(n2919), .ZN(n2857)
         );
  NAND2_X1 U3550 ( .A1(n2816), .A2(n3053), .ZN(n2859) );
  NOR2_X1 U3551 ( .A1(n3204), .A2(n2859), .ZN(n2827) );
  AOI22_X1 U3552 ( .A1(n2226), .A2(n1751), .B1(\DataP/alu_a_in[18] ), .B2(
        n2118), .ZN(n2828) );
  AOI22_X1 U3553 ( .A1(n2917), .A2(n2817), .B1(n2828), .B2(n2105), .ZN(n2839)
         );
  AOI22_X1 U3554 ( .A1(n3202), .A2(n2818), .B1(n2839), .B2(n2919), .ZN(n2862)
         );
  AOI22_X1 U3555 ( .A1(n2115), .A2(n2819), .B1(n2862), .B2(n2101), .ZN(n2821)
         );
  NOR2_X1 U3556 ( .A1(n3204), .A2(n2820), .ZN(n2884) );
  MUX2_X1 U3557 ( .A(n2821), .B(n2884), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N36 ) );
  AOI22_X1 U3558 ( .A1(n2103), .A2(\DataP/alu_a_in[18] ), .B1(
        \DataP/alu_a_in[19] ), .B2(n2118), .ZN(n2833) );
  AOI22_X1 U3559 ( .A1(n2917), .A2(n2822), .B1(n2833), .B2(n2105), .ZN(n2844)
         );
  AOI22_X1 U3560 ( .A1(n3202), .A2(n2823), .B1(n2844), .B2(n2919), .ZN(n2867)
         );
  AOI22_X1 U3561 ( .A1(n2115), .A2(n2824), .B1(n2867), .B2(n2101), .ZN(n2826)
         );
  NOR2_X1 U3562 ( .A1(n3204), .A2(n2825), .ZN(n2895) );
  MUX2_X1 U3563 ( .A(n2826), .B(n2895), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N37 ) );
  NOR2_X1 U3564 ( .A1(n3055), .A2(n2908), .ZN(\DataP/ALU_C/shifter/N19 ) );
  AOI22_X1 U3565 ( .A1(n2103), .A2(\DataP/alu_a_in[19] ), .B1(
        \DataP/alu_a_in[20] ), .B2(n2118), .ZN(n2838) );
  AOI22_X1 U3566 ( .A1(n3050), .A2(n2828), .B1(n2838), .B2(n2105), .ZN(n2849)
         );
  AOI22_X1 U3567 ( .A1(n3202), .A2(n2829), .B1(n2849), .B2(n2919), .ZN(n2874)
         );
  AOI22_X1 U3568 ( .A1(n2115), .A2(n2830), .B1(n2874), .B2(n2101), .ZN(n2832)
         );
  NOR2_X1 U3569 ( .A1(n3204), .A2(n2831), .ZN(n2896) );
  MUX2_X1 U3570 ( .A(n2832), .B(n2896), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N38 ) );
  AOI22_X1 U3571 ( .A1(n2103), .A2(\DataP/alu_a_in[20] ), .B1(
        \DataP/alu_a_in[21] ), .B2(n2118), .ZN(n2843) );
  AOI22_X1 U3572 ( .A1(n3050), .A2(n2833), .B1(n2843), .B2(n2105), .ZN(n2856)
         );
  AOI22_X1 U3573 ( .A1(n3202), .A2(n2834), .B1(n2856), .B2(n2919), .ZN(n2881)
         );
  AOI22_X1 U3574 ( .A1(n2115), .A2(n2835), .B1(n2881), .B2(n2101), .ZN(n2837)
         );
  NOR2_X1 U3575 ( .A1(n3204), .A2(n2836), .ZN(n2897) );
  MUX2_X1 U3576 ( .A(n2837), .B(n2897), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N39 ) );
  AOI22_X1 U3577 ( .A1(n2103), .A2(\DataP/alu_a_in[21] ), .B1(
        \DataP/alu_a_in[22] ), .B2(n2118), .ZN(n2848) );
  AOI22_X1 U3578 ( .A1(n2917), .A2(n2838), .B1(n2848), .B2(n2105), .ZN(n2861)
         );
  AOI22_X1 U3579 ( .A1(n3202), .A2(n2839), .B1(n2861), .B2(n2919), .ZN(n2889)
         );
  AOI22_X1 U3580 ( .A1(n2115), .A2(n2840), .B1(n2889), .B2(n2101), .ZN(n2842)
         );
  NOR2_X1 U3581 ( .A1(n3204), .A2(n2841), .ZN(n2898) );
  MUX2_X1 U3582 ( .A(n2842), .B(n2898), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N40 ) );
  AOI22_X1 U3583 ( .A1(n2103), .A2(\DataP/alu_a_in[22] ), .B1(
        \DataP/alu_a_in[23] ), .B2(n2118), .ZN(n2855) );
  AOI22_X1 U3584 ( .A1(n2917), .A2(n2843), .B1(n2855), .B2(n2105), .ZN(n2865)
         );
  AOI22_X1 U3585 ( .A1(n3202), .A2(n2844), .B1(n2865), .B2(n2919), .ZN(n2893)
         );
  AOI22_X1 U3586 ( .A1(n2115), .A2(n2845), .B1(n2893), .B2(n2101), .ZN(n2847)
         );
  NOR2_X1 U3587 ( .A1(n3204), .A2(n2846), .ZN(n2899) );
  MUX2_X1 U3588 ( .A(n2847), .B(n2899), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N41 ) );
  AOI22_X1 U3589 ( .A1(n2103), .A2(\DataP/alu_a_in[23] ), .B1(
        \DataP/alu_a_in[24] ), .B2(n2118), .ZN(n2860) );
  AOI22_X1 U3590 ( .A1(n2917), .A2(n2848), .B1(n2860), .B2(n2105), .ZN(n2872)
         );
  AOI22_X1 U3591 ( .A1(n3202), .A2(n2849), .B1(n2872), .B2(n2919), .ZN(n2850)
         );
  AOI22_X1 U3592 ( .A1(n2115), .A2(n2851), .B1(n2850), .B2(n2101), .ZN(n2854)
         );
  AOI22_X1 U3593 ( .A1(n2115), .A2(n2853), .B1(n2852), .B2(n2101), .ZN(n2900)
         );
  MUX2_X1 U3594 ( .A(n2854), .B(n2900), .S(n2138), .Z(
        \DataP/ALU_C/shifter/N42 ) );
  AOI22_X1 U3595 ( .A1(n2103), .A2(\DataP/alu_a_in[24] ), .B1(
        \DataP/alu_a_in[25] ), .B2(n2118), .ZN(n2864) );
  AOI22_X1 U3596 ( .A1(n2917), .A2(n2855), .B1(n2864), .B2(n2105), .ZN(n2879)
         );
  AOI22_X1 U3597 ( .A1(n2115), .A2(n2859), .B1(n2858), .B2(n2101), .ZN(n2901)
         );
  AOI22_X1 U3598 ( .A1(n2103), .A2(\DataP/alu_a_in[25] ), .B1(
        \DataP/alu_a_in[26] ), .B2(n2118), .ZN(n2870) );
  AOI22_X1 U3599 ( .A1(n2917), .A2(n2860), .B1(n2870), .B2(n2105), .ZN(n2888)
         );
  AOI22_X1 U3600 ( .A1(n2103), .A2(\DataP/alu_a_in[26] ), .B1(
        \DataP/alu_a_in[27] ), .B2(n2118), .ZN(n2877) );
  AOI22_X1 U3601 ( .A1(n2917), .A2(n2864), .B1(n2877), .B2(n2105), .ZN(n2892)
         );
  AOI22_X1 U3602 ( .A1(n3202), .A2(n2865), .B1(n2892), .B2(n2918), .ZN(n2866)
         );
  AOI22_X1 U3603 ( .A1(n2115), .A2(n2867), .B1(n2866), .B2(n2101), .ZN(n2869)
         );
  MUX2_X1 U3604 ( .A(n2869), .B(n2868), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N45 ) );
  AOI22_X1 U3605 ( .A1(n2103), .A2(\DataP/alu_a_in[27] ), .B1(
        \DataP/alu_a_in[28] ), .B2(n2118), .ZN(n2886) );
  AOI22_X1 U3606 ( .A1(n2917), .A2(n2870), .B1(n2886), .B2(n2105), .ZN(n2871)
         );
  AOI22_X1 U3607 ( .A1(n3202), .A2(n2872), .B1(n2871), .B2(n2918), .ZN(n2873)
         );
  AOI22_X1 U3608 ( .A1(n2115), .A2(n2874), .B1(n2873), .B2(n2101), .ZN(n2876)
         );
  MUX2_X1 U3609 ( .A(n2876), .B(n2875), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N46 ) );
  AOI22_X1 U3610 ( .A1(n2103), .A2(\DataP/alu_a_in[28] ), .B1(
        \DataP/alu_a_in[29] ), .B2(n2118), .ZN(n2891) );
  AOI22_X1 U3611 ( .A1(n2917), .A2(n2877), .B1(n2891), .B2(n2105), .ZN(n2878)
         );
  AOI22_X1 U3612 ( .A1(n3051), .A2(n2879), .B1(n2878), .B2(n2918), .ZN(n2880)
         );
  AOI22_X1 U3613 ( .A1(n2115), .A2(n2881), .B1(n2880), .B2(n2101), .ZN(n2883)
         );
  MUX2_X1 U3614 ( .A(n2883), .B(n2882), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N47 ) );
  NOR2_X1 U3615 ( .A1(n2138), .A2(n2909), .ZN(\DataP/ALU_C/shifter/N20 ) );
  AOI22_X1 U3616 ( .A1(n2103), .A2(\DataP/alu_a_in[29] ), .B1(
        \DataP/alu_a_in[30] ), .B2(n2118), .ZN(n2885) );
  AOI22_X1 U3617 ( .A1(n2917), .A2(n2886), .B1(n2885), .B2(n2105), .ZN(n2887)
         );
  INV_X1 U3618 ( .A(n2126), .ZN(n2917) );
  AOI22_X1 U3619 ( .A1(n2103), .A2(\DataP/alu_a_in[15] ), .B1(
        \DataP/alu_a_in[14] ), .B2(n2117), .ZN(n2928) );
  AOI22_X1 U3620 ( .A1(n2103), .A2(\DataP/alu_a_in[13] ), .B1(
        \DataP/alu_a_in[12] ), .B2(n2117), .ZN(n2931) );
  AOI22_X1 U3621 ( .A1(n3049), .A2(n2928), .B1(n2931), .B2(n3047), .ZN(n2939)
         );
  AOI22_X1 U3622 ( .A1(n2103), .A2(n2200), .B1(\DataP/alu_a_in[10] ), .B2(
        n2117), .ZN(n2930) );
  AOI22_X1 U3623 ( .A1(n2103), .A2(\DataP/alu_a_in[9] ), .B1(
        \DataP/alu_a_in[8] ), .B2(n2117), .ZN(n3000) );
  AOI22_X1 U3624 ( .A1(n3050), .A2(n2930), .B1(n3000), .B2(n3047), .ZN(n3017)
         );
  AOI22_X1 U3625 ( .A1(n3051), .A2(n2939), .B1(n3017), .B2(n3053), .ZN(n3038)
         );
  AOI22_X1 U3626 ( .A1(n2103), .A2(\DataP/alu_a_in[7] ), .B1(
        \DataP/alu_a_in[6] ), .B2(n2117), .ZN(n2999) );
  AOI22_X1 U3627 ( .A1(n2103), .A2(\DataP/alu_a_in[5] ), .B1(
        \DataP/alu_a_in[4] ), .B2(n2117), .ZN(n3002) );
  AOI22_X1 U3628 ( .A1(n3049), .A2(n2999), .B1(n3002), .B2(n3047), .ZN(n3016)
         );
  AOI22_X1 U3629 ( .A1(n2103), .A2(n1973), .B1(\DataP/alu_a_in[2] ), .B2(n2117), .ZN(n3001) );
  AOI22_X1 U3630 ( .A1(n2103), .A2(n2232), .B1(n2231), .B2(n2117), .ZN(n2920)
         );
  AOI221_X1 U3631 ( .B1(n3001), .B2(n3050), .C1(n2920), .C2(n3047), .A(n3051), 
        .ZN(n2921) );
  AOI21_X1 U3632 ( .B1(n3051), .B2(n3016), .A(n2921), .ZN(n2922) );
  AOI22_X1 U3633 ( .A1(n3204), .A2(n3038), .B1(n2922), .B2(n2101), .ZN(n2923)
         );
  AOI22_X1 U3634 ( .A1(n2226), .A2(\DataP/alu_a_in[31] ), .B1(
        \DataP/alu_a_in[30] ), .B2(n2117), .ZN(n2932) );
  AOI22_X1 U3635 ( .A1(n2226), .A2(\DataP/alu_a_in[29] ), .B1(
        \DataP/alu_a_in[28] ), .B2(n2117), .ZN(n2934) );
  AOI22_X1 U3636 ( .A1(n3049), .A2(n2932), .B1(n2934), .B2(n3201), .ZN(n2982)
         );
  AOI22_X1 U3637 ( .A1(n2103), .A2(\DataP/alu_a_in[27] ), .B1(
        \DataP/alu_a_in[26] ), .B2(n2117), .ZN(n2933) );
  AOI22_X1 U3638 ( .A1(n2226), .A2(\DataP/alu_a_in[25] ), .B1(
        \DataP/alu_a_in[24] ), .B2(n2117), .ZN(n2925) );
  AOI22_X1 U3639 ( .A1(n3049), .A2(n2933), .B1(n2925), .B2(n3201), .ZN(n2938)
         );
  AOI22_X1 U3640 ( .A1(n3202), .A2(n2982), .B1(n2938), .B2(n3052), .ZN(n2993)
         );
  AOI22_X1 U3641 ( .A1(n2103), .A2(\DataP/alu_a_in[23] ), .B1(
        \DataP/alu_a_in[22] ), .B2(n2117), .ZN(n2924) );
  AOI22_X1 U3642 ( .A1(n2226), .A2(\DataP/alu_a_in[21] ), .B1(
        \DataP/alu_a_in[20] ), .B2(n2117), .ZN(n2927) );
  AOI22_X1 U3643 ( .A1(n3050), .A2(n2924), .B1(n2927), .B2(n3047), .ZN(n2937)
         );
  AOI22_X1 U3644 ( .A1(n2103), .A2(\DataP/alu_a_in[19] ), .B1(
        \DataP/alu_a_in[18] ), .B2(n2117), .ZN(n2926) );
  AOI22_X1 U3645 ( .A1(n2226), .A2(\DataP/alu_a_in[17] ), .B1(
        \DataP/alu_a_in[16] ), .B2(n2117), .ZN(n2929) );
  AOI22_X1 U3646 ( .A1(n3050), .A2(n2926), .B1(n2929), .B2(n3047), .ZN(n2940)
         );
  AOI22_X1 U3647 ( .A1(n3202), .A2(n2937), .B1(n2940), .B2(n3052), .ZN(n3039)
         );
  AOI22_X1 U3648 ( .A1(n2112), .A2(n2993), .B1(n3039), .B2(n2101), .ZN(n2966)
         );
  MUX2_X1 U3649 ( .A(n2923), .B(n2966), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N50 ) );
  AOI22_X1 U3650 ( .A1(n3049), .A2(n2925), .B1(n2924), .B2(n3047), .ZN(n2954)
         );
  AOI22_X1 U3651 ( .A1(n3049), .A2(n2927), .B1(n2926), .B2(n3047), .ZN(n2957)
         );
  AOI22_X1 U3652 ( .A1(n3202), .A2(n2954), .B1(n2957), .B2(n3052), .ZN(n2971)
         );
  AOI22_X1 U3653 ( .A1(n3050), .A2(n2929), .B1(n2928), .B2(n3047), .ZN(n2956)
         );
  AOI22_X1 U3654 ( .A1(n3049), .A2(n2931), .B1(n2930), .B2(n3201), .ZN(n3028)
         );
  AOI22_X1 U3655 ( .A1(n3202), .A2(n2956), .B1(n3028), .B2(n3052), .ZN(n3005)
         );
  AOI22_X1 U3656 ( .A1(n2112), .A2(n2971), .B1(n3005), .B2(n2101), .ZN(n2935)
         );
  NOR2_X1 U3657 ( .A1(n3050), .A2(n2932), .ZN(n2987) );
  AOI22_X1 U3658 ( .A1(n3050), .A2(n2934), .B1(n2933), .B2(n3201), .ZN(n2955)
         );
  AOI22_X1 U3659 ( .A1(n3202), .A2(n2987), .B1(n2955), .B2(n3052), .ZN(n2972)
         );
  NOR2_X1 U3660 ( .A1(n2112), .A2(n2972), .ZN(n2995) );
  AOI22_X1 U3661 ( .A1(n2103), .A2(\DataP/alu_a_in[26] ), .B1(
        \DataP/alu_a_in[25] ), .B2(n2117), .ZN(n2943) );
  AOI22_X1 U3662 ( .A1(n2103), .A2(\DataP/alu_a_in[24] ), .B1(
        \DataP/alu_a_in[23] ), .B2(n2117), .ZN(n2946) );
  AOI22_X1 U3663 ( .A1(n3049), .A2(n2943), .B1(n2946), .B2(n3047), .ZN(n2960)
         );
  AOI22_X1 U3664 ( .A1(n2103), .A2(\DataP/alu_a_in[22] ), .B1(
        \DataP/alu_a_in[21] ), .B2(n2117), .ZN(n2945) );
  AOI22_X1 U3665 ( .A1(n2103), .A2(\DataP/alu_a_in[20] ), .B1(
        \DataP/alu_a_in[19] ), .B2(n2117), .ZN(n2948) );
  AOI22_X1 U3666 ( .A1(n3050), .A2(n2945), .B1(n2948), .B2(n3047), .ZN(n2963)
         );
  AOI22_X1 U3667 ( .A1(n3202), .A2(n2960), .B1(n2963), .B2(n3053), .ZN(n2973)
         );
  AOI22_X1 U3668 ( .A1(n2103), .A2(\DataP/alu_a_in[18] ), .B1(
        \DataP/alu_a_in[17] ), .B2(n2117), .ZN(n2947) );
  AOI22_X1 U3669 ( .A1(n2103), .A2(\DataP/alu_a_in[16] ), .B1(
        \DataP/alu_a_in[15] ), .B2(n2117), .ZN(n2950) );
  AOI22_X1 U3670 ( .A1(n3048), .A2(n2947), .B1(n2950), .B2(n3201), .ZN(n2962)
         );
  AOI22_X1 U3671 ( .A1(n2103), .A2(\DataP/alu_a_in[14] ), .B1(
        \DataP/alu_a_in[13] ), .B2(n2117), .ZN(n2949) );
  AOI22_X1 U3672 ( .A1(n2103), .A2(\DataP/alu_a_in[12] ), .B1(n2200), .B2(
        n2117), .ZN(n2975) );
  AOI22_X1 U3673 ( .A1(n3048), .A2(n2949), .B1(n2975), .B2(n3201), .ZN(n3034)
         );
  AOI22_X1 U3674 ( .A1(n3202), .A2(n2962), .B1(n3034), .B2(n3053), .ZN(n3014)
         );
  AOI22_X1 U3675 ( .A1(n2112), .A2(n2973), .B1(n3014), .B2(n2101), .ZN(n2936)
         );
  NAND2_X1 U3676 ( .A1(\DataP/alu_a_in[31] ), .A2(n2117), .ZN(n2952) );
  NOR2_X1 U3677 ( .A1(n3050), .A2(n2952), .ZN(n2990) );
  AOI22_X1 U3678 ( .A1(n2103), .A2(\DataP/alu_a_in[30] ), .B1(
        \DataP/alu_a_in[29] ), .B2(n2117), .ZN(n2951) );
  AOI22_X1 U3679 ( .A1(n2103), .A2(\DataP/alu_a_in[28] ), .B1(
        \DataP/alu_a_in[27] ), .B2(n2117), .ZN(n2944) );
  AOI22_X1 U3680 ( .A1(n3049), .A2(n2951), .B1(n2944), .B2(n3047), .ZN(n2961)
         );
  AOI22_X1 U3681 ( .A1(n3202), .A2(n2990), .B1(n2961), .B2(n3052), .ZN(n2974)
         );
  NOR2_X1 U3682 ( .A1(n2112), .A2(n2974), .ZN(n2996) );
  MUX2_X1 U3683 ( .A(n2936), .B(n2996), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N61 ) );
  NAND3_X1 U3684 ( .A1(n2101), .A2(n3052), .A3(n2982), .ZN(n2997) );
  AOI22_X1 U3685 ( .A1(n3202), .A2(n2938), .B1(n2937), .B2(n3053), .ZN(n2983)
         );
  AOI22_X1 U3686 ( .A1(n3202), .A2(n2940), .B1(n2939), .B2(n3053), .ZN(n3018)
         );
  AOI22_X1 U3687 ( .A1(n2112), .A2(n2983), .B1(n3018), .B2(n2101), .ZN(n2941)
         );
  NAND2_X1 U3688 ( .A1(n2102), .A2(n2941), .ZN(n2942) );
  AOI22_X1 U3689 ( .A1(n3049), .A2(n2944), .B1(n2943), .B2(n3047), .ZN(n2967)
         );
  AOI22_X1 U3690 ( .A1(n3050), .A2(n2946), .B1(n2945), .B2(n3201), .ZN(n2970)
         );
  AOI22_X1 U3691 ( .A1(n3051), .A2(n2967), .B1(n2970), .B2(n3053), .ZN(n2985)
         );
  AOI22_X1 U3692 ( .A1(n3048), .A2(n2948), .B1(n2947), .B2(n3047), .ZN(n2969)
         );
  AOI22_X1 U3693 ( .A1(n3048), .A2(n2950), .B1(n2949), .B2(n3201), .ZN(n2976)
         );
  AOI22_X1 U3694 ( .A1(n3051), .A2(n2969), .B1(n2976), .B2(n3053), .ZN(n3024)
         );
  AOI22_X1 U3695 ( .A1(n2112), .A2(n2985), .B1(n3024), .B2(n2101), .ZN(n2953)
         );
  AOI22_X1 U3696 ( .A1(n3049), .A2(n2952), .B1(n2951), .B2(n3201), .ZN(n2968)
         );
  NAND2_X1 U3697 ( .A1(n3052), .A2(n2968), .ZN(n2986) );
  NOR2_X1 U3698 ( .A1(n2112), .A2(n2986), .ZN(n2998) );
  NAND3_X1 U3699 ( .A1(n2987), .A2(n2101), .A3(n3053), .ZN(n3008) );
  AOI22_X1 U3700 ( .A1(n3051), .A2(n2955), .B1(n2954), .B2(n3053), .ZN(n2988)
         );
  AOI22_X1 U3701 ( .A1(n3051), .A2(n2957), .B1(n2956), .B2(n3053), .ZN(n3030)
         );
  AOI22_X1 U3702 ( .A1(n2112), .A2(n2988), .B1(n3030), .B2(n2101), .ZN(n2958)
         );
  NAND2_X1 U3703 ( .A1(n3206), .A2(n2958), .ZN(n2959) );
  OAI21_X1 U3704 ( .B1(n2102), .B2(n3008), .A(n2959), .ZN(
        \DataP/ALU_C/shifter/N64 ) );
  NAND3_X1 U3705 ( .A1(n2990), .A2(n2101), .A3(n3052), .ZN(n3009) );
  AOI22_X1 U3706 ( .A1(n3051), .A2(n2961), .B1(n2960), .B2(n3053), .ZN(n2991)
         );
  AOI22_X1 U3707 ( .A1(n3051), .A2(n2963), .B1(n2962), .B2(n3053), .ZN(n3035)
         );
  AOI22_X1 U3708 ( .A1(n2115), .A2(n2991), .B1(n3035), .B2(n2101), .ZN(n2964)
         );
  NAND2_X1 U3709 ( .A1(n2102), .A2(n2964), .ZN(n2965) );
  OAI21_X1 U3710 ( .B1(n3206), .B2(n3009), .A(n2965), .ZN(
        \DataP/ALU_C/shifter/N65 ) );
  AND2_X1 U3711 ( .A1(n3206), .A2(n2966), .ZN(\DataP/ALU_C/shifter/N66 ) );
  AOI22_X1 U3712 ( .A1(n3202), .A2(n2968), .B1(n2967), .B2(n3053), .ZN(n2994)
         );
  AOI22_X1 U3713 ( .A1(n3202), .A2(n2970), .B1(n2969), .B2(n3052), .ZN(n3043)
         );
  AOI22_X1 U3714 ( .A1(n3204), .A2(n2994), .B1(n3043), .B2(n2101), .ZN(n2980)
         );
  AND2_X1 U3715 ( .A1(n3206), .A2(n2980), .ZN(\DataP/ALU_C/shifter/N67 ) );
  AOI22_X1 U3716 ( .A1(n3204), .A2(n2972), .B1(n2971), .B2(n2101), .ZN(n3006)
         );
  AOI22_X1 U3717 ( .A1(n2115), .A2(n2974), .B1(n2973), .B2(n2101), .ZN(n3015)
         );
  AND2_X1 U3718 ( .A1(n2102), .A2(n3015), .ZN(\DataP/ALU_C/shifter/N69 ) );
  AOI22_X1 U3719 ( .A1(n2103), .A2(\DataP/alu_a_in[10] ), .B1(n2207), .B2(
        n2117), .ZN(n3011) );
  AOI22_X1 U3720 ( .A1(n3050), .A2(n2975), .B1(n3011), .B2(n3047), .ZN(n3022)
         );
  AOI22_X1 U3721 ( .A1(n3202), .A2(n2976), .B1(n3022), .B2(n3053), .ZN(n3042)
         );
  AOI22_X1 U3722 ( .A1(n2103), .A2(\DataP/alu_a_in[8] ), .B1(
        \DataP/alu_a_in[7] ), .B2(n2117), .ZN(n3010) );
  AOI22_X1 U3723 ( .A1(n2103), .A2(\DataP/alu_a_in[6] ), .B1(
        \DataP/alu_a_in[5] ), .B2(n2117), .ZN(n3013) );
  AOI22_X1 U3724 ( .A1(n3048), .A2(n3010), .B1(n3013), .B2(n3047), .ZN(n3021)
         );
  AOI22_X1 U3725 ( .A1(n2103), .A2(\DataP/alu_a_in[4] ), .B1(n1973), .B2(n2117), .ZN(n3012) );
  AOI22_X1 U3726 ( .A1(n2103), .A2(\DataP/alu_a_in[2] ), .B1(n2232), .B2(n2117), .ZN(n2977) );
  AOI22_X1 U3727 ( .A1(n3049), .A2(n3012), .B1(n2977), .B2(n3201), .ZN(n2978)
         );
  AOI22_X1 U3728 ( .A1(n3202), .A2(n3021), .B1(n2978), .B2(n3052), .ZN(n2979)
         );
  AOI22_X1 U3729 ( .A1(n3204), .A2(n3042), .B1(n2979), .B2(n2101), .ZN(n2981)
         );
  MUX2_X1 U3730 ( .A(n2981), .B(n2980), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N51 ) );
  NAND2_X1 U3731 ( .A1(n3052), .A2(n2982), .ZN(n2984) );
  AOI22_X1 U3732 ( .A1(n3204), .A2(n2984), .B1(n2983), .B2(n2101), .ZN(n3019)
         );
  AND2_X1 U3733 ( .A1(n2102), .A2(n3019), .ZN(\DataP/ALU_C/shifter/N70 ) );
  AOI22_X1 U3734 ( .A1(n3204), .A2(n2986), .B1(n2985), .B2(n2101), .ZN(n3025)
         );
  AND2_X1 U3735 ( .A1(n3206), .A2(n3025), .ZN(\DataP/ALU_C/shifter/N71 ) );
  NAND2_X1 U3736 ( .A1(n2987), .A2(n3052), .ZN(n2989) );
  AOI22_X1 U3737 ( .A1(n3204), .A2(n2989), .B1(n2988), .B2(n2101), .ZN(n3031)
         );
  AND2_X1 U3738 ( .A1(n3206), .A2(n3031), .ZN(\DataP/ALU_C/shifter/N72 ) );
  NAND2_X1 U3739 ( .A1(n2990), .A2(n3053), .ZN(n2992) );
  AOI22_X1 U3740 ( .A1(n3204), .A2(n2992), .B1(n2991), .B2(n2101), .ZN(n3036)
         );
  AND2_X1 U3741 ( .A1(n3206), .A2(n3036), .ZN(\DataP/ALU_C/shifter/N73 ) );
  NOR2_X1 U3742 ( .A1(n2112), .A2(n2993), .ZN(n3040) );
  AND2_X1 U3743 ( .A1(n3040), .A2(n3206), .ZN(\DataP/ALU_C/shifter/N74 ) );
  NOR2_X1 U3744 ( .A1(n2112), .A2(n2994), .ZN(n3044) );
  AND2_X1 U3745 ( .A1(n3044), .A2(n2102), .ZN(\DataP/ALU_C/shifter/N75 ) );
  AND2_X1 U3746 ( .A1(n2995), .A2(n2102), .ZN(\DataP/ALU_C/shifter/N76 ) );
  AND2_X1 U3747 ( .A1(n2996), .A2(n2102), .ZN(\DataP/ALU_C/shifter/N77 ) );
  NOR2_X1 U3748 ( .A1(n3055), .A2(n2997), .ZN(\DataP/ALU_C/shifter/N78 ) );
  AND2_X1 U3749 ( .A1(n2998), .A2(n2102), .ZN(\DataP/ALU_C/shifter/N79 ) );
  AOI22_X1 U3750 ( .A1(n3048), .A2(n3000), .B1(n2999), .B2(n3201), .ZN(n3027)
         );
  AOI22_X1 U3751 ( .A1(n3048), .A2(n3002), .B1(n3001), .B2(n3047), .ZN(n3003)
         );
  AOI22_X1 U3752 ( .A1(n3202), .A2(n3027), .B1(n3003), .B2(n3052), .ZN(n3004)
         );
  AOI22_X1 U3753 ( .A1(n2115), .A2(n3005), .B1(n3004), .B2(n2101), .ZN(n3007)
         );
  MUX2_X1 U3754 ( .A(n3007), .B(n3006), .S(n2138), .Z(
        \DataP/ALU_C/shifter/N52 ) );
  NOR2_X1 U3755 ( .A1(n2138), .A2(n3008), .ZN(\DataP/ALU_C/shifter/N80 ) );
  NOR2_X1 U3756 ( .A1(n3055), .A2(n3009), .ZN(\DataP/ALU_C/shifter/N81 ) );
  AOI22_X1 U3757 ( .A1(n3049), .A2(n3011), .B1(n3010), .B2(n3047), .ZN(n3033)
         );
  AOI22_X1 U3758 ( .A1(n3051), .A2(n3022), .B1(n3021), .B2(n3052), .ZN(n3023)
         );
  AOI22_X1 U3759 ( .A1(n2112), .A2(n3024), .B1(n3023), .B2(n2101), .ZN(n3026)
         );
  AOI22_X1 U3760 ( .A1(n3051), .A2(n3028), .B1(n3027), .B2(n3052), .ZN(n3029)
         );
  AOI22_X1 U3761 ( .A1(n2112), .A2(n3030), .B1(n3029), .B2(n2101), .ZN(n3032)
         );
  AOI22_X1 U3762 ( .A1(n2112), .A2(n3039), .B1(n3038), .B2(n2101), .ZN(n3041)
         );
  AOI22_X1 U3763 ( .A1(n2112), .A2(n3043), .B1(n3042), .B2(n2101), .ZN(n3045)
         );
  MUX2_X1 U3764 ( .A(n3045), .B(n3044), .S(n3055), .Z(
        \DataP/ALU_C/shifter/N59 ) );
  INV_X1 U3765 ( .A(n3200), .ZN(n3049) );
  INV_X1 U3766 ( .A(n3200), .ZN(n3050) );
  AOI22_X1 U3767 ( .A1(n2103), .A2(\DataP/alu_a_in[31] ), .B1(
        \DataP/alu_a_in[30] ), .B2(n3199), .ZN(n3060) );
  AOI22_X1 U3768 ( .A1(n2103), .A2(\DataP/alu_a_in[29] ), .B1(
        \DataP/alu_a_in[28] ), .B2(n3199), .ZN(n3062) );
  AOI22_X1 U3769 ( .A1(n3048), .A2(n3060), .B1(n3062), .B2(n3047), .ZN(n3073)
         );
  AOI22_X1 U3770 ( .A1(n2103), .A2(\DataP/alu_a_in[27] ), .B1(
        \DataP/alu_a_in[26] ), .B2(n3199), .ZN(n3061) );
  AOI22_X1 U3771 ( .A1(n2103), .A2(\DataP/alu_a_in[25] ), .B1(
        \DataP/alu_a_in[24] ), .B2(n3199), .ZN(n3064) );
  AOI22_X1 U3772 ( .A1(n3048), .A2(n3061), .B1(n3064), .B2(n3201), .ZN(n3075)
         );
  AOI22_X1 U3773 ( .A1(n3202), .A2(n3073), .B1(n3075), .B2(n3053), .ZN(n3126)
         );
  AOI22_X1 U3774 ( .A1(n2103), .A2(\DataP/alu_a_in[23] ), .B1(
        \DataP/alu_a_in[22] ), .B2(n3199), .ZN(n3063) );
  AOI22_X1 U3775 ( .A1(n2103), .A2(\DataP/alu_a_in[21] ), .B1(
        \DataP/alu_a_in[20] ), .B2(n3199), .ZN(n3066) );
  AOI22_X1 U3776 ( .A1(n3048), .A2(n3063), .B1(n3066), .B2(n3047), .ZN(n3074)
         );
  AOI22_X1 U3777 ( .A1(n2103), .A2(\DataP/alu_a_in[19] ), .B1(
        \DataP/alu_a_in[18] ), .B2(n3199), .ZN(n3065) );
  AOI22_X1 U3778 ( .A1(n2103), .A2(n1751), .B1(\DataP/alu_a_in[16] ), .B2(
        n3199), .ZN(n3068) );
  AOI22_X1 U3779 ( .A1(n3048), .A2(n3065), .B1(n3068), .B2(n3047), .ZN(n3077)
         );
  AOI22_X1 U3780 ( .A1(n3203), .A2(n3074), .B1(n3077), .B2(n2918), .ZN(n3189)
         );
  AOI22_X1 U3781 ( .A1(n3205), .A2(n3126), .B1(n3189), .B2(n2101), .ZN(n3101)
         );
  AOI22_X1 U3782 ( .A1(n2103), .A2(\DataP/alu_a_in[15] ), .B1(
        \DataP/alu_a_in[14] ), .B2(n3199), .ZN(n3067) );
  AOI22_X1 U3783 ( .A1(n2103), .A2(\DataP/alu_a_in[13] ), .B1(
        \DataP/alu_a_in[12] ), .B2(n3199), .ZN(n3070) );
  AOI22_X1 U3784 ( .A1(n3049), .A2(n3067), .B1(n3070), .B2(n3201), .ZN(n3076)
         );
  AOI22_X1 U3785 ( .A1(n2103), .A2(n2200), .B1(\DataP/alu_a_in[10] ), .B2(
        n2916), .ZN(n3069) );
  AOI22_X1 U3786 ( .A1(n2103), .A2(n2207), .B1(\DataP/alu_a_in[8] ), .B2(n2916), .ZN(n3141) );
  AOI22_X1 U3787 ( .A1(n3048), .A2(n3069), .B1(n3141), .B2(n3047), .ZN(n3162)
         );
  AOI22_X1 U3788 ( .A1(n3203), .A2(n3076), .B1(n3162), .B2(n2918), .ZN(n3188)
         );
  AOI22_X1 U3789 ( .A1(n2103), .A2(\DataP/alu_a_in[7] ), .B1(
        \DataP/alu_a_in[6] ), .B2(n3199), .ZN(n3140) );
  AOI22_X1 U3790 ( .A1(n2103), .A2(\DataP/alu_a_in[5] ), .B1(
        \DataP/alu_a_in[4] ), .B2(n2916), .ZN(n3143) );
  AOI22_X1 U3791 ( .A1(n3050), .A2(n3140), .B1(n3143), .B2(n3047), .ZN(n3161)
         );
  AOI22_X1 U3792 ( .A1(n2103), .A2(n1973), .B1(\DataP/alu_a_in[2] ), .B2(n3199), .ZN(n3142) );
  AOI22_X1 U3793 ( .A1(n2103), .A2(n2232), .B1(n2201), .B2(n2916), .ZN(n3056)
         );
  AOI221_X1 U3794 ( .B1(n3142), .B2(n3050), .C1(n3056), .C2(n3047), .A(n3202), 
        .ZN(n3057) );
  AOI21_X1 U3795 ( .B1(n3202), .B2(n3161), .A(n3057), .ZN(n3058) );
  AOI22_X1 U3796 ( .A1(n3205), .A2(n3188), .B1(n3058), .B2(n2101), .ZN(n3059)
         );
  MUX2_X1 U3797 ( .A(n3101), .B(n3059), .S(n3206), .Z(
        \DataP/ALU_C/shifter/N82 ) );
  AOI22_X1 U3798 ( .A1(n3050), .A2(n2073), .B1(n3060), .B2(n3047), .ZN(n3090)
         );
  AOI22_X1 U3799 ( .A1(n3048), .A2(n3062), .B1(n3061), .B2(n3047), .ZN(n3092)
         );
  AOI22_X1 U3800 ( .A1(n3203), .A2(n3090), .B1(n3092), .B2(n2918), .ZN(n3107)
         );
  NAND2_X1 U3801 ( .A1(n3204), .A2(\DataP/alu_a_in[31] ), .ZN(n3128) );
  OAI21_X1 U3802 ( .B1(n3205), .B2(n3107), .A(n3128), .ZN(n3132) );
  AOI22_X1 U3803 ( .A1(n3049), .A2(n3064), .B1(n3063), .B2(n3047), .ZN(n3091)
         );
  AOI22_X1 U3804 ( .A1(n3049), .A2(n3066), .B1(n3065), .B2(n3201), .ZN(n3094)
         );
  AOI22_X1 U3805 ( .A1(n3202), .A2(n3091), .B1(n3094), .B2(n2918), .ZN(n3106)
         );
  AOI22_X1 U3806 ( .A1(n3050), .A2(n3068), .B1(n3067), .B2(n3047), .ZN(n3093)
         );
  AOI22_X1 U3807 ( .A1(n3048), .A2(n3070), .B1(n3069), .B2(n3201), .ZN(n3176)
         );
  AOI22_X1 U3808 ( .A1(n3202), .A2(n3093), .B1(n3176), .B2(n2918), .ZN(n3146)
         );
  AOI22_X1 U3809 ( .A1(n3205), .A2(n3106), .B1(n3146), .B2(n2101), .ZN(n3071)
         );
  AOI22_X1 U3810 ( .A1(n2103), .A2(\DataP/alu_a_in[30] ), .B1(
        \DataP/alu_a_in[29] ), .B2(n2916), .ZN(n3079) );
  AOI22_X1 U3811 ( .A1(n2103), .A2(\DataP/alu_a_in[28] ), .B1(
        \DataP/alu_a_in[27] ), .B2(n3199), .ZN(n3081) );
  AOI22_X1 U3812 ( .A1(n3050), .A2(n3079), .B1(n3081), .B2(n3047), .ZN(n3097)
         );
  NOR2_X1 U3813 ( .A1(n3052), .A2(n2073), .ZN(n3089) );
  AOI21_X1 U3814 ( .B1(n2919), .B2(n3097), .A(n3089), .ZN(n3109) );
  OAI21_X1 U3815 ( .B1(n3205), .B2(n3109), .A(n3128), .ZN(n3134) );
  AOI22_X1 U3816 ( .A1(n2103), .A2(\DataP/alu_a_in[26] ), .B1(
        \DataP/alu_a_in[25] ), .B2(n2916), .ZN(n3080) );
  AOI22_X1 U3817 ( .A1(n2103), .A2(\DataP/alu_a_in[24] ), .B1(
        \DataP/alu_a_in[23] ), .B2(n3199), .ZN(n3083) );
  AOI22_X1 U3818 ( .A1(n3048), .A2(n3080), .B1(n3083), .B2(n3047), .ZN(n3096)
         );
  AOI22_X1 U3819 ( .A1(n2103), .A2(\DataP/alu_a_in[22] ), .B1(
        \DataP/alu_a_in[21] ), .B2(n3199), .ZN(n3082) );
  AOI22_X1 U3820 ( .A1(n2103), .A2(\DataP/alu_a_in[20] ), .B1(
        \DataP/alu_a_in[19] ), .B2(n3199), .ZN(n3085) );
  AOI22_X1 U3821 ( .A1(n3049), .A2(n3082), .B1(n3085), .B2(n3047), .ZN(n3099)
         );
  AOI22_X1 U3822 ( .A1(n3202), .A2(n3096), .B1(n3099), .B2(n2919), .ZN(n3108)
         );
  AOI22_X1 U3823 ( .A1(n2103), .A2(\DataP/alu_a_in[18] ), .B1(n1751), .B2(
        n3199), .ZN(n3084) );
  AOI22_X1 U3824 ( .A1(n2103), .A2(\DataP/alu_a_in[16] ), .B1(
        \DataP/alu_a_in[15] ), .B2(n2916), .ZN(n3087) );
  AOI22_X1 U3825 ( .A1(n3050), .A2(n3084), .B1(n3087), .B2(n3047), .ZN(n3098)
         );
  AOI22_X1 U3826 ( .A1(n2103), .A2(\DataP/alu_a_in[14] ), .B1(
        \DataP/alu_a_in[13] ), .B2(n3199), .ZN(n3086) );
  AOI22_X1 U3827 ( .A1(n2103), .A2(\DataP/alu_a_in[12] ), .B1(n2200), .B2(
        n2916), .ZN(n3110) );
  AOI22_X1 U3828 ( .A1(n3048), .A2(n3086), .B1(n3110), .B2(n3047), .ZN(n3183)
         );
  AOI22_X1 U3829 ( .A1(n3202), .A2(n3098), .B1(n3183), .B2(n2919), .ZN(n3157)
         );
  AOI22_X1 U3830 ( .A1(n3205), .A2(n3108), .B1(n3157), .B2(n2101), .ZN(n3072)
         );
  MUX2_X1 U3831 ( .A(n3134), .B(n3072), .S(n3206), .Z(
        \DataP/ALU_C/shifter/N93 ) );
  AOI21_X1 U3832 ( .B1(n2919), .B2(n3073), .A(n3089), .ZN(n3119) );
  OAI21_X1 U3833 ( .B1(n3205), .B2(n3119), .A(n3128), .ZN(n3136) );
  AOI22_X1 U3834 ( .A1(n3202), .A2(n3075), .B1(n3074), .B2(n2918), .ZN(n3118)
         );
  AOI22_X1 U3835 ( .A1(n3202), .A2(n3077), .B1(n3076), .B2(n2918), .ZN(n3164)
         );
  AOI22_X1 U3836 ( .A1(n3205), .A2(n3118), .B1(n3164), .B2(n2101), .ZN(n3078)
         );
  AOI22_X1 U3837 ( .A1(n3050), .A2(n2073), .B1(n3079), .B2(n3047), .ZN(n3103)
         );
  AOI21_X1 U3838 ( .B1(n2918), .B2(n3103), .A(n3089), .ZN(n3121) );
  OAI21_X1 U3839 ( .B1(n3204), .B2(n3121), .A(n3128), .ZN(n3138) );
  AOI22_X1 U3840 ( .A1(n3050), .A2(n3081), .B1(n3080), .B2(n3047), .ZN(n3102)
         );
  AOI22_X1 U3841 ( .A1(n3050), .A2(n3083), .B1(n3082), .B2(n3047), .ZN(n3105)
         );
  AOI22_X1 U3842 ( .A1(n3202), .A2(n3102), .B1(n3105), .B2(n3052), .ZN(n3120)
         );
  AOI22_X1 U3843 ( .A1(n3048), .A2(n3085), .B1(n3084), .B2(n3047), .ZN(n3104)
         );
  AOI22_X1 U3844 ( .A1(n3048), .A2(n3087), .B1(n3086), .B2(n3047), .ZN(n3111)
         );
  AOI22_X1 U3845 ( .A1(n3202), .A2(n3104), .B1(n3111), .B2(n3052), .ZN(n3171)
         );
  AOI22_X1 U3846 ( .A1(n3205), .A2(n3120), .B1(n3171), .B2(n2101), .ZN(n3088)
         );
  AOI21_X1 U3847 ( .B1(n3053), .B2(n3090), .A(n3089), .ZN(n3123) );
  OAI21_X1 U3848 ( .B1(n3204), .B2(n3123), .A(n3128), .ZN(n3150) );
  AOI22_X1 U3849 ( .A1(n3202), .A2(n3092), .B1(n3091), .B2(n2919), .ZN(n3122)
         );
  AOI22_X1 U3850 ( .A1(n3202), .A2(n3094), .B1(n3093), .B2(n2918), .ZN(n3178)
         );
  AOI22_X1 U3851 ( .A1(n3205), .A2(n3122), .B1(n3178), .B2(n2101), .ZN(n3095)
         );
  MUX2_X1 U3852 ( .A(n3150), .B(n3095), .S(n2102), .Z(
        \DataP/ALU_C/shifter/N96 ) );
  NAND2_X1 U3853 ( .A1(n3055), .A2(\DataP/alu_a_in[31] ), .ZN(n3131) );
  AOI22_X1 U3854 ( .A1(n3202), .A2(n3097), .B1(n3096), .B2(n2918), .ZN(n3124)
         );
  AOI22_X1 U3855 ( .A1(n3202), .A2(n3099), .B1(n3098), .B2(n3053), .ZN(n3185)
         );
  AOI221_X1 U3856 ( .B1(n3124), .B2(n3204), .C1(n3185), .C2(n2101), .A(n3055), 
        .ZN(n3100) );
  OR2_X1 U3857 ( .A1(n3195), .A2(n3100), .ZN(\DataP/ALU_C/shifter/N97 ) );
  AOI22_X1 U3858 ( .A1(n3202), .A2(n3103), .B1(n3102), .B2(n3052), .ZN(n3129)
         );
  AOI22_X1 U3859 ( .A1(n3202), .A2(n3105), .B1(n3104), .B2(n3052), .ZN(n3192)
         );
  MUX2_X1 U3860 ( .A(n3129), .B(n3192), .S(n2101), .Z(n3117) );
  OAI21_X1 U3861 ( .B1(n3055), .B2(n3117), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N99 ) );
  MUX2_X1 U3862 ( .A(n3107), .B(n3106), .S(n2101), .Z(n3149) );
  OAI21_X1 U3863 ( .B1(n3055), .B2(n3149), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N100 ) );
  MUX2_X1 U3864 ( .A(n3109), .B(n3108), .S(n2101), .Z(n3160) );
  OAI21_X1 U3865 ( .B1(n3055), .B2(n3160), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N101 ) );
  AOI22_X1 U3866 ( .A1(n2103), .A2(\DataP/alu_a_in[10] ), .B1(n2207), .B2(
        n2916), .ZN(n3152) );
  AOI22_X1 U3867 ( .A1(n3049), .A2(n3110), .B1(n3152), .B2(n3047), .ZN(n3169)
         );
  AOI22_X1 U3868 ( .A1(n3202), .A2(n3111), .B1(n3169), .B2(n2919), .ZN(n3191)
         );
  AOI22_X1 U3869 ( .A1(n2103), .A2(\DataP/alu_a_in[8] ), .B1(
        \DataP/alu_a_in[7] ), .B2(n3199), .ZN(n3151) );
  AOI22_X1 U3870 ( .A1(n2103), .A2(\DataP/alu_a_in[6] ), .B1(
        \DataP/alu_a_in[5] ), .B2(n3199), .ZN(n3154) );
  AOI22_X1 U3871 ( .A1(n3049), .A2(n3151), .B1(n3154), .B2(n3047), .ZN(n3168)
         );
  AOI22_X1 U3872 ( .A1(n2103), .A2(\DataP/alu_a_in[4] ), .B1(n1973), .B2(n3199), .ZN(n3153) );
  AOI22_X1 U3873 ( .A1(n2103), .A2(\DataP/alu_a_in[2] ), .B1(n2232), .B2(n3199), .ZN(n3112) );
  AOI22_X1 U3874 ( .A1(n3048), .A2(n3153), .B1(n3112), .B2(n3201), .ZN(n3113)
         );
  AOI22_X1 U3875 ( .A1(n3202), .A2(n3168), .B1(n3113), .B2(n3052), .ZN(n3114)
         );
  AOI22_X1 U3876 ( .A1(n3205), .A2(n3191), .B1(n3114), .B2(n2101), .ZN(n3115)
         );
  NAND2_X1 U3877 ( .A1(n2102), .A2(n3115), .ZN(n3116) );
  OAI21_X1 U3878 ( .B1(n2102), .B2(n3117), .A(n3116), .ZN(
        \DataP/ALU_C/shifter/N83 ) );
  MUX2_X1 U3879 ( .A(n3119), .B(n3118), .S(n2101), .Z(n3167) );
  OAI21_X1 U3880 ( .B1(n3055), .B2(n3167), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N102 ) );
  MUX2_X1 U3881 ( .A(n3121), .B(n3120), .S(n2101), .Z(n3174) );
  OAI21_X1 U3882 ( .B1(n3055), .B2(n3174), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N103 ) );
  MUX2_X1 U3883 ( .A(n3123), .B(n3122), .S(n2101), .Z(n3181) );
  OAI21_X1 U3884 ( .B1(n2138), .B2(n3181), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N104 ) );
  OAI21_X1 U3885 ( .B1(n3205), .B2(n3124), .A(n3128), .ZN(n3125) );
  OAI21_X1 U3886 ( .B1(n3055), .B2(n3196), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N105 ) );
  OAI21_X1 U3887 ( .B1(n3205), .B2(n3126), .A(n3128), .ZN(n3127) );
  OAI21_X1 U3888 ( .B1(n3055), .B2(n3197), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N106 ) );
  OAI21_X1 U3889 ( .B1(n3205), .B2(n3129), .A(n3128), .ZN(n3130) );
  OAI21_X1 U3890 ( .B1(n2138), .B2(n3198), .A(n3131), .ZN(
        \DataP/ALU_C/shifter/N107 ) );
  AOI21_X1 U3891 ( .B1(n3206), .B2(n3132), .A(n3195), .ZN(n3133) );
  AOI21_X1 U3892 ( .B1(n2102), .B2(n3134), .A(n3195), .ZN(n3135) );
  AOI21_X1 U3893 ( .B1(n3206), .B2(n3136), .A(n3195), .ZN(n3137) );
  AOI21_X1 U3894 ( .B1(n2102), .B2(n3138), .A(n3195), .ZN(n3139) );
  AOI22_X1 U3895 ( .A1(n3048), .A2(n3141), .B1(n3140), .B2(n3047), .ZN(n3175)
         );
  AOI22_X1 U3896 ( .A1(n3050), .A2(n3143), .B1(n3142), .B2(n3047), .ZN(n3144)
         );
  AOI22_X1 U3897 ( .A1(n3202), .A2(n3175), .B1(n3144), .B2(n2919), .ZN(n3145)
         );
  AOI22_X1 U3898 ( .A1(n3205), .A2(n3146), .B1(n3145), .B2(n2101), .ZN(n3147)
         );
  NAND2_X1 U3899 ( .A1(n2102), .A2(n3147), .ZN(n3148) );
  OAI21_X1 U3900 ( .B1(n3206), .B2(n3149), .A(n3148), .ZN(
        \DataP/ALU_C/shifter/N84 ) );
  AOI22_X1 U3901 ( .A1(n3048), .A2(n3152), .B1(n3151), .B2(n3047), .ZN(n3182)
         );
  AOI22_X1 U3902 ( .A1(n3049), .A2(n3154), .B1(n3153), .B2(n3047), .ZN(n3155)
         );
  AOI22_X1 U3903 ( .A1(n3202), .A2(n3182), .B1(n3155), .B2(n3052), .ZN(n3156)
         );
  AOI22_X1 U3904 ( .A1(n3205), .A2(n3157), .B1(n3156), .B2(n2101), .ZN(n3158)
         );
  NAND2_X1 U3905 ( .A1(n2102), .A2(n3158), .ZN(n3159) );
  AOI22_X1 U3906 ( .A1(n3202), .A2(n3162), .B1(n3161), .B2(n2919), .ZN(n3163)
         );
  AOI22_X1 U3907 ( .A1(n3205), .A2(n3164), .B1(n3163), .B2(n2101), .ZN(n3165)
         );
  NAND2_X1 U3908 ( .A1(n2102), .A2(n3165), .ZN(n3166) );
  AOI22_X1 U3909 ( .A1(n3202), .A2(n3169), .B1(n3168), .B2(n2918), .ZN(n3170)
         );
  AOI22_X1 U3910 ( .A1(n3205), .A2(n3171), .B1(n3170), .B2(n2101), .ZN(n3172)
         );
  NAND2_X1 U3911 ( .A1(n2102), .A2(n3172), .ZN(n3173) );
  AOI22_X1 U3912 ( .A1(n3202), .A2(n3176), .B1(n3175), .B2(n3052), .ZN(n3177)
         );
  AOI22_X1 U3913 ( .A1(n3205), .A2(n3178), .B1(n3177), .B2(n2101), .ZN(n3179)
         );
  NAND2_X1 U3914 ( .A1(n2102), .A2(n3179), .ZN(n3180) );
  AOI22_X1 U3915 ( .A1(n3203), .A2(n3183), .B1(n3182), .B2(n2918), .ZN(n3184)
         );
  AOI22_X1 U3916 ( .A1(n3204), .A2(n3185), .B1(n3184), .B2(n2101), .ZN(n3186)
         );
  NAND2_X1 U3917 ( .A1(n2102), .A2(n3186), .ZN(n3187) );
  AOI22_X1 U3918 ( .A1(n3205), .A2(n3192), .B1(n3191), .B2(n2101), .ZN(n3193)
         );
  NAND2_X1 U3919 ( .A1(n3206), .A2(n3193), .ZN(n3194) );
  INV_X1 U3920 ( .A(n3054), .ZN(n3204) );
  INV_X1 U3921 ( .A(n2072), .ZN(n3209) );
  MUX2_X1 U3922 ( .A(n3247), .B(\DataP/opcode_M[2] ), .S(\DataP/opcode_M[4] ), 
        .Z(n3248) );
  XOR2_X1 U3923 ( .A(n1625), .B(n524), .Z(n3267) );
  XOR2_X1 U3924 ( .A(n1621), .B(n523), .Z(n3266) );
  NAND3_X1 U3925 ( .A1(n3268), .A2(n3267), .A3(n3266), .ZN(n3271) );
  MUX2_X1 U3926 ( .A(\DataP/opcode_E[0] ), .B(\DataP/opcode_E[3] ), .S(
        \DataP/opcode_E[1] ), .Z(n3280) );
  MUX2_X1 U3927 ( .A(n3282), .B(n3281), .S(\DataP/opcode_E[4] ), .Z(n3287) );
  NAND3_X1 U3928 ( .A1(n3407), .A2(n443), .A3(ALU_OPCODE_i[3]), .ZN(n3408) );
  NAND3_X1 U3929 ( .A1(ALU_OPCODE_i[0]), .A2(ALU_OPCODE_i[3]), .A3(n3431), 
        .ZN(n3892) );
  MUX2_X1 U3930 ( .A(n3459), .B(n3448), .S(n2108), .Z(n3447) );
  NAND3_X1 U3931 ( .A1(n2200), .A2(n3886), .A3(n2151), .ZN(n3490) );
  NAND3_X1 U3932 ( .A1(n3563), .A2(ALU_OPCODE_i[3]), .A3(n2395), .ZN(n3570) );
  XOR2_X1 U3933 ( .A(n1741), .B(n3576), .Z(n3582) );
  XOR2_X1 U3934 ( .A(n1740), .B(n3587), .Z(n3594) );
  NAND3_X1 U3935 ( .A1(\DataP/alu_a_in[15] ), .A2(n3886), .A3(
        \DataP/alu_b_in[15] ), .ZN(n3637) );
  NAND3_X1 U3936 ( .A1(n3639), .A2(n2371), .A3(n2230), .ZN(n3640) );
  NAND3_X1 U3937 ( .A1(n3656), .A2(n3655), .A3(n3654), .ZN(n3657) );
  MUX2_X1 U3938 ( .A(n3670), .B(n2122), .S(n3886), .Z(n3671) );
  NAND3_X1 U3939 ( .A1(n3692), .A2(n2122), .A3(n2124), .ZN(n3693) );
  MUX2_X1 U3940 ( .A(n2120), .B(n3723), .S(n2108), .Z(n3816) );
  XOR2_X1 U3941 ( .A(n3729), .B(n1596), .Z(n3737) );
  NAND3_X1 U3942 ( .A1(n3735), .A2(n3734), .A3(n3733), .ZN(n3736) );
  NAND3_X1 U3943 ( .A1(n3745), .A2(n3744), .A3(n3743), .ZN(n3746) );
  XOR2_X1 U3944 ( .A(n3767), .B(n3753), .Z(n3761) );
  NAND3_X1 U3945 ( .A1(n3759), .A2(n3758), .A3(n3757), .ZN(n3760) );
  NAND3_X1 U3946 ( .A1(n3794), .A2(n3793), .A3(n3792), .ZN(n3795) );
  NAND3_X1 U3947 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3805) );
  NAND3_X1 U3948 ( .A1(n3814), .A2(n3813), .A3(n3812), .ZN(n3815) );
  MUX2_X1 U3949 ( .A(n3839), .B(n3856), .S(\DataP/alu_a_in[8] ), .Z(n3842) );
  NAND3_X1 U3950 ( .A1(\DataP/alu_a_in[13] ), .A2(n3890), .A3(n2141), .ZN(
        n3870) );
  MUX2_X1 U3951 ( .A(n3887), .B(n3898), .S(n3886), .Z(n3889) );
  NAND3_X1 U3952 ( .A1(n3893), .A2(n3892), .A3(n3891), .ZN(n3895) );
  AOI22_X1 U3953 ( .A1(n2132), .A2(\DataP/npc_pre[30] ), .B1(
        \DataP/pc_out[30] ), .B2(n3233), .ZN(n3968) );
  AOI22_X1 U3954 ( .A1(n2132), .A2(\DataP/npc_pre[28] ), .B1(
        \DataP/pc_out[28] ), .B2(n3233), .ZN(n3952) );
  AOI22_X1 U3955 ( .A1(n2132), .A2(\DataP/npc_pre[26] ), .B1(
        \DataP/pc_out[26] ), .B2(n3233), .ZN(n3953) );
  AOI22_X1 U3956 ( .A1(n2132), .A2(\DataP/npc_pre[24] ), .B1(
        \DataP/pc_out[24] ), .B2(n3233), .ZN(n3963) );
  AOI22_X1 U3957 ( .A1(n2132), .A2(\DataP/npc_pre[22] ), .B1(
        \DataP/pc_out[22] ), .B2(n3233), .ZN(n3962) );
  AOI22_X1 U3958 ( .A1(n2132), .A2(\DataP/npc_pre[20] ), .B1(
        \DataP/pc_out[20] ), .B2(n3233), .ZN(n3959) );
  AOI22_X1 U3959 ( .A1(n2132), .A2(\DataP/npc_pre[18] ), .B1(
        \DataP/pc_out[18] ), .B2(n3233), .ZN(n3964) );
  AOI22_X1 U3960 ( .A1(n2132), .A2(\DataP/npc_pre[16] ), .B1(
        \DataP/pc_out[16] ), .B2(n3233), .ZN(n3958) );
  AOI22_X1 U3961 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[14] ), .B1(
        \DataP/pc_out[14] ), .B2(n3233), .ZN(n3957) );
  AOI22_X1 U3962 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[12] ), .B1(
        \DataP/pc_out[12] ), .B2(n3233), .ZN(n3965) );
  AOI22_X1 U3963 ( .A1(n2132), .A2(\DataP/npc_pre[10] ), .B1(
        \DataP/pc_out[10] ), .B2(n3233), .ZN(n3973) );
  AOI22_X1 U3964 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[8] ), .B1(
        IRAM_ADDRESS[6]), .B2(n3233), .ZN(n3935) );
  AOI22_X1 U3965 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[6] ), .B1(
        IRAM_ADDRESS[4]), .B2(n3233), .ZN(n3941) );
  AOI22_X1 U3966 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[4] ), .B1(
        IRAM_ADDRESS[2]), .B2(n3233), .ZN(n3948) );
  AOI22_X1 U3967 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[2] ), .B1(
        IRAM_ADDRESS[0]), .B2(n3233), .ZN(\DataP/NPC_add/N3 ) );
  AOI22_X1 U3968 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[3] ), .B1(
        IRAM_ADDRESS[1]), .B2(n3233), .ZN(n3950) );
  NOR2_X1 U3969 ( .A1(\DataP/NPC_add/N3 ), .A2(n3950), .ZN(n3949) );
  INV_X1 U3970 ( .A(n3949), .ZN(n3947) );
  NOR2_X1 U3971 ( .A1(n3948), .A2(n3947), .ZN(n3946) );
  OAI221_X1 U3972 ( .B1(n2132), .B2(IRAM_ADDRESS[3]), .C1(n3233), .C2(
        \DataP/npc_pre[5] ), .A(n3946), .ZN(n3942) );
  NOR2_X1 U3973 ( .A1(n3941), .A2(n3942), .ZN(n3940) );
  OAI221_X1 U3974 ( .B1(n2132), .B2(IRAM_ADDRESS[5]), .C1(n3233), .C2(
        \DataP/npc_pre[7] ), .A(n3940), .ZN(n3936) );
  NOR2_X1 U3975 ( .A1(n3935), .A2(n3936), .ZN(n3934) );
  OAI221_X1 U3976 ( .B1(n2132), .B2(IRAM_ADDRESS[7]), .C1(n3233), .C2(
        \DataP/npc_pre[9] ), .A(n3934), .ZN(n3972) );
  NOR2_X1 U3977 ( .A1(n3973), .A2(n3972), .ZN(n3930) );
  MUX2_X1 U3978 ( .A(\DataP/pc_out[11] ), .B(\DataP/npc_pre[11] ), .S(n2132), 
        .Z(n3969) );
  NAND2_X1 U3979 ( .A1(n3930), .A2(n3969), .ZN(n3929) );
  NOR2_X1 U3980 ( .A1(n3965), .A2(n3929), .ZN(n3928) );
  MUX2_X1 U3981 ( .A(\DataP/pc_out[13] ), .B(\DataP/npc_pre[13] ), .S(n2132), 
        .Z(n3960) );
  NAND2_X1 U3982 ( .A1(n3928), .A2(n3960), .ZN(n3927) );
  NOR2_X1 U3983 ( .A1(n3957), .A2(n3927), .ZN(n3926) );
  MUX2_X1 U3984 ( .A(\DataP/pc_out[15] ), .B(\DataP/npc_pre[15] ), .S(n2132), 
        .Z(n3956) );
  NAND2_X1 U3985 ( .A1(n3926), .A2(n3956), .ZN(n3925) );
  NOR2_X1 U3986 ( .A1(n3958), .A2(n3925), .ZN(n3924) );
  MUX2_X1 U3987 ( .A(\DataP/pc_out[17] ), .B(\DataP/npc_pre[17] ), .S(n2132), 
        .Z(n3966) );
  NAND2_X1 U3988 ( .A1(n3924), .A2(n3966), .ZN(n3923) );
  NOR2_X1 U3989 ( .A1(n3964), .A2(n3923), .ZN(n3922) );
  MUX2_X1 U3990 ( .A(\DataP/pc_out[19] ), .B(\DataP/npc_pre[19] ), .S(n2132), 
        .Z(n3961) );
  NAND2_X1 U3991 ( .A1(n3922), .A2(n3961), .ZN(n3921) );
  NOR2_X1 U3992 ( .A1(n3959), .A2(n3921), .ZN(n3920) );
  MUX2_X1 U3993 ( .A(\DataP/pc_out[21] ), .B(\DataP/npc_pre[21] ), .S(n2132), 
        .Z(n3970) );
  NAND2_X1 U3994 ( .A1(n3920), .A2(n3970), .ZN(n3919) );
  NOR2_X1 U3995 ( .A1(n3962), .A2(n3919), .ZN(n3918) );
  MUX2_X1 U3996 ( .A(\DataP/pc_out[23] ), .B(\DataP/npc_pre[23] ), .S(n2132), 
        .Z(n3971) );
  NAND2_X1 U3997 ( .A1(n3918), .A2(n3971), .ZN(n3917) );
  NOR2_X1 U3998 ( .A1(n3963), .A2(n3917), .ZN(n3916) );
  MUX2_X1 U3999 ( .A(\DataP/pc_out[25] ), .B(\DataP/npc_pre[25] ), .S(n2132), 
        .Z(n3954) );
  NAND2_X1 U4000 ( .A1(n3916), .A2(n3954), .ZN(n3915) );
  NOR2_X1 U4001 ( .A1(n3953), .A2(n3915), .ZN(n3914) );
  MUX2_X1 U4002 ( .A(\DataP/pc_out[27] ), .B(\DataP/npc_pre[27] ), .S(n2132), 
        .Z(n3955) );
  NAND2_X1 U4003 ( .A1(n3914), .A2(n3955), .ZN(n3913) );
  NOR2_X1 U4004 ( .A1(n3952), .A2(n3913), .ZN(n3912) );
  MUX2_X1 U4005 ( .A(\DataP/pc_out[29] ), .B(\DataP/npc_pre[29] ), .S(n2132), 
        .Z(n3967) );
  NAND2_X1 U4006 ( .A1(n3912), .A2(n3967), .ZN(n3911) );
  NOR2_X1 U4007 ( .A1(n3968), .A2(n3911), .ZN(n3951) );
  AOI21_X1 U4008 ( .B1(n3968), .B2(n3911), .A(n3951), .ZN(\DataP/NPC_add/N31 )
         );
  XOR2_X1 U4009 ( .A(n3912), .B(n3967), .Z(\DataP/NPC_add/N30 ) );
  AOI21_X1 U4010 ( .B1(n3952), .B2(n3913), .A(n3912), .ZN(\DataP/NPC_add/N29 )
         );
  XOR2_X1 U4011 ( .A(n3914), .B(n3955), .Z(\DataP/NPC_add/N28 ) );
  AOI21_X1 U4012 ( .B1(n3953), .B2(n3915), .A(n3914), .ZN(\DataP/NPC_add/N27 )
         );
  XOR2_X1 U4013 ( .A(n3916), .B(n3954), .Z(\DataP/NPC_add/N26 ) );
  AOI21_X1 U4014 ( .B1(n3963), .B2(n3917), .A(n3916), .ZN(\DataP/NPC_add/N25 )
         );
  XOR2_X1 U4015 ( .A(n3918), .B(n3971), .Z(\DataP/NPC_add/N24 ) );
  AOI21_X1 U4016 ( .B1(n3962), .B2(n3919), .A(n3918), .ZN(\DataP/NPC_add/N23 )
         );
  XOR2_X1 U4017 ( .A(n3920), .B(n3970), .Z(\DataP/NPC_add/N22 ) );
  AOI21_X1 U4018 ( .B1(n3959), .B2(n3921), .A(n3920), .ZN(\DataP/NPC_add/N21 )
         );
  XOR2_X1 U4019 ( .A(n3922), .B(n3961), .Z(\DataP/NPC_add/N20 ) );
  AOI21_X1 U4020 ( .B1(n3964), .B2(n3923), .A(n3922), .ZN(\DataP/NPC_add/N19 )
         );
  XOR2_X1 U4021 ( .A(n3924), .B(n3966), .Z(\DataP/NPC_add/N18 ) );
  AOI21_X1 U4022 ( .B1(n3958), .B2(n3925), .A(n3924), .ZN(\DataP/NPC_add/N17 )
         );
  XOR2_X1 U4023 ( .A(n3926), .B(n3956), .Z(\DataP/NPC_add/N16 ) );
  AOI21_X1 U4024 ( .B1(n3957), .B2(n3927), .A(n3926), .ZN(\DataP/NPC_add/N15 )
         );
  XOR2_X1 U4025 ( .A(n3928), .B(n3960), .Z(\DataP/NPC_add/N14 ) );
  AOI21_X1 U4026 ( .B1(n3965), .B2(n3929), .A(n3928), .ZN(\DataP/NPC_add/N13 )
         );
  XOR2_X1 U4027 ( .A(n3930), .B(n3969), .Z(\DataP/NPC_add/N12 ) );
  AOI21_X1 U4028 ( .B1(n3973), .B2(n3972), .A(n3930), .ZN(\DataP/NPC_add/N11 )
         );
  AOI22_X1 U4029 ( .A1(n2132), .A2(\DataP/npc_pre[9] ), .B1(IRAM_ADDRESS[7]), 
        .B2(n3233), .ZN(n3933) );
  INV_X1 U4030 ( .A(n3934), .ZN(n3932) );
  INV_X1 U4031 ( .A(n3972), .ZN(n3931) );
  AOI21_X1 U4032 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(\DataP/NPC_add/N10 )
         );
  AOI21_X1 U4033 ( .B1(n3935), .B2(n3936), .A(n3934), .ZN(\DataP/NPC_add/N9 )
         );
  AOI22_X1 U4034 ( .A1(n2132), .A2(\DataP/npc_pre[7] ), .B1(IRAM_ADDRESS[5]), 
        .B2(n3233), .ZN(n3939) );
  INV_X1 U4035 ( .A(n3940), .ZN(n3938) );
  INV_X1 U4036 ( .A(n3936), .ZN(n3937) );
  AOI21_X1 U4037 ( .B1(n3939), .B2(n3938), .A(n3937), .ZN(\DataP/NPC_add/N8 )
         );
  AOI21_X1 U4038 ( .B1(n3941), .B2(n3942), .A(n3940), .ZN(\DataP/NPC_add/N7 )
         );
  AOI22_X1 U4039 ( .A1(n2132), .A2(\DataP/npc_pre[5] ), .B1(IRAM_ADDRESS[3]), 
        .B2(n3233), .ZN(n3945) );
  INV_X1 U4040 ( .A(n3946), .ZN(n3944) );
  INV_X1 U4041 ( .A(n3942), .ZN(n3943) );
  AOI21_X1 U4042 ( .B1(n3945), .B2(n3944), .A(n3943), .ZN(\DataP/NPC_add/N6 )
         );
  AOI21_X1 U4043 ( .B1(n3948), .B2(n3947), .A(n3946), .ZN(\DataP/NPC_add/N5 )
         );
  AOI21_X1 U4044 ( .B1(n3950), .B2(\DataP/NPC_add/N3 ), .A(n3949), .ZN(
        \DataP/NPC_add/N4 ) );
  AOI22_X1 U4045 ( .A1(n2132), .A2(\DataP/npc_pre[31] ), .B1(
        \DataP/pc_out[31] ), .B2(n3233), .ZN(n3974) );
  XNOR2_X1 U4046 ( .A(n3974), .B(n3951), .ZN(\DataP/NPC_add/N32 ) );
  NAND2_X1 U4049 ( .A1(n514), .A2(n515), .ZN(n4155) );
  NAND2_X1 U4050 ( .A1(IR_CU_28), .A2(n516), .ZN(n3980) );
  NOR2_X1 U4051 ( .A1(n4155), .A2(n3980), .ZN(n607) );
  NAND2_X1 U4052 ( .A1(IR_CU_27), .A2(n497), .ZN(n4151) );
  NOR2_X1 U4053 ( .A1(n514), .A2(n515), .ZN(n4176) );
  NAND3_X1 U4054 ( .A1(IR_CU_31), .A2(n4176), .A3(n1960), .ZN(n4012) );
  NOR2_X1 U4055 ( .A1(IR_CU_27), .A2(n497), .ZN(n3996) );
  INV_X1 U4056 ( .A(n4176), .ZN(n4177) );
  NOR2_X1 U4057 ( .A1(n3980), .A2(n4177), .ZN(n4013) );
  NOR3_X1 U4058 ( .A1(IR_CU_27), .A2(n4155), .A3(n516), .ZN(n4046) );
  AOI22_X1 U4059 ( .A1(IR_CU_31), .A2(n4166), .B1(n2374), .B2(n504), .ZN(n3975) );
  NAND2_X1 U4060 ( .A1(n515), .A2(n1960), .ZN(n4044) );
  NOR3_X1 U4061 ( .A1(n514), .A2(n2377), .A3(n3980), .ZN(n3995) );
  AOI22_X1 U4062 ( .A1(n4055), .A2(n607), .B1(n4052), .B2(n3995), .ZN(n3997)
         );
  NAND3_X1 U4063 ( .A1(n4166), .A2(n16), .A3(n2377), .ZN(n4156) );
  OAI211_X1 U4064 ( .C1(n3975), .C2(n4044), .A(n3997), .B(n4156), .ZN(n3976)
         );
  AOI211_X1 U4065 ( .C1(n3996), .C2(n4013), .A(n4046), .B(n3976), .ZN(n3987)
         );
  NOR4_X1 U4066 ( .A1(IR_CU[8]), .A2(IR_CU[6]), .A3(IR_CU[7]), .A4(IR_CU[9]), 
        .ZN(n3977) );
  NAND3_X1 U4067 ( .A1(n4153), .A2(n484), .A3(n3977), .ZN(n3989) );
  NOR2_X1 U4068 ( .A1(n479), .A2(n3989), .ZN(n4023) );
  NAND2_X1 U4069 ( .A1(IR_CU[5]), .A2(n4023), .ZN(n4001) );
  NOR3_X1 U4070 ( .A1(n477), .A2(n2375), .A3(n4001), .ZN(n3985) );
  NOR3_X1 U4071 ( .A1(n478), .A2(n3989), .A3(n2399), .ZN(n4003) );
  NAND2_X1 U4072 ( .A1(n4003), .A2(n476), .ZN(n4005) );
  OAI21_X1 U4073 ( .B1(n476), .B2(n479), .A(n2375), .ZN(n3978) );
  OAI211_X1 U4074 ( .C1(n479), .C2(n2375), .A(n3978), .B(n477), .ZN(n3979) );
  NAND2_X1 U4075 ( .A1(IR_CU[5]), .A2(n480), .ZN(n4035) );
  AOI221_X1 U4076 ( .B1(n3989), .B2(n4005), .C1(n3979), .C2(n4005), .A(n4035), 
        .ZN(n3984) );
  INV_X1 U4077 ( .A(n3985), .ZN(n4032) );
  NOR3_X1 U4078 ( .A1(n3994), .A2(n4155), .A3(n4151), .ZN(n4020) );
  INV_X1 U4079 ( .A(n3980), .ZN(n3981) );
  NAND3_X1 U4080 ( .A1(n514), .A2(n3981), .A3(n2377), .ZN(n4016) );
  NAND4_X1 U4081 ( .A1(n4003), .A2(IR_CU[1]), .A3(n480), .A4(n482), .ZN(n4026)
         );
  OAI21_X1 U4082 ( .B1(n504), .B2(n4016), .A(n4026), .ZN(n4000) );
  AOI211_X1 U4083 ( .C1(n4055), .C2(n3995), .A(n4020), .B(n4000), .ZN(n3983)
         );
  NAND3_X1 U4084 ( .A1(n4166), .A2(n4176), .A3(n1960), .ZN(n3982) );
  OAI211_X1 U4085 ( .C1(n4032), .C2(n476), .A(n3983), .B(n3982), .ZN(n3991) );
  AOI211_X1 U4086 ( .C1(n3985), .C2(IR_CU[4]), .A(n3984), .B(n3991), .ZN(n3986) );
  OAI211_X1 U4087 ( .C1(n4151), .C2(n4012), .A(n3987), .B(n3986), .ZN(
        \CU_I/aluOpcode_i[0] ) );
  INV_X1 U4088 ( .A(n3994), .ZN(n4168) );
  NAND2_X1 U4089 ( .A1(n4168), .A2(IR_CU_27), .ZN(n4154) );
  NOR2_X1 U4090 ( .A1(IR_CU[1]), .A2(n478), .ZN(n3988) );
  AOI22_X1 U4091 ( .A1(IR_CU[1]), .A2(n478), .B1(n3988), .B2(n476), .ZN(n4002)
         );
  NOR3_X1 U4092 ( .A1(n4002), .A2(n4035), .A3(n3989), .ZN(n3990) );
  AOI21_X1 U4093 ( .B1(n4013), .B2(n4055), .A(n3990), .ZN(n3993) );
  NOR3_X1 U4094 ( .A1(IR_CU[1]), .A2(n478), .A3(n4001), .ZN(n4031) );
  NOR2_X1 U4095 ( .A1(n516), .A2(n1960), .ZN(n4174) );
  NAND2_X1 U4096 ( .A1(n4176), .A2(n4174), .ZN(n4027) );
  AOI211_X1 U4097 ( .C1(n4031), .C2(n476), .A(n3991), .B(n4006), .ZN(n3992) );
  OAI211_X1 U4098 ( .C1(n514), .C2(n4154), .A(n3993), .B(n3992), .ZN(
        \CU_I/aluOpcode_i[1] ) );
  INV_X1 U4099 ( .A(n4166), .ZN(n4048) );
  NOR3_X1 U4100 ( .A1(n3994), .A2(n4155), .A3(n4048), .ZN(n4019) );
  NOR3_X1 U4101 ( .A1(n3994), .A2(n4036), .A3(n4177), .ZN(n4030) );
  INV_X1 U4102 ( .A(n3995), .ZN(n3998) );
  INV_X1 U4103 ( .A(n3996), .ZN(n4170) );
  OAI21_X1 U4104 ( .B1(n3998), .B2(n4170), .A(n3997), .ZN(n3999) );
  NOR4_X1 U4105 ( .A1(n4019), .A2(n4030), .A3(n4000), .A4(n3999), .ZN(n4011)
         );
  NOR3_X1 U4106 ( .A1(n4002), .A2(n4001), .A3(n480), .ZN(n4009) );
  NAND3_X1 U4107 ( .A1(n478), .A2(n4023), .A3(n476), .ZN(n4034) );
  NAND2_X1 U4108 ( .A1(n4003), .A2(IR_CU[0]), .ZN(n4004) );
  AOI211_X1 U4109 ( .C1(n4034), .C2(n4004), .A(IR_CU[1]), .B(n4035), .ZN(n4008) );
  NOR3_X1 U4110 ( .A1(IR_CU[4]), .A2(n477), .A3(n4005), .ZN(n4007) );
  NOR4_X1 U4111 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  OAI211_X1 U4112 ( .C1(n504), .C2(n4012), .A(n4011), .B(n4010), .ZN(
        \CU_I/aluOpcode_i[2] ) );
  AOI211_X1 U4113 ( .C1(IR_CU_31), .C2(n1960), .A(n4177), .B(n4170), .ZN(n4018) );
  NAND2_X1 U4114 ( .A1(n4055), .A2(n4013), .ZN(n4015) );
  NAND2_X1 U4115 ( .A1(n607), .A2(n504), .ZN(n4014) );
  OAI211_X1 U4116 ( .C1(n4048), .C2(n4016), .A(n4015), .B(n4014), .ZN(n4017)
         );
  NOR4_X1 U4117 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4025)
         );
  OAI211_X1 U4118 ( .C1(n2375), .C2(n480), .A(IR_CU[5]), .B(IR_CU[0]), .ZN(
        n4021) );
  OAI21_X1 U4119 ( .B1(n478), .B2(n4035), .A(n4021), .ZN(n4022) );
  NAND3_X1 U4120 ( .A1(n4023), .A2(n477), .A3(n4022), .ZN(n4024) );
  OAI211_X1 U4121 ( .C1(n476), .C2(n4026), .A(n4025), .B(n4024), .ZN(
        \CU_I/aluOpcode_i[3] ) );
  OAI211_X1 U4122 ( .C1(n516), .C2(n2374), .A(n1960), .B(n2377), .ZN(n4028) );
  AOI22_X1 U4123 ( .A1(IR_CU_27), .A2(n4028), .B1(n4027), .B2(n504), .ZN(n4029) );
  AOI211_X1 U4124 ( .C1(n4031), .C2(IR_CU[4]), .A(n4030), .B(n4029), .ZN(n4033) );
  OAI211_X1 U4125 ( .C1(n4035), .C2(n4034), .A(n4033), .B(n4032), .ZN(
        \CU_I/aluOpcode_i[4] ) );
  OAI211_X1 U4126 ( .C1(IR_CU_26), .C2(n2377), .A(IR_CU_28), .B(IR_CU_27), 
        .ZN(n4038) );
  NOR3_X1 U4127 ( .A1(n515), .A2(n1960), .A3(n4036), .ZN(n4037) );
  AOI21_X1 U4128 ( .B1(n2374), .B2(n4038), .A(n4037), .ZN(n4056) );
  NOR3_X1 U4129 ( .A1(n515), .A2(n2374), .A3(n504), .ZN(n4058) );
  INV_X1 U4130 ( .A(n4044), .ZN(n4039) );
  AOI22_X1 U4131 ( .A1(IR_CU_28), .A2(n4058), .B1(n4055), .B2(n4039), .ZN(
        n4040) );
  AOI22_X1 U4132 ( .A1(IR_CU_28), .A2(IR_CU_27), .B1(n504), .B2(n1960), .ZN(
        n4043) );
  NAND2_X1 U4133 ( .A1(n4176), .A2(n4043), .ZN(n4059) );
  OAI221_X1 U4134 ( .B1(IR_CU_31), .B2(n4056), .C1(IR_CU_31), .C2(n4040), .A(
        n4059), .ZN(n4045) );
  AOI21_X1 U4135 ( .B1(n4168), .B2(n4166), .A(n4045), .ZN(n1372) );
  AOI21_X1 U4136 ( .B1(IR_CU_26), .B2(n1960), .A(n504), .ZN(n4042) );
  INV_X1 U4137 ( .A(n4155), .ZN(n4173) );
  NAND2_X1 U4138 ( .A1(IR_CU_31), .A2(n4173), .ZN(n4041) );
  OAI21_X1 U4139 ( .B1(n4042), .B2(n4041), .A(n1372), .ZN(\CU_I/cw[0] ) );
  AND3_X1 U4140 ( .A1(n4173), .A2(n4043), .A3(n516), .ZN(\CU_I/cw[10] ) );
  AOI21_X1 U4141 ( .B1(n4151), .B2(n4049), .A(n4046), .ZN(n4061) );
  INV_X1 U4142 ( .A(n4061), .ZN(\CU_I/cw[6] ) );
  OR2_X1 U4143 ( .A1(n4045), .A2(\CU_I/cw[6] ), .ZN(\CU_I/cw[1] ) );
  NAND2_X1 U4144 ( .A1(n4049), .A2(n2374), .ZN(n4051) );
  AOI22_X1 U4145 ( .A1(n4049), .A2(n4055), .B1(n4046), .B2(n1960), .ZN(n4047)
         );
  OAI21_X1 U4146 ( .B1(n4048), .B2(n4051), .A(n4047), .ZN(\CU_I/cw[3] ) );
  NAND2_X1 U4147 ( .A1(n4173), .A2(n4174), .ZN(n4053) );
  OAI211_X1 U4148 ( .C1(n2374), .C2(n497), .A(n4049), .B(n504), .ZN(n4050) );
  OAI21_X1 U4149 ( .B1(n4170), .B2(n4053), .A(n4050), .ZN(\CU_I/cw[4] ) );
  INV_X1 U4150 ( .A(n4053), .ZN(n4054) );
  AOI21_X1 U4151 ( .B1(n4055), .B2(n4054), .A(\CU_I/cw[7] ), .ZN(n1358) );
  INV_X1 U4152 ( .A(n4056), .ZN(n4057) );
  AOI221_X1 U4153 ( .B1(n4058), .B2(n516), .C1(n4057), .C2(n516), .A(
        \CU_I/cw[10] ), .ZN(n4060) );
  NAND3_X1 U4154 ( .A1(n443), .A2(ALU_OPCODE_i[2]), .A3(ALU_OPCODE_i[1]), .ZN(
        n4101) );
  NOR4_X1 U4155 ( .A1(\DataP/alu_out_W[12] ), .A2(\DataP/alu_out_W[11] ), .A3(
        \DataP/alu_out_W[10] ), .A4(\DataP/alu_out_W[0] ), .ZN(n4065) );
  NOR4_X1 U4156 ( .A1(\DataP/alu_out_W[15] ), .A2(\DataP/alu_out_W[14] ), .A3(
        \DataP/alu_out_W[13] ), .A4(\DataP/alu_out_W[16] ), .ZN(n4064) );
  NOR4_X1 U4157 ( .A1(\DataP/alu_out_W[17] ), .A2(\DataP/alu_out_W[19] ), .A3(
        \DataP/alu_out_W[18] ), .A4(\DataP/alu_out_W[1] ), .ZN(n4063) );
  NOR4_X1 U4158 ( .A1(\DataP/alu_out_W[23] ), .A2(\DataP/alu_out_W[21] ), .A3(
        \DataP/alu_out_W[20] ), .A4(\DataP/alu_out_W[22] ), .ZN(n4062) );
  NAND4_X1 U4159 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4098)
         );
  INV_X1 U4160 ( .A(\DataP/FWD_MUX_BR_S[0] ), .ZN(n4070) );
  NAND2_X1 U4161 ( .A1(n4070), .A2(\DataP/FWD_MUX_BR_S[1] ), .ZN(n4079) );
  INV_X1 U4162 ( .A(n4079), .ZN(n4097) );
  NOR4_X1 U4163 ( .A1(\DataP/alu_out_W[27] ), .A2(\DataP/alu_out_W[26] ), .A3(
        \DataP/alu_out_W[25] ), .A4(\DataP/alu_out_W[24] ), .ZN(n4069) );
  NOR4_X1 U4164 ( .A1(\DataP/alu_out_W[30] ), .A2(\DataP/alu_out_W[29] ), .A3(
        \DataP/alu_out_W[28] ), .A4(\DataP/alu_out_W[2] ), .ZN(n4068) );
  NOR4_X1 U4165 ( .A1(\DataP/alu_out_W[31] ), .A2(\DataP/alu_out_W[5] ), .A3(
        \DataP/alu_out_W[4] ), .A4(\DataP/alu_out_W[3] ), .ZN(n4067) );
  NOR4_X1 U4166 ( .A1(\DataP/alu_out_W[9] ), .A2(\DataP/alu_out_W[8] ), .A3(
        \DataP/alu_out_W[7] ), .A4(\DataP/alu_out_W[6] ), .ZN(n4066) );
  NAND4_X1 U4167 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4096)
         );
  NOR2_X1 U4168 ( .A1(\DataP/FWD_MUX_BR_S[1] ), .A2(n4070), .ZN(n4094) );
  NOR4_X1 U4169 ( .A1(\DataP/A_s[27] ), .A2(\DataP/A_s[26] ), .A3(
        \DataP/A_s[25] ), .A4(\DataP/A_s[24] ), .ZN(n4074) );
  NOR4_X1 U4170 ( .A1(\DataP/A_s[30] ), .A2(\DataP/A_s[29] ), .A3(
        \DataP/A_s[28] ), .A4(\DataP/A_s[2] ), .ZN(n4073) );
  NOR4_X1 U4171 ( .A1(\DataP/A_s[31] ), .A2(\DataP/A_s[5] ), .A3(
        \DataP/A_s[4] ), .A4(\DataP/A_s[3] ), .ZN(n4072) );
  NOR4_X1 U4172 ( .A1(\DataP/A_s[9] ), .A2(\DataP/A_s[8] ), .A3(\DataP/A_s[7] ), .A4(\DataP/A_s[6] ), .ZN(n4071) );
  NAND4_X1 U4173 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4081)
         );
  NOR4_X1 U4174 ( .A1(\DataP/A_s[12] ), .A2(\DataP/A_s[11] ), .A3(
        \DataP/A_s[10] ), .A4(\DataP/A_s[0] ), .ZN(n4078) );
  NOR4_X1 U4175 ( .A1(\DataP/A_s[15] ), .A2(\DataP/A_s[14] ), .A3(
        \DataP/A_s[13] ), .A4(\DataP/A_s[16] ), .ZN(n4077) );
  NOR4_X1 U4176 ( .A1(\DataP/A_s[17] ), .A2(\DataP/A_s[19] ), .A3(
        \DataP/A_s[18] ), .A4(\DataP/A_s[1] ), .ZN(n4076) );
  NOR4_X1 U4177 ( .A1(\DataP/A_s[23] ), .A2(\DataP/A_s[21] ), .A3(
        \DataP/A_s[20] ), .A4(\DataP/A_s[22] ), .ZN(n4075) );
  NAND4_X1 U4178 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4080)
         );
  OAI21_X1 U4179 ( .B1(n4081), .B2(n4080), .A(n4079), .ZN(n4093) );
  NOR4_X1 U4180 ( .A1(DRAM_ADDRESS[11]), .A2(DRAM_ADDRESS[10]), .A3(
        DRAM_ADDRESS[1]), .A4(DRAM_ADDRESS[0]), .ZN(n4085) );
  NOR4_X1 U4181 ( .A1(DRAM_ADDRESS[5]), .A2(DRAM_ADDRESS[4]), .A3(
        DRAM_ADDRESS[3]), .A4(DRAM_ADDRESS[2]), .ZN(n4084) );
  NOR4_X1 U4182 ( .A1(DRAM_ADDRESS[9]), .A2(DRAM_ADDRESS[8]), .A3(
        DRAM_ADDRESS[7]), .A4(DRAM_ADDRESS[6]), .ZN(n4083) );
  NOR4_X1 U4183 ( .A1(\DataP/alu_out_M[15] ), .A2(\DataP/alu_out_M[14] ), .A3(
        \DataP/alu_out_M[13] ), .A4(\DataP/alu_out_M[12] ), .ZN(n4082) );
  NAND4_X1 U4184 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4091)
         );
  NOR4_X1 U4185 ( .A1(\DataP/alu_out_M[16] ), .A2(\DataP/alu_out_M[17] ), .A3(
        \DataP/alu_out_M[19] ), .A4(\DataP/alu_out_M[18] ), .ZN(n4089) );
  NOR4_X1 U4186 ( .A1(\DataP/alu_out_M[23] ), .A2(\DataP/alu_out_M[21] ), .A3(
        \DataP/alu_out_M[20] ), .A4(\DataP/alu_out_M[22] ), .ZN(n4088) );
  NOR4_X1 U4187 ( .A1(\DataP/alu_out_M[27] ), .A2(\DataP/alu_out_M[26] ), .A3(
        \DataP/alu_out_M[25] ), .A4(\DataP/alu_out_M[24] ), .ZN(n4087) );
  NOR4_X1 U4188 ( .A1(\DataP/alu_out_M[31] ), .A2(\DataP/alu_out_M[30] ), .A3(
        \DataP/alu_out_M[29] ), .A4(\DataP/alu_out_M[28] ), .ZN(n4086) );
  NAND4_X1 U4189 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  OAI21_X1 U4190 ( .B1(n4091), .B2(n4090), .A(n4094), .ZN(n4092) );
  OAI21_X1 U4191 ( .B1(n4094), .B2(n4093), .A(n4092), .ZN(n4095) );
  AOI221_X1 U4192 ( .B1(n4098), .B2(n4097), .C1(n4096), .C2(n4097), .A(n4095), 
        .ZN(n4099) );
  XNOR2_X1 U4193 ( .A(\DataP/pr_E ), .B(n4099), .ZN(n4183) );
  NAND2_X1 U4194 ( .A1(BR_EN_i), .A2(ALU_OPCODE_i[3]), .ZN(n4182) );
  NAND2_X1 U4195 ( .A1(ALU_OPCODE_i[1]), .A2(ALU_OPCODE_i[0]), .ZN(n4100) );
  INV_X1 U4196 ( .A(\DataP/npc[8] ), .ZN(n4214) );
  INV_X1 U4197 ( .A(\DataP/npc[9] ), .ZN(n4213) );
  OAI22_X1 U4198 ( .A1(n341), .A2(n4111), .B1(n4110), .B2(n4213), .ZN(
        \DataP/PC_reg/N11 ) );
  INV_X1 U4199 ( .A(\DataP/npc[10] ), .ZN(n4212) );
  OAI22_X1 U4200 ( .A1(n340), .A2(n4111), .B1(n4110), .B2(n4212), .ZN(
        \DataP/PC_reg/N12 ) );
  INV_X1 U4201 ( .A(\DataP/npc[11] ), .ZN(n4211) );
  OAI22_X1 U4202 ( .A1(n2386), .A2(n4111), .B1(n4110), .B2(n4211), .ZN(
        \DataP/PC_reg/N13 ) );
  INV_X1 U4203 ( .A(\DataP/npc[12] ), .ZN(n4210) );
  OAI22_X1 U4204 ( .A1(n337), .A2(n4111), .B1(n4110), .B2(n4210), .ZN(
        \DataP/PC_reg/N14 ) );
  NAND3_X1 U4205 ( .A1(n2434), .A2(n4107), .A3(n4106), .ZN(n4105) );
  INV_X1 U4206 ( .A(\DataP/npc[0] ), .ZN(n4223) );
  OAI22_X1 U4207 ( .A1(n296), .A2(n4111), .B1(n4110), .B2(n4223), .ZN(
        \DataP/PC_reg/N2 ) );
  INV_X1 U4208 ( .A(\DataP/npc[1] ), .ZN(n4221) );
  OAI22_X1 U4209 ( .A1(n358), .A2(n4111), .B1(n4110), .B2(n4221), .ZN(
        \DataP/PC_reg/N3 ) );
  INV_X1 U4210 ( .A(\DataP/npc[2] ), .ZN(n4220) );
  OAI22_X1 U4211 ( .A1(n357), .A2(n4111), .B1(n4110), .B2(n4220), .ZN(
        \DataP/PC_reg/N4 ) );
  INV_X1 U4212 ( .A(\DataP/npc[3] ), .ZN(n4219) );
  INV_X1 U4213 ( .A(\DataP/npc[4] ), .ZN(n4218) );
  INV_X1 U4214 ( .A(\DataP/npc[5] ), .ZN(n4217) );
  OAI22_X1 U4215 ( .A1(n354), .A2(n4111), .B1(n4110), .B2(n4217), .ZN(
        \DataP/PC_reg/N7 ) );
  INV_X1 U4216 ( .A(\DataP/npc[6] ), .ZN(n4216) );
  INV_X1 U4217 ( .A(\DataP/npc[7] ), .ZN(n4215) );
  OAI22_X1 U4218 ( .A1(n350), .A2(n4111), .B1(n4110), .B2(n4215), .ZN(
        \DataP/PC_reg/N9 ) );
  AOI22_X1 U4219 ( .A1(n3229), .A2(\DataP/LMD_out[0] ), .B1(n4143), .B2(
        \DataP/link_addr_W[0] ), .ZN(n4112) );
  OAI21_X1 U4220 ( .B1(n2521), .B2(n4146), .A(n4112), .ZN(\DataP/WB[0] ) );
  AOI22_X1 U4221 ( .A1(n3229), .A2(\DataP/LMD_out[10] ), .B1(n4143), .B2(
        \DataP/link_addr_W[10] ), .ZN(n4113) );
  OAI21_X1 U4222 ( .B1(n2503), .B2(n4146), .A(n4113), .ZN(\DataP/WB[10] ) );
  AOI22_X1 U4223 ( .A1(n3229), .A2(\DataP/LMD_out[11] ), .B1(n4143), .B2(
        \DataP/link_addr_W[11] ), .ZN(n4114) );
  OAI21_X1 U4224 ( .B1(n2518), .B2(n4146), .A(n4114), .ZN(\DataP/WB[11] ) );
  AOI22_X1 U4225 ( .A1(n3229), .A2(\DataP/LMD_out[12] ), .B1(n4143), .B2(
        \DataP/link_addr_W[12] ), .ZN(n4115) );
  OAI21_X1 U4226 ( .B1(n2492), .B2(n4146), .A(n4115), .ZN(\DataP/WB[12] ) );
  AOI22_X1 U4227 ( .A1(n3229), .A2(\DataP/LMD_out[13] ), .B1(n4143), .B2(
        \DataP/link_addr_W[13] ), .ZN(n4116) );
  OAI21_X1 U4228 ( .B1(n2504), .B2(n4146), .A(n4116), .ZN(\DataP/WB[13] ) );
  AOI22_X1 U4229 ( .A1(n3229), .A2(\DataP/LMD_out[14] ), .B1(n4143), .B2(
        \DataP/link_addr_W[14] ), .ZN(n4117) );
  OAI21_X1 U4230 ( .B1(n2497), .B2(n4146), .A(n4117), .ZN(\DataP/WB[14] ) );
  AOI22_X1 U4231 ( .A1(n3229), .A2(\DataP/LMD_out[15] ), .B1(n4143), .B2(
        \DataP/link_addr_W[15] ), .ZN(n4118) );
  OAI21_X1 U4232 ( .B1(n2516), .B2(n4146), .A(n4118), .ZN(\DataP/WB[15] ) );
  AOI22_X1 U4233 ( .A1(n3229), .A2(\DataP/LMD_out[16] ), .B1(n4143), .B2(
        \DataP/link_addr_W[16] ), .ZN(n4119) );
  OAI21_X1 U4234 ( .B1(n2511), .B2(n4146), .A(n4119), .ZN(\DataP/WB[16] ) );
  AOI22_X1 U4235 ( .A1(n4144), .A2(\DataP/LMD_out[17] ), .B1(n4143), .B2(
        \DataP/link_addr_W[17] ), .ZN(n4120) );
  OAI21_X1 U4236 ( .B1(n2493), .B2(n4146), .A(n4120), .ZN(\DataP/WB[17] ) );
  AOI22_X1 U4237 ( .A1(n4144), .A2(\DataP/LMD_out[18] ), .B1(n4143), .B2(
        \DataP/link_addr_W[18] ), .ZN(n4121) );
  OAI21_X1 U4238 ( .B1(n2505), .B2(n4146), .A(n4121), .ZN(\DataP/WB[18] ) );
  AOI22_X1 U4239 ( .A1(n3229), .A2(\DataP/LMD_out[19] ), .B1(n4143), .B2(
        \DataP/link_addr_W[19] ), .ZN(n4122) );
  OAI21_X1 U4240 ( .B1(n2498), .B2(n4146), .A(n4122), .ZN(\DataP/WB[19] ) );
  AOI22_X1 U4241 ( .A1(n3229), .A2(\DataP/LMD_out[1] ), .B1(n4143), .B2(
        \DataP/link_addr_W[1] ), .ZN(n4123) );
  OAI21_X1 U4242 ( .B1(n2522), .B2(n4146), .A(n4123), .ZN(\DataP/WB[1] ) );
  AOI22_X1 U4243 ( .A1(n3229), .A2(\DataP/LMD_out[20] ), .B1(n4143), .B2(
        \DataP/link_addr_W[20] ), .ZN(n4124) );
  OAI21_X1 U4244 ( .B1(n2506), .B2(n4146), .A(n4124), .ZN(\DataP/WB[20] ) );
  AOI22_X1 U4245 ( .A1(n3229), .A2(\DataP/LMD_out[21] ), .B1(n4143), .B2(
        \DataP/link_addr_W[21] ), .ZN(n4125) );
  OAI21_X1 U4246 ( .B1(n2499), .B2(n4146), .A(n4125), .ZN(\DataP/WB[21] ) );
  AOI22_X1 U4247 ( .A1(n3229), .A2(\DataP/LMD_out[22] ), .B1(n4143), .B2(
        \DataP/link_addr_W[22] ), .ZN(n4126) );
  OAI21_X1 U4248 ( .B1(n2512), .B2(n4146), .A(n4126), .ZN(\DataP/WB[22] ) );
  AOI22_X1 U4249 ( .A1(n3229), .A2(\DataP/LMD_out[23] ), .B1(n4143), .B2(
        \DataP/link_addr_W[23] ), .ZN(n4127) );
  OAI21_X1 U4250 ( .B1(n2494), .B2(n4146), .A(n4127), .ZN(\DataP/WB[23] ) );
  AOI22_X1 U4251 ( .A1(n3229), .A2(\DataP/LMD_out[24] ), .B1(n4143), .B2(
        \DataP/link_addr_W[24] ), .ZN(n4128) );
  OAI21_X1 U4252 ( .B1(n2513), .B2(n4146), .A(n4128), .ZN(\DataP/WB[24] ) );
  AOI22_X1 U4253 ( .A1(n3229), .A2(\DataP/LMD_out[25] ), .B1(n4143), .B2(
        \DataP/link_addr_W[25] ), .ZN(n4129) );
  OAI21_X1 U4254 ( .B1(n2507), .B2(n4146), .A(n4129), .ZN(\DataP/WB[25] ) );
  AOI22_X1 U4255 ( .A1(n3229), .A2(\DataP/LMD_out[26] ), .B1(n4143), .B2(
        \DataP/link_addr_W[26] ), .ZN(n4130) );
  OAI21_X1 U4256 ( .B1(n2500), .B2(n4146), .A(n4130), .ZN(\DataP/WB[26] ) );
  AOI22_X1 U4257 ( .A1(n3229), .A2(\DataP/LMD_out[27] ), .B1(n4143), .B2(
        \DataP/link_addr_W[27] ), .ZN(n4131) );
  OAI21_X1 U4258 ( .B1(n2495), .B2(n4146), .A(n4131), .ZN(\DataP/WB[27] ) );
  AOI22_X1 U4259 ( .A1(n4144), .A2(\DataP/LMD_out[28] ), .B1(n4143), .B2(
        \DataP/link_addr_W[28] ), .ZN(n4132) );
  OAI21_X1 U4260 ( .B1(n2508), .B2(n4146), .A(n4132), .ZN(\DataP/WB[28] ) );
  AOI22_X1 U4261 ( .A1(n4144), .A2(\DataP/LMD_out[29] ), .B1(n4143), .B2(
        \DataP/link_addr_W[29] ), .ZN(n4133) );
  OAI21_X1 U4262 ( .B1(n2501), .B2(n4146), .A(n4133), .ZN(\DataP/WB[29] ) );
  AOI22_X1 U4263 ( .A1(n4144), .A2(\DataP/LMD_out[2] ), .B1(n4143), .B2(
        \DataP/link_addr_W[2] ), .ZN(n4134) );
  OAI21_X1 U4264 ( .B1(n2514), .B2(n4146), .A(n4134), .ZN(\DataP/WB[2] ) );
  AOI22_X1 U4265 ( .A1(n4144), .A2(\DataP/LMD_out[30] ), .B1(n4143), .B2(
        \DataP/link_addr_W[30] ), .ZN(n4135) );
  OAI21_X1 U4266 ( .B1(n2496), .B2(n4146), .A(n4135), .ZN(\DataP/WB[30] ) );
  AOI22_X1 U4267 ( .A1(n4144), .A2(\DataP/LMD_out[31] ), .B1(n4143), .B2(
        \DataP/link_addr_W[31] ), .ZN(n4136) );
  OAI21_X1 U4268 ( .B1(n2517), .B2(n4146), .A(n4136), .ZN(\DataP/WB[31] ) );
  AOI22_X1 U4269 ( .A1(n4144), .A2(\DataP/LMD_out[3] ), .B1(n4143), .B2(
        \DataP/link_addr_W[3] ), .ZN(n4137) );
  OAI21_X1 U4270 ( .B1(n2523), .B2(n4146), .A(n4137), .ZN(\DataP/WB[3] ) );
  AOI22_X1 U4271 ( .A1(n4144), .A2(\DataP/LMD_out[4] ), .B1(n4143), .B2(
        \DataP/link_addr_W[4] ), .ZN(n4138) );
  OAI21_X1 U4272 ( .B1(n2509), .B2(n4146), .A(n4138), .ZN(\DataP/WB[4] ) );
  AOI22_X1 U4273 ( .A1(n3229), .A2(\DataP/LMD_out[5] ), .B1(n4143), .B2(
        \DataP/link_addr_W[5] ), .ZN(n4139) );
  OAI21_X1 U4274 ( .B1(n2520), .B2(n4146), .A(n4139), .ZN(\DataP/WB[5] ) );
  AOI22_X1 U4275 ( .A1(n4144), .A2(\DataP/LMD_out[6] ), .B1(n4143), .B2(
        \DataP/link_addr_W[6] ), .ZN(n4140) );
  OAI21_X1 U4276 ( .B1(n2515), .B2(n4146), .A(n4140), .ZN(\DataP/WB[6] ) );
  AOI22_X1 U4277 ( .A1(n3229), .A2(\DataP/LMD_out[7] ), .B1(n4143), .B2(
        \DataP/link_addr_W[7] ), .ZN(n4141) );
  OAI21_X1 U4278 ( .B1(n2510), .B2(n4146), .A(n4141), .ZN(\DataP/WB[7] ) );
  AOI22_X1 U4279 ( .A1(n4144), .A2(\DataP/LMD_out[8] ), .B1(n4143), .B2(
        \DataP/link_addr_W[8] ), .ZN(n4142) );
  OAI21_X1 U4280 ( .B1(n2502), .B2(n4146), .A(n4142), .ZN(\DataP/WB[8] ) );
  AOI22_X1 U4281 ( .A1(n3229), .A2(\DataP/LMD_out[9] ), .B1(n4143), .B2(
        \DataP/link_addr_W[9] ), .ZN(n4145) );
  OAI21_X1 U4282 ( .B1(n2519), .B2(n4146), .A(n4145), .ZN(\DataP/WB[9] ) );
  INV_X1 U4283 ( .A(n16), .ZN(n4152) );
  AOI211_X1 U4284 ( .C1(n607), .C2(n504), .A(\CU_I/cw[7] ), .B(n4153), .ZN(
        n4150) );
  OAI211_X1 U4285 ( .C1(n4152), .C2(n4151), .A(Rst), .B(n4150), .ZN(n4164) );
  AND2_X1 U4286 ( .A1(Rst), .A2(n4153), .ZN(n4162) );
  NOR2_X1 U4287 ( .A1(n4155), .A2(n4154), .ZN(n4165) );
  NAND2_X1 U4288 ( .A1(Rst), .A2(n4165), .ZN(n4179) );
  OAI22_X1 U4289 ( .A1(n497), .A2(n4179), .B1(n4156), .B2(n4164), .ZN(n4161)
         );
  AOI21_X1 U4290 ( .B1(n4162), .B2(\DataP/IR1[11] ), .A(n4161), .ZN(n4157) );
  OAI21_X1 U4291 ( .B1(n485), .B2(n4164), .A(n4157), .ZN(\DataP/dest_D[0] ) );
  AOI21_X1 U4292 ( .B1(n4162), .B2(\DataP/IR1[12] ), .A(n4161), .ZN(n4158) );
  OAI21_X1 U4293 ( .B1(n486), .B2(n4164), .A(n4158), .ZN(\DataP/dest_D[1] ) );
  AOI21_X1 U4294 ( .B1(n4162), .B2(\DataP/IR1[13] ), .A(n4161), .ZN(n4159) );
  OAI21_X1 U4295 ( .B1(n487), .B2(n4164), .A(n4159), .ZN(\DataP/dest_D[2] ) );
  AOI21_X1 U4296 ( .B1(n4162), .B2(\DataP/IR1[14] ), .A(n4161), .ZN(n4160) );
  OAI21_X1 U4297 ( .B1(n488), .B2(n4164), .A(n4160), .ZN(\DataP/dest_D[3] ) );
  AOI21_X1 U4298 ( .B1(n4162), .B2(\DataP/IR1[15] ), .A(n4161), .ZN(n4163) );
  OAI21_X1 U4299 ( .B1(n489), .B2(n4164), .A(n4163), .ZN(\DataP/dest_D[4] ) );
  NAND2_X1 U4300 ( .A1(IR_CU_28), .A2(n4166), .ZN(n4171) );
  OAI21_X1 U4301 ( .B1(n515), .B2(IR_CU_27), .A(n2374), .ZN(n4167) );
  AOI22_X1 U4302 ( .A1(n4168), .A2(n497), .B1(n1960), .B2(n4167), .ZN(n4169)
         );
  OAI221_X1 U4303 ( .B1(n514), .B2(n4171), .C1(n2374), .C2(n4170), .A(n4169), 
        .ZN(n4172) );
  AOI211_X1 U4304 ( .C1(IR_CU_27), .C2(n4174), .A(n4173), .B(n4172), .ZN(n4175) );
  OAI221_X1 U4305 ( .B1(IR_CU_31), .B2(n4177), .C1(n516), .C2(n4176), .A(n4175), .ZN(n4178) );
  NAND4_X1 U4306 ( .A1(Rst), .A2(\DataP/IR1[15] ), .A3(n4181), .A4(n4178), 
        .ZN(n4180) );
  OAI21_X1 U4307 ( .B1(n485), .B2(n4179), .A(n4180), .ZN(\DataP/imm_out[16] )
         );
  OAI21_X1 U4308 ( .B1(n486), .B2(n4179), .A(n4180), .ZN(\DataP/imm_out[17] )
         );
  OAI21_X1 U4309 ( .B1(n487), .B2(n4179), .A(n4180), .ZN(\DataP/imm_out[18] )
         );
  OAI21_X1 U4310 ( .B1(n488), .B2(n4179), .A(n4180), .ZN(\DataP/imm_out[19] )
         );
  OAI21_X1 U4311 ( .B1(n489), .B2(n4179), .A(n4180), .ZN(\DataP/imm_out[20] )
         );
  NAND2_X1 U4312 ( .A1(Rst), .A2(\DataP/IR1[21] ), .ZN(n4189) );
  OAI21_X1 U4313 ( .B1(n4181), .B2(n4189), .A(n4180), .ZN(\DataP/imm_out[21] )
         );
  NAND2_X1 U4314 ( .A1(Rst), .A2(\DataP/IR1[22] ), .ZN(n4188) );
  OAI21_X1 U4315 ( .B1(n4181), .B2(n4188), .A(n4180), .ZN(\DataP/imm_out[22] )
         );
  NAND2_X1 U4316 ( .A1(Rst), .A2(\DataP/IR1[23] ), .ZN(n4187) );
  OAI21_X1 U4317 ( .B1(n4181), .B2(n4187), .A(n4180), .ZN(\DataP/imm_out[23] )
         );
  NAND2_X1 U4318 ( .A1(Rst), .A2(\DataP/IR1[24] ), .ZN(n4186) );
  OAI21_X1 U4319 ( .B1(n4181), .B2(n4186), .A(n4180), .ZN(\DataP/imm_out[24] )
         );
  NAND2_X1 U4320 ( .A1(Rst), .A2(\DataP/IR1[25] ), .ZN(n4185) );
  OAI21_X1 U4321 ( .B1(n4181), .B2(n4185), .A(n4180), .ZN(\DataP/imm_out[31] )
         );
  MUX2_X1 U4322 ( .A(\DataP/pc_out_0 ), .B(\DataP/npc_pre[0] ), .S(n2132), .Z(
        \DataP/NPC_add/N1 ) );
  MUX2_X1 U4323 ( .A(\DataP/pc_out_1 ), .B(\DataP/npc_pre[1] ), .S(n2132), .Z(
        \DataP/NPC_add/N2 ) );
  MUX2_X1 U4324 ( .A(\DataP/link_addr_D[31] ), .B(\DataP/link_addr_F[31] ), 
        .S(n3230), .Z(n1481) );
  MUX2_X1 U4325 ( .A(\DataP/link_addr_D[0] ), .B(\DataP/link_addr_F[0] ), .S(
        n3230), .Z(n1480) );
  MUX2_X1 U4326 ( .A(\DataP/link_addr_D[1] ), .B(\DataP/link_addr_F[1] ), .S(
        n3230), .Z(n1479) );
  MUX2_X1 U4327 ( .A(\DataP/link_addr_D[2] ), .B(\DataP/link_addr_F[2] ), .S(
        n3230), .Z(n1478) );
  MUX2_X1 U4328 ( .A(\DataP/link_addr_D[3] ), .B(\DataP/link_addr_F[3] ), .S(
        n3230), .Z(n1477) );
  MUX2_X1 U4329 ( .A(\DataP/link_addr_D[4] ), .B(\DataP/link_addr_F[4] ), .S(
        n3230), .Z(n1476) );
  MUX2_X1 U4330 ( .A(\DataP/link_addr_D[5] ), .B(\DataP/link_addr_F[5] ), .S(
        n3230), .Z(n1475) );
  MUX2_X1 U4331 ( .A(\DataP/link_addr_D[6] ), .B(\DataP/link_addr_F[6] ), .S(
        n3230), .Z(n1474) );
  MUX2_X1 U4332 ( .A(\DataP/link_addr_D[7] ), .B(\DataP/link_addr_F[7] ), .S(
        n3230), .Z(n1473) );
  MUX2_X1 U4333 ( .A(\DataP/link_addr_D[8] ), .B(\DataP/link_addr_F[8] ), .S(
        n3230), .Z(n1472) );
  MUX2_X1 U4334 ( .A(\DataP/link_addr_D[9] ), .B(\DataP/link_addr_F[9] ), .S(
        n3230), .Z(n1471) );
  MUX2_X1 U4335 ( .A(\DataP/link_addr_D[10] ), .B(\DataP/link_addr_F[10] ), 
        .S(n3230), .Z(n1470) );
  MUX2_X1 U4336 ( .A(\DataP/link_addr_D[11] ), .B(\DataP/link_addr_F[11] ), 
        .S(n3231), .Z(n1469) );
  MUX2_X1 U4337 ( .A(\DataP/link_addr_D[12] ), .B(\DataP/link_addr_F[12] ), 
        .S(n3231), .Z(n1468) );
  MUX2_X1 U4338 ( .A(\DataP/link_addr_D[13] ), .B(\DataP/link_addr_F[13] ), 
        .S(n3231), .Z(n1467) );
  MUX2_X1 U4339 ( .A(\DataP/link_addr_D[14] ), .B(\DataP/link_addr_F[14] ), 
        .S(n3231), .Z(n1466) );
  MUX2_X1 U4340 ( .A(\DataP/link_addr_D[15] ), .B(\DataP/link_addr_F[15] ), 
        .S(n3231), .Z(n1465) );
  MUX2_X1 U4341 ( .A(\DataP/link_addr_D[16] ), .B(\DataP/link_addr_F[16] ), 
        .S(n3231), .Z(n1464) );
  MUX2_X1 U4342 ( .A(\DataP/link_addr_D[17] ), .B(\DataP/link_addr_F[17] ), 
        .S(n3231), .Z(n1463) );
  MUX2_X1 U4343 ( .A(\DataP/link_addr_D[18] ), .B(\DataP/link_addr_F[18] ), 
        .S(n3231), .Z(n1462) );
  MUX2_X1 U4344 ( .A(\DataP/link_addr_D[19] ), .B(\DataP/link_addr_F[19] ), 
        .S(n3231), .Z(n1461) );
  MUX2_X1 U4345 ( .A(\DataP/link_addr_D[20] ), .B(\DataP/link_addr_F[20] ), 
        .S(n3231), .Z(n1460) );
  MUX2_X1 U4346 ( .A(\DataP/link_addr_D[21] ), .B(\DataP/link_addr_F[21] ), 
        .S(n3231), .Z(n1459) );
  MUX2_X1 U4347 ( .A(\DataP/link_addr_D[22] ), .B(\DataP/link_addr_F[22] ), 
        .S(n3231), .Z(n1458) );
  MUX2_X1 U4348 ( .A(\DataP/link_addr_D[23] ), .B(\DataP/link_addr_F[23] ), 
        .S(n3230), .Z(n1457) );
  MUX2_X1 U4349 ( .A(\DataP/link_addr_D[24] ), .B(\DataP/link_addr_F[24] ), 
        .S(n3231), .Z(n1456) );
  MUX2_X1 U4350 ( .A(\DataP/link_addr_D[25] ), .B(\DataP/link_addr_F[25] ), 
        .S(n3230), .Z(n1455) );
  MUX2_X1 U4351 ( .A(\DataP/link_addr_D[26] ), .B(\DataP/link_addr_F[26] ), 
        .S(n3231), .Z(n1454) );
  MUX2_X1 U4352 ( .A(\DataP/link_addr_D[27] ), .B(\DataP/link_addr_F[27] ), 
        .S(n3230), .Z(n1453) );
  MUX2_X1 U4353 ( .A(\DataP/link_addr_D[28] ), .B(\DataP/link_addr_F[28] ), 
        .S(n3231), .Z(n1452) );
  MUX2_X1 U4354 ( .A(\DataP/link_addr_D[29] ), .B(\DataP/link_addr_F[29] ), 
        .S(n3230), .Z(n1451) );
  MUX2_X1 U4355 ( .A(\DataP/link_addr_D[30] ), .B(\DataP/link_addr_F[30] ), 
        .S(n3231), .Z(n1450) );
  MUX2_X1 U4356 ( .A(\DataP/pr_D ), .B(\DataP/prediction ), .S(n3230), .Z(
        n1449) );
  NAND2_X1 U4357 ( .A1(\DataP/npc[31] ), .A2(n3232), .ZN(n163) );
  AOI21_X1 U4358 ( .B1(n4191), .B2(n2104), .A(n3235), .ZN(n162) );
  NAND2_X1 U4359 ( .A1(\DataP/npc[30] ), .A2(n3232), .ZN(n159) );
  AOI21_X1 U4360 ( .B1(n4192), .B2(n2104), .A(n3235), .ZN(n158) );
  NAND2_X1 U4361 ( .A1(\DataP/npc[29] ), .A2(n3232), .ZN(n155) );
  AOI21_X1 U4362 ( .B1(n4193), .B2(n2104), .A(n3235), .ZN(n154) );
  NAND2_X1 U4363 ( .A1(\DataP/npc[28] ), .A2(n3232), .ZN(n151) );
  AOI21_X1 U4364 ( .B1(n4194), .B2(n2104), .A(n3235), .ZN(n150) );
  NAND2_X1 U4365 ( .A1(\DataP/npc[27] ), .A2(n3232), .ZN(n147) );
  AOI21_X1 U4366 ( .B1(n4195), .B2(n2104), .A(n3235), .ZN(n146) );
  NAND2_X1 U4367 ( .A1(\DataP/npc[26] ), .A2(n3232), .ZN(n143) );
  AOI21_X1 U4368 ( .B1(n4196), .B2(n2104), .A(n3235), .ZN(n142) );
  NAND2_X1 U4369 ( .A1(\DataP/npc[25] ), .A2(n3232), .ZN(n139) );
  AOI21_X1 U4370 ( .B1(n4197), .B2(n2104), .A(n3235), .ZN(n138) );
  NAND2_X1 U4371 ( .A1(\DataP/npc[24] ), .A2(n3232), .ZN(n135) );
  AOI21_X1 U4372 ( .B1(n4198), .B2(n2104), .A(n3235), .ZN(n134) );
  NAND2_X1 U4373 ( .A1(\DataP/npc[23] ), .A2(n3232), .ZN(n131) );
  AOI21_X1 U4374 ( .B1(n4199), .B2(n2104), .A(n3235), .ZN(n130) );
  NAND2_X1 U4375 ( .A1(\DataP/npc[22] ), .A2(n3232), .ZN(n127) );
  AOI21_X1 U4376 ( .B1(n4200), .B2(n2104), .A(n3235), .ZN(n126) );
  NAND2_X1 U4377 ( .A1(\DataP/npc[21] ), .A2(n4222), .ZN(n123) );
  AOI21_X1 U4378 ( .B1(n4201), .B2(n2104), .A(n3235), .ZN(n122) );
  NAND2_X1 U4379 ( .A1(\DataP/npc[20] ), .A2(n4222), .ZN(n119) );
  AOI21_X1 U4380 ( .B1(n4202), .B2(n2104), .A(n3236), .ZN(n118) );
  NAND2_X1 U4381 ( .A1(\DataP/npc[19] ), .A2(n4222), .ZN(n115) );
  AOI21_X1 U4382 ( .B1(n4203), .B2(n2104), .A(n3235), .ZN(n114) );
  NAND2_X1 U4383 ( .A1(\DataP/npc[18] ), .A2(n3232), .ZN(n111) );
  AOI21_X1 U4384 ( .B1(n4204), .B2(n2104), .A(n3235), .ZN(n110) );
  NAND2_X1 U4385 ( .A1(\DataP/npc[17] ), .A2(n4222), .ZN(n107) );
  AOI21_X1 U4386 ( .B1(n4205), .B2(n2104), .A(n3235), .ZN(n106) );
  NAND2_X1 U4387 ( .A1(\DataP/npc[16] ), .A2(n3232), .ZN(n103) );
  AOI21_X1 U4388 ( .B1(n4206), .B2(n2104), .A(n3236), .ZN(n102) );
  NAND2_X1 U4389 ( .A1(\DataP/npc[15] ), .A2(n4222), .ZN(n99) );
  AOI21_X1 U4390 ( .B1(n4207), .B2(n2104), .A(n3236), .ZN(n98) );
  NAND2_X1 U4391 ( .A1(\DataP/npc[14] ), .A2(n3232), .ZN(n95) );
  AOI21_X1 U4392 ( .B1(n4208), .B2(n2104), .A(n3236), .ZN(n94) );
  NAND2_X1 U4393 ( .A1(\DataP/npc[13] ), .A2(n4222), .ZN(n91) );
  AOI21_X1 U4394 ( .B1(n4209), .B2(n2104), .A(n3236), .ZN(n90) );
  NAND2_X1 U4395 ( .A1(\DataP/npc[12] ), .A2(n4222), .ZN(n87) );
  AOI21_X1 U4396 ( .B1(n4210), .B2(n2104), .A(n3236), .ZN(n86) );
  NAND2_X1 U4397 ( .A1(\DataP/npc[11] ), .A2(n4222), .ZN(n83) );
  AOI21_X1 U4398 ( .B1(n4211), .B2(n2104), .A(n3236), .ZN(n82) );
  NAND2_X1 U4399 ( .A1(\DataP/npc[10] ), .A2(n4222), .ZN(n79) );
  AOI21_X1 U4400 ( .B1(n4212), .B2(n2104), .A(n3236), .ZN(n78) );
  NAND2_X1 U4401 ( .A1(\DataP/npc[9] ), .A2(n4222), .ZN(n75) );
  AOI21_X1 U4402 ( .B1(n4213), .B2(n2104), .A(n3236), .ZN(n74) );
  NAND2_X1 U4403 ( .A1(\DataP/npc[8] ), .A2(n4222), .ZN(n71) );
  AOI21_X1 U4404 ( .B1(n4214), .B2(n2104), .A(n3236), .ZN(n70) );
  NAND2_X1 U4405 ( .A1(\DataP/npc[7] ), .A2(n3232), .ZN(n67) );
  AOI21_X1 U4406 ( .B1(n4215), .B2(n2104), .A(n3236), .ZN(n66) );
  NAND2_X1 U4407 ( .A1(\DataP/npc[6] ), .A2(n3232), .ZN(n63) );
  AOI21_X1 U4408 ( .B1(n4216), .B2(n2104), .A(n3236), .ZN(n62) );
  NAND2_X1 U4409 ( .A1(\DataP/npc[5] ), .A2(n3232), .ZN(n59) );
  AOI21_X1 U4410 ( .B1(n4217), .B2(n2104), .A(n3236), .ZN(n58) );
  NAND2_X1 U4411 ( .A1(\DataP/npc[4] ), .A2(n3232), .ZN(n55) );
  AOI21_X1 U4412 ( .B1(n4218), .B2(n2104), .A(n3236), .ZN(n54) );
  NAND2_X1 U4413 ( .A1(\DataP/npc[3] ), .A2(n3232), .ZN(n51) );
  AOI21_X1 U4414 ( .B1(n4219), .B2(n2104), .A(n3236), .ZN(n50) );
  NAND2_X1 U4415 ( .A1(\DataP/npc[2] ), .A2(n3232), .ZN(n47) );
  AOI21_X1 U4416 ( .B1(n4220), .B2(n2104), .A(n3236), .ZN(n46) );
  NAND2_X1 U4417 ( .A1(\DataP/npc[1] ), .A2(n3232), .ZN(n43) );
  AOI21_X1 U4418 ( .B1(n4221), .B2(n2104), .A(n3236), .ZN(n42) );
  NAND2_X1 U4419 ( .A1(\DataP/npc[0] ), .A2(n3232), .ZN(n39) );
  AOI21_X1 U4420 ( .B1(n4223), .B2(n2104), .A(n3235), .ZN(n38) );
endmodule

