
module register_file_N32_addBit5 ( RESET, RE, WE, ADD_WR, ADD_RDA, ADD_RDB, 
        DATAIN, OUTA, OUTB );
  input [4:0] ADD_WR;
  input [4:0] ADD_RDA;
  input [4:0] ADD_RDB;
  input [31:0] DATAIN;
  output [31:0] OUTA;
  output [31:0] OUTB;
  input RESET, RE, WE;
  wire   \REGISTERS[1][31] , \REGISTERS[1][30] , \REGISTERS[1][29] ,
         \REGISTERS[1][28] , \REGISTERS[1][27] , \REGISTERS[1][26] ,
         \REGISTERS[1][25] , \REGISTERS[1][24] , \REGISTERS[1][23] ,
         \REGISTERS[1][22] , \REGISTERS[1][21] , \REGISTERS[1][20] ,
         \REGISTERS[1][19] , \REGISTERS[1][18] , \REGISTERS[1][17] ,
         \REGISTERS[1][16] , \REGISTERS[1][15] , \REGISTERS[1][14] ,
         \REGISTERS[1][13] , \REGISTERS[1][12] , \REGISTERS[1][11] ,
         \REGISTERS[1][10] , \REGISTERS[1][9] , \REGISTERS[1][8] ,
         \REGISTERS[1][7] , \REGISTERS[1][6] , \REGISTERS[1][5] ,
         \REGISTERS[1][4] , \REGISTERS[1][3] , \REGISTERS[1][2] ,
         \REGISTERS[1][1] , \REGISTERS[1][0] , \REGISTERS[2][31] ,
         \REGISTERS[2][30] , \REGISTERS[2][29] , \REGISTERS[2][28] ,
         \REGISTERS[2][27] , \REGISTERS[2][26] , \REGISTERS[2][25] ,
         \REGISTERS[2][24] , \REGISTERS[2][23] , \REGISTERS[2][22] ,
         \REGISTERS[2][21] , \REGISTERS[2][20] , \REGISTERS[2][19] ,
         \REGISTERS[2][18] , \REGISTERS[2][17] , \REGISTERS[2][16] ,
         \REGISTERS[2][15] , \REGISTERS[2][14] , \REGISTERS[2][13] ,
         \REGISTERS[2][12] , \REGISTERS[2][11] , \REGISTERS[2][10] ,
         \REGISTERS[2][9] , \REGISTERS[2][8] , \REGISTERS[2][7] ,
         \REGISTERS[2][6] , \REGISTERS[2][5] , \REGISTERS[2][4] ,
         \REGISTERS[2][3] , \REGISTERS[2][2] , \REGISTERS[2][1] ,
         \REGISTERS[2][0] , \REGISTERS[3][31] , \REGISTERS[3][30] ,
         \REGISTERS[3][29] , \REGISTERS[3][28] , \REGISTERS[3][27] ,
         \REGISTERS[3][26] , \REGISTERS[3][25] , \REGISTERS[3][24] ,
         \REGISTERS[3][23] , \REGISTERS[3][22] , \REGISTERS[3][21] ,
         \REGISTERS[3][20] , \REGISTERS[3][19] , \REGISTERS[3][18] ,
         \REGISTERS[3][17] , \REGISTERS[3][16] , \REGISTERS[3][15] ,
         \REGISTERS[3][14] , \REGISTERS[3][13] , \REGISTERS[3][12] ,
         \REGISTERS[3][11] , \REGISTERS[3][10] , \REGISTERS[3][9] ,
         \REGISTERS[3][8] , \REGISTERS[3][7] , \REGISTERS[3][6] ,
         \REGISTERS[3][5] , \REGISTERS[3][4] , \REGISTERS[3][3] ,
         \REGISTERS[3][2] , \REGISTERS[3][1] , \REGISTERS[3][0] ,
         \REGISTERS[4][31] , \REGISTERS[4][30] , \REGISTERS[4][29] ,
         \REGISTERS[4][28] , \REGISTERS[4][27] , \REGISTERS[4][26] ,
         \REGISTERS[4][25] , \REGISTERS[4][24] , \REGISTERS[4][23] ,
         \REGISTERS[4][22] , \REGISTERS[4][21] , \REGISTERS[4][20] ,
         \REGISTERS[4][19] , \REGISTERS[4][18] , \REGISTERS[4][17] ,
         \REGISTERS[4][16] , \REGISTERS[4][15] , \REGISTERS[4][14] ,
         \REGISTERS[4][13] , \REGISTERS[4][12] , \REGISTERS[4][11] ,
         \REGISTERS[4][10] , \REGISTERS[4][9] , \REGISTERS[4][8] ,
         \REGISTERS[4][7] , \REGISTERS[4][6] , \REGISTERS[4][5] ,
         \REGISTERS[4][4] , \REGISTERS[4][3] , \REGISTERS[4][2] ,
         \REGISTERS[4][1] , \REGISTERS[4][0] , \REGISTERS[5][31] ,
         \REGISTERS[5][30] , \REGISTERS[5][29] , \REGISTERS[5][28] ,
         \REGISTERS[5][27] , \REGISTERS[5][26] , \REGISTERS[5][25] ,
         \REGISTERS[5][24] , \REGISTERS[5][23] , \REGISTERS[5][22] ,
         \REGISTERS[5][21] , \REGISTERS[5][20] , \REGISTERS[5][19] ,
         \REGISTERS[5][18] , \REGISTERS[5][17] , \REGISTERS[5][16] ,
         \REGISTERS[5][15] , \REGISTERS[5][14] , \REGISTERS[5][13] ,
         \REGISTERS[5][12] , \REGISTERS[5][11] , \REGISTERS[5][10] ,
         \REGISTERS[5][9] , \REGISTERS[5][8] , \REGISTERS[5][7] ,
         \REGISTERS[5][6] , \REGISTERS[5][5] , \REGISTERS[5][4] ,
         \REGISTERS[5][3] , \REGISTERS[5][2] , \REGISTERS[5][1] ,
         \REGISTERS[5][0] , \REGISTERS[6][31] , \REGISTERS[6][30] ,
         \REGISTERS[6][29] , \REGISTERS[6][28] , \REGISTERS[6][27] ,
         \REGISTERS[6][26] , \REGISTERS[6][25] , \REGISTERS[6][24] ,
         \REGISTERS[6][23] , \REGISTERS[6][22] , \REGISTERS[6][21] ,
         \REGISTERS[6][20] , \REGISTERS[6][19] , \REGISTERS[6][18] ,
         \REGISTERS[6][17] , \REGISTERS[6][16] , \REGISTERS[6][15] ,
         \REGISTERS[6][14] , \REGISTERS[6][13] , \REGISTERS[6][12] ,
         \REGISTERS[6][11] , \REGISTERS[6][10] , \REGISTERS[6][9] ,
         \REGISTERS[6][8] , \REGISTERS[6][7] , \REGISTERS[6][6] ,
         \REGISTERS[6][5] , \REGISTERS[6][4] , \REGISTERS[6][3] ,
         \REGISTERS[6][2] , \REGISTERS[6][1] , \REGISTERS[6][0] ,
         \REGISTERS[7][31] , \REGISTERS[7][30] , \REGISTERS[7][29] ,
         \REGISTERS[7][28] , \REGISTERS[7][27] , \REGISTERS[7][26] ,
         \REGISTERS[7][25] , \REGISTERS[7][24] , \REGISTERS[7][23] ,
         \REGISTERS[7][22] , \REGISTERS[7][21] , \REGISTERS[7][20] ,
         \REGISTERS[7][19] , \REGISTERS[7][18] , \REGISTERS[7][17] ,
         \REGISTERS[7][16] , \REGISTERS[7][15] , \REGISTERS[7][14] ,
         \REGISTERS[7][13] , \REGISTERS[7][12] , \REGISTERS[7][11] ,
         \REGISTERS[7][10] , \REGISTERS[7][9] , \REGISTERS[7][8] ,
         \REGISTERS[7][7] , \REGISTERS[7][6] , \REGISTERS[7][5] ,
         \REGISTERS[7][4] , \REGISTERS[7][3] , \REGISTERS[7][2] ,
         \REGISTERS[7][1] , \REGISTERS[7][0] , \REGISTERS[8][31] ,
         \REGISTERS[8][30] , \REGISTERS[8][29] , \REGISTERS[8][28] ,
         \REGISTERS[8][27] , \REGISTERS[8][26] , \REGISTERS[8][25] ,
         \REGISTERS[8][24] , \REGISTERS[8][23] , \REGISTERS[8][22] ,
         \REGISTERS[8][21] , \REGISTERS[8][20] , \REGISTERS[8][19] ,
         \REGISTERS[8][18] , \REGISTERS[8][17] , \REGISTERS[8][16] ,
         \REGISTERS[8][15] , \REGISTERS[8][14] , \REGISTERS[8][13] ,
         \REGISTERS[8][12] , \REGISTERS[8][11] , \REGISTERS[8][10] ,
         \REGISTERS[8][9] , \REGISTERS[8][8] , \REGISTERS[8][7] ,
         \REGISTERS[8][6] , \REGISTERS[8][5] , \REGISTERS[8][4] ,
         \REGISTERS[8][3] , \REGISTERS[8][2] , \REGISTERS[8][1] ,
         \REGISTERS[8][0] , \REGISTERS[9][31] , \REGISTERS[9][30] ,
         \REGISTERS[9][29] , \REGISTERS[9][28] , \REGISTERS[9][27] ,
         \REGISTERS[9][26] , \REGISTERS[9][25] , \REGISTERS[9][24] ,
         \REGISTERS[9][23] , \REGISTERS[9][22] , \REGISTERS[9][21] ,
         \REGISTERS[9][20] , \REGISTERS[9][19] , \REGISTERS[9][18] ,
         \REGISTERS[9][17] , \REGISTERS[9][16] , \REGISTERS[9][15] ,
         \REGISTERS[9][14] , \REGISTERS[9][13] , \REGISTERS[9][12] ,
         \REGISTERS[9][11] , \REGISTERS[9][10] , \REGISTERS[9][9] ,
         \REGISTERS[9][8] , \REGISTERS[9][7] , \REGISTERS[9][6] ,
         \REGISTERS[9][5] , \REGISTERS[9][4] , \REGISTERS[9][3] ,
         \REGISTERS[9][2] , \REGISTERS[9][1] , \REGISTERS[9][0] ,
         \REGISTERS[10][31] , \REGISTERS[10][30] , \REGISTERS[10][29] ,
         \REGISTERS[10][28] , \REGISTERS[10][27] , \REGISTERS[10][26] ,
         \REGISTERS[10][25] , \REGISTERS[10][24] , \REGISTERS[10][23] ,
         \REGISTERS[10][22] , \REGISTERS[10][21] , \REGISTERS[10][20] ,
         \REGISTERS[10][19] , \REGISTERS[10][18] , \REGISTERS[10][17] ,
         \REGISTERS[10][16] , \REGISTERS[10][15] , \REGISTERS[10][14] ,
         \REGISTERS[10][13] , \REGISTERS[10][12] , \REGISTERS[10][11] ,
         \REGISTERS[10][10] , \REGISTERS[10][9] , \REGISTERS[10][8] ,
         \REGISTERS[10][7] , \REGISTERS[10][6] , \REGISTERS[10][5] ,
         \REGISTERS[10][4] , \REGISTERS[10][3] , \REGISTERS[10][2] ,
         \REGISTERS[10][1] , \REGISTERS[10][0] , \REGISTERS[11][31] ,
         \REGISTERS[11][30] , \REGISTERS[11][29] , \REGISTERS[11][28] ,
         \REGISTERS[11][27] , \REGISTERS[11][26] , \REGISTERS[11][25] ,
         \REGISTERS[11][24] , \REGISTERS[11][23] , \REGISTERS[11][22] ,
         \REGISTERS[11][21] , \REGISTERS[11][20] , \REGISTERS[11][19] ,
         \REGISTERS[11][18] , \REGISTERS[11][17] , \REGISTERS[11][16] ,
         \REGISTERS[11][15] , \REGISTERS[11][14] , \REGISTERS[11][13] ,
         \REGISTERS[11][12] , \REGISTERS[11][11] , \REGISTERS[11][10] ,
         \REGISTERS[11][9] , \REGISTERS[11][8] , \REGISTERS[11][7] ,
         \REGISTERS[11][6] , \REGISTERS[11][5] , \REGISTERS[11][4] ,
         \REGISTERS[11][3] , \REGISTERS[11][2] , \REGISTERS[11][1] ,
         \REGISTERS[11][0] , \REGISTERS[12][31] , \REGISTERS[12][30] ,
         \REGISTERS[12][29] , \REGISTERS[12][28] , \REGISTERS[12][27] ,
         \REGISTERS[12][26] , \REGISTERS[12][25] , \REGISTERS[12][24] ,
         \REGISTERS[12][23] , \REGISTERS[12][22] , \REGISTERS[12][21] ,
         \REGISTERS[12][20] , \REGISTERS[12][19] , \REGISTERS[12][18] ,
         \REGISTERS[12][17] , \REGISTERS[12][16] , \REGISTERS[12][15] ,
         \REGISTERS[12][14] , \REGISTERS[12][13] , \REGISTERS[12][12] ,
         \REGISTERS[12][11] , \REGISTERS[12][10] , \REGISTERS[12][9] ,
         \REGISTERS[12][8] , \REGISTERS[12][7] , \REGISTERS[12][6] ,
         \REGISTERS[12][5] , \REGISTERS[12][4] , \REGISTERS[12][3] ,
         \REGISTERS[12][2] , \REGISTERS[12][1] , \REGISTERS[12][0] ,
         \REGISTERS[13][31] , \REGISTERS[13][30] , \REGISTERS[13][29] ,
         \REGISTERS[13][28] , \REGISTERS[13][27] , \REGISTERS[13][26] ,
         \REGISTERS[13][25] , \REGISTERS[13][24] , \REGISTERS[13][23] ,
         \REGISTERS[13][22] , \REGISTERS[13][21] , \REGISTERS[13][20] ,
         \REGISTERS[13][19] , \REGISTERS[13][18] , \REGISTERS[13][17] ,
         \REGISTERS[13][16] , \REGISTERS[13][15] , \REGISTERS[13][14] ,
         \REGISTERS[13][13] , \REGISTERS[13][12] , \REGISTERS[13][11] ,
         \REGISTERS[13][10] , \REGISTERS[13][9] , \REGISTERS[13][8] ,
         \REGISTERS[13][7] , \REGISTERS[13][6] , \REGISTERS[13][5] ,
         \REGISTERS[13][4] , \REGISTERS[13][3] , \REGISTERS[13][2] ,
         \REGISTERS[13][1] , \REGISTERS[13][0] , \REGISTERS[14][31] ,
         \REGISTERS[14][30] , \REGISTERS[14][29] , \REGISTERS[14][28] ,
         \REGISTERS[14][27] , \REGISTERS[14][26] , \REGISTERS[14][25] ,
         \REGISTERS[14][24] , \REGISTERS[14][23] , \REGISTERS[14][22] ,
         \REGISTERS[14][21] , \REGISTERS[14][20] , \REGISTERS[14][19] ,
         \REGISTERS[14][18] , \REGISTERS[14][17] , \REGISTERS[14][16] ,
         \REGISTERS[14][15] , \REGISTERS[14][14] , \REGISTERS[14][13] ,
         \REGISTERS[14][12] , \REGISTERS[14][11] , \REGISTERS[14][10] ,
         \REGISTERS[14][9] , \REGISTERS[14][8] , \REGISTERS[14][7] ,
         \REGISTERS[14][6] , \REGISTERS[14][5] , \REGISTERS[14][4] ,
         \REGISTERS[14][3] , \REGISTERS[14][2] , \REGISTERS[14][1] ,
         \REGISTERS[14][0] , \REGISTERS[15][31] , \REGISTERS[15][30] ,
         \REGISTERS[15][29] , \REGISTERS[15][28] , \REGISTERS[15][27] ,
         \REGISTERS[15][26] , \REGISTERS[15][25] , \REGISTERS[15][24] ,
         \REGISTERS[15][23] , \REGISTERS[15][22] , \REGISTERS[15][21] ,
         \REGISTERS[15][20] , \REGISTERS[15][19] , \REGISTERS[15][18] ,
         \REGISTERS[15][17] , \REGISTERS[15][16] , \REGISTERS[15][15] ,
         \REGISTERS[15][14] , \REGISTERS[15][13] , \REGISTERS[15][12] ,
         \REGISTERS[15][11] , \REGISTERS[15][10] , \REGISTERS[15][9] ,
         \REGISTERS[15][8] , \REGISTERS[15][7] , \REGISTERS[15][6] ,
         \REGISTERS[15][5] , \REGISTERS[15][4] , \REGISTERS[15][3] ,
         \REGISTERS[15][2] , \REGISTERS[15][1] , \REGISTERS[15][0] ,
         \REGISTERS[16][31] , \REGISTERS[16][30] , \REGISTERS[16][29] ,
         \REGISTERS[16][28] , \REGISTERS[16][27] , \REGISTERS[16][26] ,
         \REGISTERS[16][25] , \REGISTERS[16][24] , \REGISTERS[16][23] ,
         \REGISTERS[16][22] , \REGISTERS[16][21] , \REGISTERS[16][20] ,
         \REGISTERS[16][19] , \REGISTERS[16][18] , \REGISTERS[16][17] ,
         \REGISTERS[16][16] , \REGISTERS[16][15] , \REGISTERS[16][14] ,
         \REGISTERS[16][13] , \REGISTERS[16][12] , \REGISTERS[16][11] ,
         \REGISTERS[16][10] , \REGISTERS[16][9] , \REGISTERS[16][8] ,
         \REGISTERS[16][7] , \REGISTERS[16][6] , \REGISTERS[16][5] ,
         \REGISTERS[16][4] , \REGISTERS[16][3] , \REGISTERS[16][2] ,
         \REGISTERS[16][1] , \REGISTERS[16][0] , \REGISTERS[17][31] ,
         \REGISTERS[17][30] , \REGISTERS[17][29] , \REGISTERS[17][28] ,
         \REGISTERS[17][27] , \REGISTERS[17][26] , \REGISTERS[17][25] ,
         \REGISTERS[17][24] , \REGISTERS[17][23] , \REGISTERS[17][22] ,
         \REGISTERS[17][21] , \REGISTERS[17][20] , \REGISTERS[17][19] ,
         \REGISTERS[17][18] , \REGISTERS[17][17] , \REGISTERS[17][16] ,
         \REGISTERS[17][15] , \REGISTERS[17][14] , \REGISTERS[17][13] ,
         \REGISTERS[17][12] , \REGISTERS[17][11] , \REGISTERS[17][10] ,
         \REGISTERS[17][9] , \REGISTERS[17][8] , \REGISTERS[17][7] ,
         \REGISTERS[17][6] , \REGISTERS[17][5] , \REGISTERS[17][4] ,
         \REGISTERS[17][3] , \REGISTERS[17][2] , \REGISTERS[17][1] ,
         \REGISTERS[17][0] , \REGISTERS[18][31] , \REGISTERS[18][30] ,
         \REGISTERS[18][29] , \REGISTERS[18][28] , \REGISTERS[18][27] ,
         \REGISTERS[18][26] , \REGISTERS[18][25] , \REGISTERS[18][24] ,
         \REGISTERS[18][23] , \REGISTERS[18][22] , \REGISTERS[18][21] ,
         \REGISTERS[18][20] , \REGISTERS[18][19] , \REGISTERS[18][18] ,
         \REGISTERS[18][17] , \REGISTERS[18][16] , \REGISTERS[18][15] ,
         \REGISTERS[18][14] , \REGISTERS[18][13] , \REGISTERS[18][12] ,
         \REGISTERS[18][11] , \REGISTERS[18][10] , \REGISTERS[18][9] ,
         \REGISTERS[18][8] , \REGISTERS[18][7] , \REGISTERS[18][6] ,
         \REGISTERS[18][5] , \REGISTERS[18][4] , \REGISTERS[18][3] ,
         \REGISTERS[18][2] , \REGISTERS[18][1] , \REGISTERS[18][0] ,
         \REGISTERS[19][31] , \REGISTERS[19][30] , \REGISTERS[19][29] ,
         \REGISTERS[19][28] , \REGISTERS[19][27] , \REGISTERS[19][26] ,
         \REGISTERS[19][25] , \REGISTERS[19][24] , \REGISTERS[19][23] ,
         \REGISTERS[19][22] , \REGISTERS[19][21] , \REGISTERS[19][20] ,
         \REGISTERS[19][19] , \REGISTERS[19][18] , \REGISTERS[19][17] ,
         \REGISTERS[19][16] , \REGISTERS[19][15] , \REGISTERS[19][14] ,
         \REGISTERS[19][13] , \REGISTERS[19][12] , \REGISTERS[19][11] ,
         \REGISTERS[19][10] , \REGISTERS[19][9] , \REGISTERS[19][8] ,
         \REGISTERS[19][7] , \REGISTERS[19][6] , \REGISTERS[19][5] ,
         \REGISTERS[19][4] , \REGISTERS[19][3] , \REGISTERS[19][2] ,
         \REGISTERS[19][1] , \REGISTERS[19][0] , \REGISTERS[20][31] ,
         \REGISTERS[20][30] , \REGISTERS[20][29] , \REGISTERS[20][28] ,
         \REGISTERS[20][27] , \REGISTERS[20][26] , \REGISTERS[20][25] ,
         \REGISTERS[20][24] , \REGISTERS[20][23] , \REGISTERS[20][22] ,
         \REGISTERS[20][21] , \REGISTERS[20][20] , \REGISTERS[20][19] ,
         \REGISTERS[20][18] , \REGISTERS[20][17] , \REGISTERS[20][16] ,
         \REGISTERS[20][15] , \REGISTERS[20][14] , \REGISTERS[20][13] ,
         \REGISTERS[20][12] , \REGISTERS[20][11] , \REGISTERS[20][10] ,
         \REGISTERS[20][9] , \REGISTERS[20][8] , \REGISTERS[20][7] ,
         \REGISTERS[20][6] , \REGISTERS[20][5] , \REGISTERS[20][4] ,
         \REGISTERS[20][3] , \REGISTERS[20][2] , \REGISTERS[20][1] ,
         \REGISTERS[20][0] , \REGISTERS[21][31] , \REGISTERS[21][30] ,
         \REGISTERS[21][29] , \REGISTERS[21][28] , \REGISTERS[21][27] ,
         \REGISTERS[21][26] , \REGISTERS[21][25] , \REGISTERS[21][24] ,
         \REGISTERS[21][23] , \REGISTERS[21][22] , \REGISTERS[21][21] ,
         \REGISTERS[21][20] , \REGISTERS[21][19] , \REGISTERS[21][18] ,
         \REGISTERS[21][17] , \REGISTERS[21][16] , \REGISTERS[21][15] ,
         \REGISTERS[21][14] , \REGISTERS[21][13] , \REGISTERS[21][12] ,
         \REGISTERS[21][11] , \REGISTERS[21][10] , \REGISTERS[21][9] ,
         \REGISTERS[21][8] , \REGISTERS[21][7] , \REGISTERS[21][6] ,
         \REGISTERS[21][5] , \REGISTERS[21][4] , \REGISTERS[21][3] ,
         \REGISTERS[21][2] , \REGISTERS[21][1] , \REGISTERS[21][0] ,
         \REGISTERS[22][31] , \REGISTERS[22][30] , \REGISTERS[22][29] ,
         \REGISTERS[22][28] , \REGISTERS[22][27] , \REGISTERS[22][26] ,
         \REGISTERS[22][25] , \REGISTERS[22][24] , \REGISTERS[22][23] ,
         \REGISTERS[22][22] , \REGISTERS[22][21] , \REGISTERS[22][20] ,
         \REGISTERS[22][19] , \REGISTERS[22][18] , \REGISTERS[22][17] ,
         \REGISTERS[22][16] , \REGISTERS[22][15] , \REGISTERS[22][14] ,
         \REGISTERS[22][13] , \REGISTERS[22][12] , \REGISTERS[22][11] ,
         \REGISTERS[22][10] , \REGISTERS[22][9] , \REGISTERS[22][8] ,
         \REGISTERS[22][7] , \REGISTERS[22][6] , \REGISTERS[22][5] ,
         \REGISTERS[22][4] , \REGISTERS[22][3] , \REGISTERS[22][2] ,
         \REGISTERS[22][1] , \REGISTERS[22][0] , \REGISTERS[23][31] ,
         \REGISTERS[23][30] , \REGISTERS[23][29] , \REGISTERS[23][28] ,
         \REGISTERS[23][27] , \REGISTERS[23][26] , \REGISTERS[23][25] ,
         \REGISTERS[23][24] , \REGISTERS[23][23] , \REGISTERS[23][22] ,
         \REGISTERS[23][21] , \REGISTERS[23][20] , \REGISTERS[23][19] ,
         \REGISTERS[23][18] , \REGISTERS[23][17] , \REGISTERS[23][16] ,
         \REGISTERS[23][15] , \REGISTERS[23][14] , \REGISTERS[23][13] ,
         \REGISTERS[23][12] , \REGISTERS[23][11] , \REGISTERS[23][10] ,
         \REGISTERS[23][9] , \REGISTERS[23][8] , \REGISTERS[23][7] ,
         \REGISTERS[23][6] , \REGISTERS[23][5] , \REGISTERS[23][4] ,
         \REGISTERS[23][3] , \REGISTERS[23][2] , \REGISTERS[23][1] ,
         \REGISTERS[23][0] , \REGISTERS[24][31] , \REGISTERS[24][30] ,
         \REGISTERS[24][29] , \REGISTERS[24][28] , \REGISTERS[24][27] ,
         \REGISTERS[24][26] , \REGISTERS[24][25] , \REGISTERS[24][24] ,
         \REGISTERS[24][23] , \REGISTERS[24][22] , \REGISTERS[24][21] ,
         \REGISTERS[24][20] , \REGISTERS[24][19] , \REGISTERS[24][18] ,
         \REGISTERS[24][17] , \REGISTERS[24][16] , \REGISTERS[24][15] ,
         \REGISTERS[24][14] , \REGISTERS[24][13] , \REGISTERS[24][12] ,
         \REGISTERS[24][11] , \REGISTERS[24][10] , \REGISTERS[24][9] ,
         \REGISTERS[24][8] , \REGISTERS[24][7] , \REGISTERS[24][6] ,
         \REGISTERS[24][5] , \REGISTERS[24][4] , \REGISTERS[24][3] ,
         \REGISTERS[24][2] , \REGISTERS[24][1] , \REGISTERS[24][0] ,
         \REGISTERS[25][31] , \REGISTERS[25][30] , \REGISTERS[25][29] ,
         \REGISTERS[25][28] , \REGISTERS[25][27] , \REGISTERS[25][26] ,
         \REGISTERS[25][25] , \REGISTERS[25][24] , \REGISTERS[25][23] ,
         \REGISTERS[25][22] , \REGISTERS[25][21] , \REGISTERS[25][20] ,
         \REGISTERS[25][19] , \REGISTERS[25][18] , \REGISTERS[25][17] ,
         \REGISTERS[25][16] , \REGISTERS[25][15] , \REGISTERS[25][14] ,
         \REGISTERS[25][13] , \REGISTERS[25][12] , \REGISTERS[25][11] ,
         \REGISTERS[25][10] , \REGISTERS[25][9] , \REGISTERS[25][8] ,
         \REGISTERS[25][7] , \REGISTERS[25][6] , \REGISTERS[25][5] ,
         \REGISTERS[25][4] , \REGISTERS[25][3] , \REGISTERS[25][2] ,
         \REGISTERS[25][1] , \REGISTERS[25][0] , \REGISTERS[26][31] ,
         \REGISTERS[26][30] , \REGISTERS[26][29] , \REGISTERS[26][28] ,
         \REGISTERS[26][27] , \REGISTERS[26][26] , \REGISTERS[26][25] ,
         \REGISTERS[26][24] , \REGISTERS[26][23] , \REGISTERS[26][22] ,
         \REGISTERS[26][21] , \REGISTERS[26][20] , \REGISTERS[26][19] ,
         \REGISTERS[26][18] , \REGISTERS[26][17] , \REGISTERS[26][16] ,
         \REGISTERS[26][15] , \REGISTERS[26][14] , \REGISTERS[26][13] ,
         \REGISTERS[26][12] , \REGISTERS[26][11] , \REGISTERS[26][10] ,
         \REGISTERS[26][9] , \REGISTERS[26][8] , \REGISTERS[26][7] ,
         \REGISTERS[26][6] , \REGISTERS[26][5] , \REGISTERS[26][4] ,
         \REGISTERS[26][3] , \REGISTERS[26][2] , \REGISTERS[26][1] ,
         \REGISTERS[26][0] , \REGISTERS[27][31] , \REGISTERS[27][30] ,
         \REGISTERS[27][29] , \REGISTERS[27][28] , \REGISTERS[27][27] ,
         \REGISTERS[27][26] , \REGISTERS[27][25] , \REGISTERS[27][24] ,
         \REGISTERS[27][23] , \REGISTERS[27][22] , \REGISTERS[27][21] ,
         \REGISTERS[27][20] , \REGISTERS[27][19] , \REGISTERS[27][18] ,
         \REGISTERS[27][17] , \REGISTERS[27][16] , \REGISTERS[27][15] ,
         \REGISTERS[27][14] , \REGISTERS[27][13] , \REGISTERS[27][12] ,
         \REGISTERS[27][11] , \REGISTERS[27][10] , \REGISTERS[27][9] ,
         \REGISTERS[27][8] , \REGISTERS[27][7] , \REGISTERS[27][6] ,
         \REGISTERS[27][5] , \REGISTERS[27][4] , \REGISTERS[27][3] ,
         \REGISTERS[27][2] , \REGISTERS[27][1] , \REGISTERS[27][0] ,
         \REGISTERS[28][31] , \REGISTERS[28][30] , \REGISTERS[28][29] ,
         \REGISTERS[28][28] , \REGISTERS[28][27] , \REGISTERS[28][26] ,
         \REGISTERS[28][25] , \REGISTERS[28][24] , \REGISTERS[28][23] ,
         \REGISTERS[28][22] , \REGISTERS[28][21] , \REGISTERS[28][20] ,
         \REGISTERS[28][19] , \REGISTERS[28][18] , \REGISTERS[28][17] ,
         \REGISTERS[28][16] , \REGISTERS[28][15] , \REGISTERS[28][14] ,
         \REGISTERS[28][13] , \REGISTERS[28][12] , \REGISTERS[28][11] ,
         \REGISTERS[28][10] , \REGISTERS[28][9] , \REGISTERS[28][8] ,
         \REGISTERS[28][7] , \REGISTERS[28][6] , \REGISTERS[28][5] ,
         \REGISTERS[28][4] , \REGISTERS[28][3] , \REGISTERS[28][2] ,
         \REGISTERS[28][1] , \REGISTERS[28][0] , \REGISTERS[29][31] ,
         \REGISTERS[29][30] , \REGISTERS[29][29] , \REGISTERS[29][28] ,
         \REGISTERS[29][27] , \REGISTERS[29][26] , \REGISTERS[29][25] ,
         \REGISTERS[29][24] , \REGISTERS[29][23] , \REGISTERS[29][22] ,
         \REGISTERS[29][21] , \REGISTERS[29][20] , \REGISTERS[29][19] ,
         \REGISTERS[29][18] , \REGISTERS[29][17] , \REGISTERS[29][16] ,
         \REGISTERS[29][15] , \REGISTERS[29][14] , \REGISTERS[29][13] ,
         \REGISTERS[29][12] , \REGISTERS[29][11] , \REGISTERS[29][10] ,
         \REGISTERS[29][9] , \REGISTERS[29][8] , \REGISTERS[29][7] ,
         \REGISTERS[29][6] , \REGISTERS[29][5] , \REGISTERS[29][4] ,
         \REGISTERS[29][3] , \REGISTERS[29][2] , \REGISTERS[29][1] ,
         \REGISTERS[29][0] , \REGISTERS[30][31] , \REGISTERS[30][30] ,
         \REGISTERS[30][29] , \REGISTERS[30][28] , \REGISTERS[30][27] ,
         \REGISTERS[30][26] , \REGISTERS[30][25] , \REGISTERS[30][24] ,
         \REGISTERS[30][23] , \REGISTERS[30][22] , \REGISTERS[30][21] ,
         \REGISTERS[30][20] , \REGISTERS[30][19] , \REGISTERS[30][18] ,
         \REGISTERS[30][17] , \REGISTERS[30][16] , \REGISTERS[30][15] ,
         \REGISTERS[30][14] , \REGISTERS[30][13] , \REGISTERS[30][12] ,
         \REGISTERS[30][11] , \REGISTERS[30][10] , \REGISTERS[30][9] ,
         \REGISTERS[30][8] , \REGISTERS[30][7] , \REGISTERS[30][6] ,
         \REGISTERS[30][5] , \REGISTERS[30][4] , \REGISTERS[30][3] ,
         \REGISTERS[30][2] , \REGISTERS[30][1] , \REGISTERS[30][0] ,
         \REGISTERS[31][31] , \REGISTERS[31][30] , \REGISTERS[31][29] ,
         \REGISTERS[31][28] , \REGISTERS[31][27] , \REGISTERS[31][26] ,
         \REGISTERS[31][25] , \REGISTERS[31][24] , \REGISTERS[31][23] ,
         \REGISTERS[31][22] , \REGISTERS[31][21] , \REGISTERS[31][20] ,
         \REGISTERS[31][19] , \REGISTERS[31][18] , \REGISTERS[31][17] ,
         \REGISTERS[31][16] , \REGISTERS[31][15] , \REGISTERS[31][14] ,
         \REGISTERS[31][13] , \REGISTERS[31][12] , \REGISTERS[31][11] ,
         \REGISTERS[31][10] , \REGISTERS[31][9] , \REGISTERS[31][8] ,
         \REGISTERS[31][7] , \REGISTERS[31][6] , \REGISTERS[31][5] ,
         \REGISTERS[31][4] , \REGISTERS[31][3] , \REGISTERS[31][2] ,
         \REGISTERS[31][1] , \REGISTERS[31][0] , N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, n36859, n36860, n36861, n36862, n36863, n36864,
         n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872,
         n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880,
         n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888,
         n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896,
         n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904,
         n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912,
         n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920,
         n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
         n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936,
         n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
         n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952,
         n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960,
         n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968,
         n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976,
         n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984,
         n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992,
         n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
         n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008,
         n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016,
         n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024,
         n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032,
         n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040,
         n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048,
         n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056,
         n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064,
         n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
         n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080,
         n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
         n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096,
         n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104,
         n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112,
         n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120,
         n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128,
         n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136,
         n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
         n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152,
         n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160,
         n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168,
         n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176,
         n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184,
         n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192,
         n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200,
         n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208,
         n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
         n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224,
         n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232,
         n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240,
         n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248,
         n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256,
         n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264,
         n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272,
         n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280,
         n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
         n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296,
         n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
         n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312,
         n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320,
         n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328,
         n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
         n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344,
         n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352,
         n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
         n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368,
         n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
         n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
         n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392,
         n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
         n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408,
         n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416,
         n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424,
         n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
         n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440,
         n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
         n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456,
         n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
         n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472,
         n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480,
         n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488,
         n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496,
         n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
         n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512,
         n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
         n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528,
         n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
         n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544,
         n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552,
         n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560,
         n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
         n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
         n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584,
         n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
         n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
         n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608,
         n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616,
         n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624,
         n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632,
         n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640,
         n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
         n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656,
         n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
         n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
         n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680,
         n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688,
         n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696,
         n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704,
         n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712,
         n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720,
         n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728,
         n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
         n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744,
         n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752,
         n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760,
         n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768,
         n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776,
         n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784,
         n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
         n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
         n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
         n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816,
         n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824,
         n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832,
         n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840,
         n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848,
         n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856,
         n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
         n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872,
         n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880,
         n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888,
         n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896,
         n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904,
         n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912,
         n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920,
         n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928,
         n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936,
         n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944,
         n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
         n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960,
         n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968,
         n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976,
         n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984,
         n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992,
         n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000,
         n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008,
         n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016,
         n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
         n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032,
         n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040,
         n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048,
         n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056,
         n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064,
         n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072,
         n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080,
         n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088,
         n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
         n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104,
         n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112,
         n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120,
         n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128,
         n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136,
         n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144,
         n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
         n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160,
         n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
         n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176,
         n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184,
         n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
         n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
         n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208,
         n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
         n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
         n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232,
         n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
         n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248,
         n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256,
         n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264,
         n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272,
         n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280,
         n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288,
         n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
         n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304,
         n38305;

  DLH_X1 \REGISTERS_reg[1][31]  ( .G(n37757), .D(N275), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(n37757), .D(N274), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(n37757), .D(N273), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(N305), .D(N272), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(n37757), .D(N271), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(N305), .D(N270), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(n37757), .D(N269), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(n37757), .D(N268), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(n37757), .D(N267), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(n37757), .D(N266), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(N305), .D(N265), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n37757), .D(N264), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n37757), .D(N263), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(N305), .D(N262), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(N305), .D(N261), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(n37757), .D(N260), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(N305), .D(N259), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(N305), .D(N258), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(N305), .D(N257), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(N305), .D(N256), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n37757), .D(N255), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(N305), .D(N254), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(N305), .D(N253), .Q(\REGISTERS[1][9] ) );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(N305), .D(N252), .Q(\REGISTERS[1][8] ) );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n37757), .D(N251), .Q(\REGISTERS[1][7] )
         );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(n37757), .D(N250), .Q(\REGISTERS[1][6] )
         );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n37757), .D(N249), .Q(\REGISTERS[1][5] )
         );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(N305), .D(N248), .Q(\REGISTERS[1][4] ) );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(N305), .D(N247), .Q(\REGISTERS[1][3] ) );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(N305), .D(N246), .Q(\REGISTERS[1][2] ) );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(n37757), .D(N245), .Q(\REGISTERS[1][1] )
         );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n37757), .D(N244), .Q(\REGISTERS[1][0] )
         );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(n37758), .D(N275), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(n37758), .D(N274), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(n37758), .D(N273), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(n37758), .D(N272), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(n37758), .D(N271), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(n37758), .D(N270), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(N304), .D(N269), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(N304), .D(N268), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n37758), .D(N267), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n37758), .D(N266), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(n37758), .D(N265), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(n37758), .D(N264), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n37758), .D(N263), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(N304), .D(N262), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n37758), .D(N261), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(N304), .D(N260), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(n37758), .D(N259), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(N304), .D(N258), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(N304), .D(N257), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(N304), .D(N256), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(N304), .D(N255), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n37758), .D(N254), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(N304), .D(N253), .Q(\REGISTERS[2][9] ) );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(N304), .D(N252), .Q(\REGISTERS[2][8] ) );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n37758), .D(N251), .Q(\REGISTERS[2][7] )
         );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(n37758), .D(N250), .Q(\REGISTERS[2][6] )
         );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(N304), .D(N249), .Q(\REGISTERS[2][5] ) );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(N304), .D(N248), .Q(\REGISTERS[2][4] ) );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(N304), .D(N247), .Q(\REGISTERS[2][3] ) );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(N304), .D(N246), .Q(\REGISTERS[2][2] ) );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(n37758), .D(N245), .Q(\REGISTERS[2][1] )
         );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(N304), .D(N244), .Q(\REGISTERS[2][0] ) );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(n37759), .D(N275), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(n37759), .D(N274), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(n37759), .D(N273), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(n37759), .D(N272), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(n37759), .D(N271), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(n37759), .D(N270), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(N303), .D(N269), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(N303), .D(N268), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n37759), .D(N267), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n37759), .D(N266), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(n37759), .D(N265), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(n37759), .D(N264), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n37759), .D(N263), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(N303), .D(N262), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n37759), .D(N261), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(N303), .D(N260), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(n37759), .D(N259), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(N303), .D(N258), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(N303), .D(N257), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(N303), .D(N256), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(N303), .D(N255), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n37759), .D(N254), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(N303), .D(N253), .Q(\REGISTERS[3][9] ) );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(N303), .D(N252), .Q(\REGISTERS[3][8] ) );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n37759), .D(N251), .Q(\REGISTERS[3][7] )
         );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(n37759), .D(N250), .Q(\REGISTERS[3][6] )
         );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(N303), .D(N249), .Q(\REGISTERS[3][5] ) );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(N303), .D(N248), .Q(\REGISTERS[3][4] ) );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(N303), .D(N247), .Q(\REGISTERS[3][3] ) );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(N303), .D(N246), .Q(\REGISTERS[3][2] ) );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(n37759), .D(N245), .Q(\REGISTERS[3][1] )
         );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(N303), .D(N244), .Q(\REGISTERS[3][0] ) );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(n37760), .D(N275), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(n37760), .D(N274), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(n37760), .D(N273), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(n37760), .D(N272), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(n37760), .D(N271), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(n37760), .D(N270), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(N302), .D(N269), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(N302), .D(N268), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n37760), .D(N267), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n37760), .D(N266), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(n37760), .D(N265), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(n37760), .D(N264), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n37760), .D(N263), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(N302), .D(N262), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n37760), .D(N261), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(N302), .D(N260), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(n37760), .D(N259), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(N302), .D(N258), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(N302), .D(N257), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(N302), .D(N256), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(N302), .D(N255), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n37760), .D(N254), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(N302), .D(N253), .Q(\REGISTERS[4][9] ) );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(N302), .D(N252), .Q(\REGISTERS[4][8] ) );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(N302), .D(N251), .Q(\REGISTERS[4][7] ) );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(n37760), .D(N250), .Q(\REGISTERS[4][6] )
         );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(N302), .D(N249), .Q(\REGISTERS[4][5] ) );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(N302), .D(N248), .Q(\REGISTERS[4][4] ) );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(N302), .D(N247), .Q(\REGISTERS[4][3] ) );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(N302), .D(N246), .Q(\REGISTERS[4][2] ) );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(n37760), .D(N245), .Q(\REGISTERS[4][1] )
         );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n37760), .D(N244), .Q(\REGISTERS[4][0] )
         );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(n37761), .D(N275), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(n37761), .D(N274), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(n37761), .D(N273), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(n37761), .D(N272), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(n37761), .D(N271), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(n37761), .D(N270), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(N301), .D(N269), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(N301), .D(N268), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n37761), .D(N267), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n37761), .D(N266), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(n37761), .D(N265), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(n37761), .D(N264), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n37761), .D(N263), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(N301), .D(N262), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n37761), .D(N261), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(N301), .D(N260), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(n37761), .D(N259), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(N301), .D(N258), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(N301), .D(N257), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(N301), .D(N256), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(N301), .D(N255), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n37761), .D(N254), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(N301), .D(N253), .Q(\REGISTERS[5][9] ) );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(N301), .D(N252), .Q(\REGISTERS[5][8] ) );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n37761), .D(N251), .Q(\REGISTERS[5][7] )
         );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(n37761), .D(N250), .Q(\REGISTERS[5][6] )
         );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(N301), .D(N249), .Q(\REGISTERS[5][5] ) );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(N301), .D(N248), .Q(\REGISTERS[5][4] ) );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(N301), .D(N247), .Q(\REGISTERS[5][3] ) );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(N301), .D(N246), .Q(\REGISTERS[5][2] ) );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(n37761), .D(N245), .Q(\REGISTERS[5][1] )
         );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(N301), .D(N244), .Q(\REGISTERS[5][0] ) );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(n37762), .D(N275), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(n37762), .D(N274), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(n37762), .D(N273), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(n37762), .D(N272), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(n37762), .D(N271), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(n37762), .D(N270), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(N300), .D(N269), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(N300), .D(N268), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n37762), .D(N267), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n37762), .D(N266), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(n37762), .D(N265), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(n37762), .D(N264), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n37762), .D(N263), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(N300), .D(N262), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n37762), .D(N261), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(N300), .D(N260), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(n37762), .D(N259), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(N300), .D(N258), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(N300), .D(N257), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(N300), .D(N256), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(N300), .D(N255), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n37762), .D(N254), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(N300), .D(N253), .Q(\REGISTERS[6][9] ) );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(N300), .D(N252), .Q(\REGISTERS[6][8] ) );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(N300), .D(N251), .Q(\REGISTERS[6][7] ) );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(n37762), .D(N250), .Q(\REGISTERS[6][6] )
         );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(N300), .D(N249), .Q(\REGISTERS[6][5] ) );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(N300), .D(N248), .Q(\REGISTERS[6][4] ) );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(N300), .D(N247), .Q(\REGISTERS[6][3] ) );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(N300), .D(N246), .Q(\REGISTERS[6][2] ) );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(n37762), .D(N245), .Q(\REGISTERS[6][1] )
         );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n37762), .D(N244), .Q(\REGISTERS[6][0] )
         );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(n37763), .D(N275), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(n37763), .D(N274), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(n37763), .D(N273), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(n37763), .D(N272), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(n37763), .D(N271), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(n37763), .D(N270), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(N299), .D(N269), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(N299), .D(N268), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n37763), .D(N267), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n37763), .D(N266), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(n37763), .D(N265), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(n37763), .D(N264), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n37763), .D(N263), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(N299), .D(N262), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n37763), .D(N261), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(N299), .D(N260), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(n37763), .D(N259), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(N299), .D(N258), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(N299), .D(N257), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(N299), .D(N256), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(N299), .D(N255), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n37763), .D(N254), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(N299), .D(N253), .Q(\REGISTERS[7][9] ) );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(N299), .D(N252), .Q(\REGISTERS[7][8] ) );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n37763), .D(N251), .Q(\REGISTERS[7][7] )
         );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(n37763), .D(N250), .Q(\REGISTERS[7][6] )
         );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(N299), .D(N249), .Q(\REGISTERS[7][5] ) );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(N299), .D(N248), .Q(\REGISTERS[7][4] ) );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(N299), .D(N247), .Q(\REGISTERS[7][3] ) );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(N299), .D(N246), .Q(\REGISTERS[7][2] ) );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(n37763), .D(N245), .Q(\REGISTERS[7][1] )
         );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(N299), .D(N244), .Q(\REGISTERS[7][0] ) );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(n37764), .D(N275), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(n37764), .D(N274), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(n37764), .D(N273), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(n37764), .D(N272), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(n37764), .D(N271), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(n37764), .D(N270), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(N298), .D(N269), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(N298), .D(N268), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n37764), .D(N267), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n37764), .D(N266), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(n37764), .D(N265), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(n37764), .D(N264), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n37764), .D(N263), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(N298), .D(N262), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n37764), .D(N261), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(N298), .D(N260), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(n37764), .D(N259), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(N298), .D(N258), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(N298), .D(N257), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(N298), .D(N256), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(N298), .D(N255), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n37764), .D(N254), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(N298), .D(N253), .Q(\REGISTERS[8][9] ) );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(N298), .D(N252), .Q(\REGISTERS[8][8] ) );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n37764), .D(N251), .Q(\REGISTERS[8][7] )
         );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(n37764), .D(N250), .Q(\REGISTERS[8][6] )
         );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(N298), .D(N249), .Q(\REGISTERS[8][5] ) );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(N298), .D(N248), .Q(\REGISTERS[8][4] ) );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(N298), .D(N247), .Q(\REGISTERS[8][3] ) );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(N298), .D(N246), .Q(\REGISTERS[8][2] ) );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(n37764), .D(N245), .Q(\REGISTERS[8][1] )
         );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(N298), .D(N244), .Q(\REGISTERS[8][0] ) );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(n37765), .D(N275), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(n37765), .D(N274), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(n37765), .D(N273), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(n37765), .D(N272), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(n37765), .D(N271), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(n37765), .D(N270), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(N297), .D(N269), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(N297), .D(N268), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n37765), .D(N267), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n37765), .D(N266), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(n37765), .D(N265), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(n37765), .D(N264), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n37765), .D(N263), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(N297), .D(N262), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n37765), .D(N261), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(N297), .D(N260), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(n37765), .D(N259), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(N297), .D(N258), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(N297), .D(N257), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(N297), .D(N256), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(N297), .D(N255), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n37765), .D(N254), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(N297), .D(N253), .Q(\REGISTERS[9][9] ) );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(N297), .D(N252), .Q(\REGISTERS[9][8] ) );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n37765), .D(N251), .Q(\REGISTERS[9][7] )
         );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(n37765), .D(N250), .Q(\REGISTERS[9][6] )
         );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(N297), .D(N249), .Q(\REGISTERS[9][5] ) );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(N297), .D(N248), .Q(\REGISTERS[9][4] ) );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(N297), .D(N247), .Q(\REGISTERS[9][3] ) );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(N297), .D(N246), .Q(\REGISTERS[9][2] ) );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(n37765), .D(N245), .Q(\REGISTERS[9][1] )
         );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(N297), .D(N244), .Q(\REGISTERS[9][0] ) );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(n37766), .D(N275), .Q(
        \REGISTERS[10][31] ) );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(n37766), .D(N274), .Q(
        \REGISTERS[10][30] ) );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(n37766), .D(N273), .Q(
        \REGISTERS[10][29] ) );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(n37766), .D(N272), .Q(
        \REGISTERS[10][28] ) );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(n37766), .D(N271), .Q(
        \REGISTERS[10][27] ) );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(n37766), .D(N270), .Q(
        \REGISTERS[10][26] ) );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(N296), .D(N269), .Q(\REGISTERS[10][25] )
         );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(N296), .D(N268), .Q(\REGISTERS[10][24] )
         );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n37766), .D(N267), .Q(
        \REGISTERS[10][23] ) );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(N296), .D(N266), .Q(\REGISTERS[10][22] )
         );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(n37766), .D(N265), .Q(
        \REGISTERS[10][21] ) );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(n37766), .D(N264), .Q(
        \REGISTERS[10][20] ) );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n37766), .D(N263), .Q(
        \REGISTERS[10][19] ) );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(N296), .D(N262), .Q(\REGISTERS[10][18] )
         );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(N296), .D(N261), .Q(\REGISTERS[10][17] )
         );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n37766), .D(N260), .Q(
        \REGISTERS[10][16] ) );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(N296), .D(N259), .Q(\REGISTERS[10][15] )
         );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(n37766), .D(N258), .Q(
        \REGISTERS[10][14] ) );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n37766), .D(N257), .Q(
        \REGISTERS[10][13] ) );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(N296), .D(N256), .Q(\REGISTERS[10][12] )
         );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n37766), .D(N255), .Q(
        \REGISTERS[10][11] ) );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n37766), .D(N254), .Q(
        \REGISTERS[10][10] ) );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(N296), .D(N253), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(N296), .D(N252), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(N296), .D(N251), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(n37766), .D(N250), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(N296), .D(N249), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(N296), .D(N248), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(N296), .D(N247), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(N296), .D(N246), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(n37766), .D(N245), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(N296), .D(N244), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(n37767), .D(N275), .Q(
        \REGISTERS[11][31] ) );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(n37767), .D(N274), .Q(
        \REGISTERS[11][30] ) );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(n37767), .D(N273), .Q(
        \REGISTERS[11][29] ) );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(n37767), .D(N272), .Q(
        \REGISTERS[11][28] ) );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(n37767), .D(N271), .Q(
        \REGISTERS[11][27] ) );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(n37767), .D(N270), .Q(
        \REGISTERS[11][26] ) );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(N295), .D(N269), .Q(\REGISTERS[11][25] )
         );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(N295), .D(N268), .Q(\REGISTERS[11][24] )
         );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n37767), .D(N267), .Q(
        \REGISTERS[11][23] ) );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n37767), .D(N266), .Q(
        \REGISTERS[11][22] ) );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(n37767), .D(N265), .Q(
        \REGISTERS[11][21] ) );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(n37767), .D(N264), .Q(
        \REGISTERS[11][20] ) );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n37767), .D(N263), .Q(
        \REGISTERS[11][19] ) );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(N295), .D(N262), .Q(\REGISTERS[11][18] )
         );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n37767), .D(N261), .Q(
        \REGISTERS[11][17] ) );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(N295), .D(N260), .Q(\REGISTERS[11][16] )
         );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(n37767), .D(N259), .Q(
        \REGISTERS[11][15] ) );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(N295), .D(N258), .Q(\REGISTERS[11][14] )
         );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(N295), .D(N257), .Q(\REGISTERS[11][13] )
         );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(N295), .D(N256), .Q(\REGISTERS[11][12] )
         );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(N295), .D(N255), .Q(\REGISTERS[11][11] )
         );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n37767), .D(N254), .Q(
        \REGISTERS[11][10] ) );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(N295), .D(N253), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(N295), .D(N252), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n37767), .D(N251), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(n37767), .D(N250), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(N295), .D(N249), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(N295), .D(N248), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(N295), .D(N247), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(N295), .D(N246), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(n37767), .D(N245), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(N295), .D(N244), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(n37768), .D(N275), .Q(
        \REGISTERS[12][31] ) );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(n37768), .D(N274), .Q(
        \REGISTERS[12][30] ) );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(n37768), .D(N273), .Q(
        \REGISTERS[12][29] ) );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(n37768), .D(N272), .Q(
        \REGISTERS[12][28] ) );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(n37768), .D(N271), .Q(
        \REGISTERS[12][27] ) );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(n37768), .D(N270), .Q(
        \REGISTERS[12][26] ) );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(N294), .D(N269), .Q(\REGISTERS[12][25] )
         );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(N294), .D(N268), .Q(\REGISTERS[12][24] )
         );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n37768), .D(N267), .Q(
        \REGISTERS[12][23] ) );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n37768), .D(N266), .Q(
        \REGISTERS[12][22] ) );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(n37768), .D(N265), .Q(
        \REGISTERS[12][21] ) );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(n37768), .D(N264), .Q(
        \REGISTERS[12][20] ) );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n37768), .D(N263), .Q(
        \REGISTERS[12][19] ) );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(N294), .D(N262), .Q(\REGISTERS[12][18] )
         );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n37768), .D(N261), .Q(
        \REGISTERS[12][17] ) );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(N294), .D(N260), .Q(\REGISTERS[12][16] )
         );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(n37768), .D(N259), .Q(
        \REGISTERS[12][15] ) );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(N294), .D(N258), .Q(\REGISTERS[12][14] )
         );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(N294), .D(N257), .Q(\REGISTERS[12][13] )
         );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(N294), .D(N256), .Q(\REGISTERS[12][12] )
         );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n37768), .D(N255), .Q(
        \REGISTERS[12][11] ) );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n37768), .D(N254), .Q(
        \REGISTERS[12][10] ) );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(N294), .D(N253), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(N294), .D(N252), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(N294), .D(N251), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(n37768), .D(N250), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(N294), .D(N249), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(N294), .D(N248), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(N294), .D(N247), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(N294), .D(N246), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(n37768), .D(N245), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(N294), .D(N244), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(n37769), .D(N275), .Q(
        \REGISTERS[13][31] ) );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(n37769), .D(N274), .Q(
        \REGISTERS[13][30] ) );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(n37769), .D(N273), .Q(
        \REGISTERS[13][29] ) );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(n37769), .D(N272), .Q(
        \REGISTERS[13][28] ) );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(n37769), .D(N271), .Q(
        \REGISTERS[13][27] ) );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(n37769), .D(N270), .Q(
        \REGISTERS[13][26] ) );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(N293), .D(N269), .Q(\REGISTERS[13][25] )
         );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(N293), .D(N268), .Q(\REGISTERS[13][24] )
         );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n37769), .D(N267), .Q(
        \REGISTERS[13][23] ) );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n37769), .D(N266), .Q(
        \REGISTERS[13][22] ) );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(n37769), .D(N265), .Q(
        \REGISTERS[13][21] ) );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(n37769), .D(N264), .Q(
        \REGISTERS[13][20] ) );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n37769), .D(N263), .Q(
        \REGISTERS[13][19] ) );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(N293), .D(N262), .Q(\REGISTERS[13][18] )
         );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n37769), .D(N261), .Q(
        \REGISTERS[13][17] ) );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(N293), .D(N260), .Q(\REGISTERS[13][16] )
         );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(n37769), .D(N259), .Q(
        \REGISTERS[13][15] ) );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(N293), .D(N258), .Q(\REGISTERS[13][14] )
         );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(N293), .D(N257), .Q(\REGISTERS[13][13] )
         );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(N293), .D(N256), .Q(\REGISTERS[13][12] )
         );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(N293), .D(N255), .Q(\REGISTERS[13][11] )
         );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n37769), .D(N254), .Q(
        \REGISTERS[13][10] ) );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(N293), .D(N253), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(N293), .D(N252), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n37769), .D(N251), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(n37769), .D(N250), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(N293), .D(N249), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(N293), .D(N248), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(N293), .D(N247), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(N293), .D(N246), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(n37769), .D(N245), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(N293), .D(N244), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(n37770), .D(N275), .Q(
        \REGISTERS[14][31] ) );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(n37770), .D(N274), .Q(
        \REGISTERS[14][30] ) );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(n37770), .D(N273), .Q(
        \REGISTERS[14][29] ) );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(n37770), .D(N272), .Q(
        \REGISTERS[14][28] ) );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(n37770), .D(N271), .Q(
        \REGISTERS[14][27] ) );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(n37770), .D(N270), .Q(
        \REGISTERS[14][26] ) );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(N292), .D(N269), .Q(\REGISTERS[14][25] )
         );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(N292), .D(N268), .Q(\REGISTERS[14][24] )
         );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n37770), .D(N267), .Q(
        \REGISTERS[14][23] ) );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n37770), .D(N266), .Q(
        \REGISTERS[14][22] ) );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(n37770), .D(N265), .Q(
        \REGISTERS[14][21] ) );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(n37770), .D(N264), .Q(
        \REGISTERS[14][20] ) );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n37770), .D(N263), .Q(
        \REGISTERS[14][19] ) );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(N292), .D(N262), .Q(\REGISTERS[14][18] )
         );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n37770), .D(N261), .Q(
        \REGISTERS[14][17] ) );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(N292), .D(N260), .Q(\REGISTERS[14][16] )
         );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(n37770), .D(N259), .Q(
        \REGISTERS[14][15] ) );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(N292), .D(N258), .Q(\REGISTERS[14][14] )
         );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(N292), .D(N257), .Q(\REGISTERS[14][13] )
         );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(N292), .D(N256), .Q(\REGISTERS[14][12] )
         );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(N292), .D(N255), .Q(\REGISTERS[14][11] )
         );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n37770), .D(N254), .Q(
        \REGISTERS[14][10] ) );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(N292), .D(N253), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(N292), .D(N252), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n37770), .D(N251), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(n37770), .D(N250), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(N292), .D(N249), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(N292), .D(N248), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(N292), .D(N247), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(N292), .D(N246), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(n37770), .D(N245), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(N292), .D(N244), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(n37771), .D(N275), .Q(
        \REGISTERS[15][31] ) );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(n37771), .D(N274), .Q(
        \REGISTERS[15][30] ) );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(n37771), .D(N273), .Q(
        \REGISTERS[15][29] ) );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(n37771), .D(N272), .Q(
        \REGISTERS[15][28] ) );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(n37771), .D(N271), .Q(
        \REGISTERS[15][27] ) );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(n37771), .D(N270), .Q(
        \REGISTERS[15][26] ) );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(N291), .D(N269), .Q(\REGISTERS[15][25] )
         );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(N291), .D(N268), .Q(\REGISTERS[15][24] )
         );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n37771), .D(N267), .Q(
        \REGISTERS[15][23] ) );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n37771), .D(N266), .Q(
        \REGISTERS[15][22] ) );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(n37771), .D(N265), .Q(
        \REGISTERS[15][21] ) );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(n37771), .D(N264), .Q(
        \REGISTERS[15][20] ) );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n37771), .D(N263), .Q(
        \REGISTERS[15][19] ) );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(N291), .D(N262), .Q(\REGISTERS[15][18] )
         );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n37771), .D(N261), .Q(
        \REGISTERS[15][17] ) );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(N291), .D(N260), .Q(\REGISTERS[15][16] )
         );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(n37771), .D(N259), .Q(
        \REGISTERS[15][15] ) );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(N291), .D(N258), .Q(\REGISTERS[15][14] )
         );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(N291), .D(N257), .Q(\REGISTERS[15][13] )
         );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(N291), .D(N256), .Q(\REGISTERS[15][12] )
         );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(N291), .D(N255), .Q(\REGISTERS[15][11] )
         );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n37771), .D(N254), .Q(
        \REGISTERS[15][10] ) );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(N291), .D(N253), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(N291), .D(N252), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n37771), .D(N251), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(n37771), .D(N250), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(N291), .D(N249), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(N291), .D(N248), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(N291), .D(N247), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(N291), .D(N246), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(n37771), .D(N245), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(N291), .D(N244), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(n37772), .D(N275), .Q(
        \REGISTERS[16][31] ) );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(n37772), .D(N274), .Q(
        \REGISTERS[16][30] ) );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(n37772), .D(N273), .Q(
        \REGISTERS[16][29] ) );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(n37772), .D(N272), .Q(
        \REGISTERS[16][28] ) );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(n37772), .D(N271), .Q(
        \REGISTERS[16][27] ) );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(n37772), .D(N270), .Q(
        \REGISTERS[16][26] ) );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(N290), .D(N269), .Q(\REGISTERS[16][25] )
         );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(N290), .D(N268), .Q(\REGISTERS[16][24] )
         );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n37772), .D(N267), .Q(
        \REGISTERS[16][23] ) );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n37772), .D(N266), .Q(
        \REGISTERS[16][22] ) );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(n37772), .D(N265), .Q(
        \REGISTERS[16][21] ) );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(n37772), .D(N264), .Q(
        \REGISTERS[16][20] ) );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n37772), .D(N263), .Q(
        \REGISTERS[16][19] ) );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(N290), .D(N262), .Q(\REGISTERS[16][18] )
         );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n37772), .D(N261), .Q(
        \REGISTERS[16][17] ) );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(N290), .D(N260), .Q(\REGISTERS[16][16] )
         );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(n37772), .D(N259), .Q(
        \REGISTERS[16][15] ) );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(N290), .D(N258), .Q(\REGISTERS[16][14] )
         );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(N290), .D(N257), .Q(\REGISTERS[16][13] )
         );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(N290), .D(N256), .Q(\REGISTERS[16][12] )
         );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(N290), .D(N255), .Q(\REGISTERS[16][11] )
         );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n37772), .D(N254), .Q(
        \REGISTERS[16][10] ) );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(N290), .D(N253), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(N290), .D(N252), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n37772), .D(N251), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(n37772), .D(N250), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(N290), .D(N249), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(N290), .D(N248), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(N290), .D(N247), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(N290), .D(N246), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(n37772), .D(N245), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(N290), .D(N244), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(n37773), .D(N275), .Q(
        \REGISTERS[17][31] ) );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(n37773), .D(N274), .Q(
        \REGISTERS[17][30] ) );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(n37773), .D(N273), .Q(
        \REGISTERS[17][29] ) );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(n37773), .D(N272), .Q(
        \REGISTERS[17][28] ) );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(n37773), .D(N271), .Q(
        \REGISTERS[17][27] ) );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(n37773), .D(N270), .Q(
        \REGISTERS[17][26] ) );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(N289), .D(N269), .Q(\REGISTERS[17][25] )
         );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(N289), .D(N268), .Q(\REGISTERS[17][24] )
         );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n37773), .D(N267), .Q(
        \REGISTERS[17][23] ) );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n37773), .D(N266), .Q(
        \REGISTERS[17][22] ) );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(n37773), .D(N265), .Q(
        \REGISTERS[17][21] ) );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(n37773), .D(N264), .Q(
        \REGISTERS[17][20] ) );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n37773), .D(N263), .Q(
        \REGISTERS[17][19] ) );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(N289), .D(N262), .Q(\REGISTERS[17][18] )
         );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n37773), .D(N261), .Q(
        \REGISTERS[17][17] ) );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(N289), .D(N260), .Q(\REGISTERS[17][16] )
         );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(n37773), .D(N259), .Q(
        \REGISTERS[17][15] ) );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(N289), .D(N258), .Q(\REGISTERS[17][14] )
         );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(N289), .D(N257), .Q(\REGISTERS[17][13] )
         );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(N289), .D(N256), .Q(\REGISTERS[17][12] )
         );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(N289), .D(N255), .Q(\REGISTERS[17][11] )
         );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n37773), .D(N254), .Q(
        \REGISTERS[17][10] ) );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(N289), .D(N253), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(N289), .D(N252), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n37773), .D(N251), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(n37773), .D(N250), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(N289), .D(N249), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(N289), .D(N248), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(N289), .D(N247), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(N289), .D(N246), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(n37773), .D(N245), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(N289), .D(N244), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(n37774), .D(N275), .Q(
        \REGISTERS[18][31] ) );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(n37774), .D(N274), .Q(
        \REGISTERS[18][30] ) );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(n37774), .D(N273), .Q(
        \REGISTERS[18][29] ) );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(n37774), .D(N272), .Q(
        \REGISTERS[18][28] ) );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(n37774), .D(N271), .Q(
        \REGISTERS[18][27] ) );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(n37774), .D(N270), .Q(
        \REGISTERS[18][26] ) );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(N288), .D(N269), .Q(\REGISTERS[18][25] )
         );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(N288), .D(N268), .Q(\REGISTERS[18][24] )
         );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n37774), .D(N267), .Q(
        \REGISTERS[18][23] ) );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n37774), .D(N266), .Q(
        \REGISTERS[18][22] ) );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(n37774), .D(N265), .Q(
        \REGISTERS[18][21] ) );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(n37774), .D(N264), .Q(
        \REGISTERS[18][20] ) );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n37774), .D(N263), .Q(
        \REGISTERS[18][19] ) );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(N288), .D(N262), .Q(\REGISTERS[18][18] )
         );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n37774), .D(N261), .Q(
        \REGISTERS[18][17] ) );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(N288), .D(N260), .Q(\REGISTERS[18][16] )
         );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(n37774), .D(N259), .Q(
        \REGISTERS[18][15] ) );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(N288), .D(N258), .Q(\REGISTERS[18][14] )
         );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(N288), .D(N257), .Q(\REGISTERS[18][13] )
         );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(N288), .D(N256), .Q(\REGISTERS[18][12] )
         );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(N288), .D(N255), .Q(\REGISTERS[18][11] )
         );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n37774), .D(N254), .Q(
        \REGISTERS[18][10] ) );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(N288), .D(N253), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(N288), .D(N252), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n37774), .D(N251), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(n37774), .D(N250), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(N288), .D(N249), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(N288), .D(N248), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(N288), .D(N247), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(N288), .D(N246), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(n37774), .D(N245), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(N288), .D(N244), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(n37775), .D(N275), .Q(
        \REGISTERS[19][31] ) );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(n37775), .D(N274), .Q(
        \REGISTERS[19][30] ) );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(n37775), .D(N273), .Q(
        \REGISTERS[19][29] ) );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(n37775), .D(N272), .Q(
        \REGISTERS[19][28] ) );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(n37775), .D(N271), .Q(
        \REGISTERS[19][27] ) );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(n37775), .D(N270), .Q(
        \REGISTERS[19][26] ) );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(N287), .D(N269), .Q(\REGISTERS[19][25] )
         );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(N287), .D(N268), .Q(\REGISTERS[19][24] )
         );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n37775), .D(N267), .Q(
        \REGISTERS[19][23] ) );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n37775), .D(N266), .Q(
        \REGISTERS[19][22] ) );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(n37775), .D(N265), .Q(
        \REGISTERS[19][21] ) );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(n37775), .D(N264), .Q(
        \REGISTERS[19][20] ) );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n37775), .D(N263), .Q(
        \REGISTERS[19][19] ) );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(N287), .D(N262), .Q(\REGISTERS[19][18] )
         );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n37775), .D(N261), .Q(
        \REGISTERS[19][17] ) );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(N287), .D(N260), .Q(\REGISTERS[19][16] )
         );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(n37775), .D(N259), .Q(
        \REGISTERS[19][15] ) );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(N287), .D(N258), .Q(\REGISTERS[19][14] )
         );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(N287), .D(N257), .Q(\REGISTERS[19][13] )
         );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(N287), .D(N256), .Q(\REGISTERS[19][12] )
         );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(N287), .D(N255), .Q(\REGISTERS[19][11] )
         );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n37775), .D(N254), .Q(
        \REGISTERS[19][10] ) );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(N287), .D(N253), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(N287), .D(N252), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n37775), .D(N251), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(n37775), .D(N250), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(N287), .D(N249), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(N287), .D(N248), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(N287), .D(N247), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(N287), .D(N246), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(n37775), .D(N245), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(N287), .D(N244), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(n37776), .D(N275), .Q(
        \REGISTERS[20][31] ) );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(n37776), .D(N274), .Q(
        \REGISTERS[20][30] ) );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(n37776), .D(N273), .Q(
        \REGISTERS[20][29] ) );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(n37776), .D(N272), .Q(
        \REGISTERS[20][28] ) );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(n37776), .D(N271), .Q(
        \REGISTERS[20][27] ) );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(n37776), .D(N270), .Q(
        \REGISTERS[20][26] ) );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(N286), .D(N269), .Q(\REGISTERS[20][25] )
         );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(N286), .D(N268), .Q(\REGISTERS[20][24] )
         );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n37776), .D(N267), .Q(
        \REGISTERS[20][23] ) );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n37776), .D(N266), .Q(
        \REGISTERS[20][22] ) );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(n37776), .D(N265), .Q(
        \REGISTERS[20][21] ) );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(n37776), .D(N264), .Q(
        \REGISTERS[20][20] ) );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n37776), .D(N263), .Q(
        \REGISTERS[20][19] ) );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(N286), .D(N262), .Q(\REGISTERS[20][18] )
         );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n37776), .D(N261), .Q(
        \REGISTERS[20][17] ) );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(N286), .D(N260), .Q(\REGISTERS[20][16] )
         );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(n37776), .D(N259), .Q(
        \REGISTERS[20][15] ) );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(N286), .D(N258), .Q(\REGISTERS[20][14] )
         );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(N286), .D(N257), .Q(\REGISTERS[20][13] )
         );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(N286), .D(N256), .Q(\REGISTERS[20][12] )
         );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(N286), .D(N255), .Q(\REGISTERS[20][11] )
         );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n37776), .D(N254), .Q(
        \REGISTERS[20][10] ) );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(N286), .D(N253), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(N286), .D(N252), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n37776), .D(N251), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(n37776), .D(N250), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(N286), .D(N249), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(N286), .D(N248), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(N286), .D(N247), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(N286), .D(N246), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(n37776), .D(N245), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(N286), .D(N244), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(n37777), .D(N275), .Q(
        \REGISTERS[21][31] ) );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(n37777), .D(N274), .Q(
        \REGISTERS[21][30] ) );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(n37777), .D(N273), .Q(
        \REGISTERS[21][29] ) );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(n37777), .D(N272), .Q(
        \REGISTERS[21][28] ) );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(n37777), .D(N271), .Q(
        \REGISTERS[21][27] ) );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(n37777), .D(N270), .Q(
        \REGISTERS[21][26] ) );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(N285), .D(N269), .Q(\REGISTERS[21][25] )
         );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(N285), .D(N268), .Q(\REGISTERS[21][24] )
         );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n37777), .D(N267), .Q(
        \REGISTERS[21][23] ) );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n37777), .D(N266), .Q(
        \REGISTERS[21][22] ) );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(n37777), .D(N265), .Q(
        \REGISTERS[21][21] ) );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(n37777), .D(N264), .Q(
        \REGISTERS[21][20] ) );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n37777), .D(N263), .Q(
        \REGISTERS[21][19] ) );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(N285), .D(N262), .Q(\REGISTERS[21][18] )
         );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n37777), .D(N261), .Q(
        \REGISTERS[21][17] ) );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(N285), .D(N260), .Q(\REGISTERS[21][16] )
         );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(n37777), .D(N259), .Q(
        \REGISTERS[21][15] ) );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(N285), .D(N258), .Q(\REGISTERS[21][14] )
         );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(N285), .D(N257), .Q(\REGISTERS[21][13] )
         );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(N285), .D(N256), .Q(\REGISTERS[21][12] )
         );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(N285), .D(N255), .Q(\REGISTERS[21][11] )
         );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n37777), .D(N254), .Q(
        \REGISTERS[21][10] ) );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(N285), .D(N253), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(N285), .D(N252), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n37777), .D(N251), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(n37777), .D(N250), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(N285), .D(N249), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(N285), .D(N248), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(N285), .D(N247), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(N285), .D(N246), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(n37777), .D(N245), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(N285), .D(N244), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(n37778), .D(N275), .Q(
        \REGISTERS[22][31] ) );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(n37778), .D(N274), .Q(
        \REGISTERS[22][30] ) );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(n37778), .D(N273), .Q(
        \REGISTERS[22][29] ) );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(n37778), .D(N272), .Q(
        \REGISTERS[22][28] ) );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(n37778), .D(N271), .Q(
        \REGISTERS[22][27] ) );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(n37778), .D(N270), .Q(
        \REGISTERS[22][26] ) );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(N284), .D(N269), .Q(\REGISTERS[22][25] )
         );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(N284), .D(N268), .Q(\REGISTERS[22][24] )
         );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n37778), .D(N267), .Q(
        \REGISTERS[22][23] ) );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n37778), .D(N266), .Q(
        \REGISTERS[22][22] ) );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(n37778), .D(N265), .Q(
        \REGISTERS[22][21] ) );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(n37778), .D(N264), .Q(
        \REGISTERS[22][20] ) );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n37778), .D(N263), .Q(
        \REGISTERS[22][19] ) );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(N284), .D(N262), .Q(\REGISTERS[22][18] )
         );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n37778), .D(N261), .Q(
        \REGISTERS[22][17] ) );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(N284), .D(N260), .Q(\REGISTERS[22][16] )
         );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(n37778), .D(N259), .Q(
        \REGISTERS[22][15] ) );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(N284), .D(N258), .Q(\REGISTERS[22][14] )
         );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(N284), .D(N257), .Q(\REGISTERS[22][13] )
         );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(N284), .D(N256), .Q(\REGISTERS[22][12] )
         );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(N284), .D(N255), .Q(\REGISTERS[22][11] )
         );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n37778), .D(N254), .Q(
        \REGISTERS[22][10] ) );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(N284), .D(N253), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(N284), .D(N252), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n37778), .D(N251), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(n37778), .D(N250), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(N284), .D(N249), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(N284), .D(N248), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(N284), .D(N247), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(N284), .D(N246), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(n37778), .D(N245), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(N284), .D(N244), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(n37779), .D(N275), .Q(
        \REGISTERS[23][31] ) );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(n37779), .D(N274), .Q(
        \REGISTERS[23][30] ) );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(n37779), .D(N273), .Q(
        \REGISTERS[23][29] ) );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(n37779), .D(N272), .Q(
        \REGISTERS[23][28] ) );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(n37779), .D(N271), .Q(
        \REGISTERS[23][27] ) );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(n37779), .D(N270), .Q(
        \REGISTERS[23][26] ) );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(N283), .D(N269), .Q(\REGISTERS[23][25] )
         );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(N283), .D(N268), .Q(\REGISTERS[23][24] )
         );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n37779), .D(N267), .Q(
        \REGISTERS[23][23] ) );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n37779), .D(N266), .Q(
        \REGISTERS[23][22] ) );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(n37779), .D(N265), .Q(
        \REGISTERS[23][21] ) );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(n37779), .D(N264), .Q(
        \REGISTERS[23][20] ) );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n37779), .D(N263), .Q(
        \REGISTERS[23][19] ) );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(N283), .D(N262), .Q(\REGISTERS[23][18] )
         );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n37779), .D(N261), .Q(
        \REGISTERS[23][17] ) );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(N283), .D(N260), .Q(\REGISTERS[23][16] )
         );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(n37779), .D(N259), .Q(
        \REGISTERS[23][15] ) );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(N283), .D(N258), .Q(\REGISTERS[23][14] )
         );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(N283), .D(N257), .Q(\REGISTERS[23][13] )
         );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(N283), .D(N256), .Q(\REGISTERS[23][12] )
         );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(N283), .D(N255), .Q(\REGISTERS[23][11] )
         );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n37779), .D(N254), .Q(
        \REGISTERS[23][10] ) );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(N283), .D(N253), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(N283), .D(N252), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n37779), .D(N251), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(n37779), .D(N250), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(N283), .D(N249), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(N283), .D(N248), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(N283), .D(N247), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(N283), .D(N246), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(n37779), .D(N245), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(N283), .D(N244), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(n37780), .D(N275), .Q(
        \REGISTERS[24][31] ) );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(n37780), .D(N274), .Q(
        \REGISTERS[24][30] ) );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(n37780), .D(N273), .Q(
        \REGISTERS[24][29] ) );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(n37780), .D(N272), .Q(
        \REGISTERS[24][28] ) );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(n37780), .D(N271), .Q(
        \REGISTERS[24][27] ) );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(n37780), .D(N270), .Q(
        \REGISTERS[24][26] ) );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(n37780), .D(N269), .Q(
        \REGISTERS[24][25] ) );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n37780), .D(N268), .Q(
        \REGISTERS[24][24] ) );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n37780), .D(N267), .Q(
        \REGISTERS[24][23] ) );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(N282), .D(N266), .Q(\REGISTERS[24][22] )
         );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n37780), .D(N265), .Q(
        \REGISTERS[24][21] ) );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n37780), .D(N264), .Q(
        \REGISTERS[24][20] ) );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(n37780), .D(N263), .Q(
        \REGISTERS[24][19] ) );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(N282), .D(N262), .Q(\REGISTERS[24][18] )
         );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(N282), .D(N261), .Q(\REGISTERS[24][17] )
         );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(N282), .D(N260), .Q(\REGISTERS[24][16] )
         );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n37780), .D(N259), .Q(
        \REGISTERS[24][15] ) );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(N282), .D(N258), .Q(\REGISTERS[24][14] )
         );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(N282), .D(N257), .Q(\REGISTERS[24][13] )
         );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(N282), .D(N256), .Q(\REGISTERS[24][12] )
         );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(n37780), .D(N255), .Q(
        \REGISTERS[24][11] ) );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(n37780), .D(N254), .Q(
        \REGISTERS[24][10] ) );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(N282), .D(N253), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(N282), .D(N252), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(n37780), .D(N251), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n37780), .D(N250), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(N282), .D(N249), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(N282), .D(N248), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(N282), .D(N247), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(N282), .D(N246), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(N282), .D(N245), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(N282), .D(N244), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(n37781), .D(N275), .Q(
        \REGISTERS[25][31] ) );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(n37781), .D(N274), .Q(
        \REGISTERS[25][30] ) );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(n37781), .D(N273), .Q(
        \REGISTERS[25][29] ) );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(n37781), .D(N272), .Q(
        \REGISTERS[25][28] ) );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(n37781), .D(N271), .Q(
        \REGISTERS[25][27] ) );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(n37781), .D(N270), .Q(
        \REGISTERS[25][26] ) );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(N281), .D(N269), .Q(\REGISTERS[25][25] )
         );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(N281), .D(N268), .Q(\REGISTERS[25][24] )
         );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n37781), .D(N267), .Q(
        \REGISTERS[25][23] ) );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n37781), .D(N266), .Q(
        \REGISTERS[25][22] ) );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(n37781), .D(N265), .Q(
        \REGISTERS[25][21] ) );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(n37781), .D(N264), .Q(
        \REGISTERS[25][20] ) );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n37781), .D(N263), .Q(
        \REGISTERS[25][19] ) );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(N281), .D(N262), .Q(\REGISTERS[25][18] )
         );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n37781), .D(N261), .Q(
        \REGISTERS[25][17] ) );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(N281), .D(N260), .Q(\REGISTERS[25][16] )
         );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(n37781), .D(N259), .Q(
        \REGISTERS[25][15] ) );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(N281), .D(N258), .Q(\REGISTERS[25][14] )
         );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(N281), .D(N257), .Q(\REGISTERS[25][13] )
         );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(N281), .D(N256), .Q(\REGISTERS[25][12] )
         );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(N281), .D(N255), .Q(\REGISTERS[25][11] )
         );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n37781), .D(N254), .Q(
        \REGISTERS[25][10] ) );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(N281), .D(N253), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(N281), .D(N252), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n37781), .D(N251), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(n37781), .D(N250), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(N281), .D(N249), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(N281), .D(N248), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(N281), .D(N247), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(N281), .D(N246), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(n37781), .D(N245), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(N281), .D(N244), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(n37782), .D(N275), .Q(
        \REGISTERS[26][31] ) );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(n37782), .D(N274), .Q(
        \REGISTERS[26][30] ) );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(n37782), .D(N273), .Q(
        \REGISTERS[26][29] ) );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(n37782), .D(N272), .Q(
        \REGISTERS[26][28] ) );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(n37782), .D(N271), .Q(
        \REGISTERS[26][27] ) );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(n37782), .D(N270), .Q(
        \REGISTERS[26][26] ) );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(N280), .D(N269), .Q(\REGISTERS[26][25] )
         );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(N280), .D(N268), .Q(\REGISTERS[26][24] )
         );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n37782), .D(N267), .Q(
        \REGISTERS[26][23] ) );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n37782), .D(N266), .Q(
        \REGISTERS[26][22] ) );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(n37782), .D(N265), .Q(
        \REGISTERS[26][21] ) );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(n37782), .D(N264), .Q(
        \REGISTERS[26][20] ) );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n37782), .D(N263), .Q(
        \REGISTERS[26][19] ) );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(N280), .D(N262), .Q(\REGISTERS[26][18] )
         );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n37782), .D(N261), .Q(
        \REGISTERS[26][17] ) );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(N280), .D(N260), .Q(\REGISTERS[26][16] )
         );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(n37782), .D(N259), .Q(
        \REGISTERS[26][15] ) );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(N280), .D(N258), .Q(\REGISTERS[26][14] )
         );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(N280), .D(N257), .Q(\REGISTERS[26][13] )
         );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(N280), .D(N256), .Q(\REGISTERS[26][12] )
         );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(N280), .D(N255), .Q(\REGISTERS[26][11] )
         );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n37782), .D(N254), .Q(
        \REGISTERS[26][10] ) );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(N280), .D(N253), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(N280), .D(N252), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n37782), .D(N251), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(n37782), .D(N250), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(N280), .D(N249), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(N280), .D(N248), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(N280), .D(N247), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(N280), .D(N246), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(n37782), .D(N245), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(N280), .D(N244), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(n37783), .D(N275), .Q(
        \REGISTERS[27][31] ) );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(n37783), .D(N274), .Q(
        \REGISTERS[27][30] ) );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(n37783), .D(N273), .Q(
        \REGISTERS[27][29] ) );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(n37783), .D(N272), .Q(
        \REGISTERS[27][28] ) );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(n37783), .D(N271), .Q(
        \REGISTERS[27][27] ) );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(n37783), .D(N270), .Q(
        \REGISTERS[27][26] ) );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(N279), .D(N269), .Q(\REGISTERS[27][25] )
         );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(N279), .D(N268), .Q(\REGISTERS[27][24] )
         );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n37783), .D(N267), .Q(
        \REGISTERS[27][23] ) );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n37783), .D(N266), .Q(
        \REGISTERS[27][22] ) );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(n37783), .D(N265), .Q(
        \REGISTERS[27][21] ) );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(n37783), .D(N264), .Q(
        \REGISTERS[27][20] ) );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n37783), .D(N263), .Q(
        \REGISTERS[27][19] ) );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(N279), .D(N262), .Q(\REGISTERS[27][18] )
         );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n37783), .D(N261), .Q(
        \REGISTERS[27][17] ) );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(N279), .D(N260), .Q(\REGISTERS[27][16] )
         );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(n37783), .D(N259), .Q(
        \REGISTERS[27][15] ) );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(N279), .D(N258), .Q(\REGISTERS[27][14] )
         );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(N279), .D(N257), .Q(\REGISTERS[27][13] )
         );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(N279), .D(N256), .Q(\REGISTERS[27][12] )
         );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(N279), .D(N255), .Q(\REGISTERS[27][11] )
         );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n37783), .D(N254), .Q(
        \REGISTERS[27][10] ) );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(N279), .D(N253), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(N279), .D(N252), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n37783), .D(N251), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(n37783), .D(N250), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(N279), .D(N249), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(N279), .D(N248), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(N279), .D(N247), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(N279), .D(N246), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(n37783), .D(N245), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(N279), .D(N244), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(n37784), .D(N275), .Q(
        \REGISTERS[28][31] ) );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(n37784), .D(N274), .Q(
        \REGISTERS[28][30] ) );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(n37784), .D(N273), .Q(
        \REGISTERS[28][29] ) );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(n37784), .D(N272), .Q(
        \REGISTERS[28][28] ) );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(n37784), .D(N271), .Q(
        \REGISTERS[28][27] ) );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(n37784), .D(N270), .Q(
        \REGISTERS[28][26] ) );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(N278), .D(N269), .Q(\REGISTERS[28][25] )
         );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(N278), .D(N268), .Q(\REGISTERS[28][24] )
         );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n37784), .D(N267), .Q(
        \REGISTERS[28][23] ) );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n37784), .D(N266), .Q(
        \REGISTERS[28][22] ) );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(n37784), .D(N265), .Q(
        \REGISTERS[28][21] ) );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(n37784), .D(N264), .Q(
        \REGISTERS[28][20] ) );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n37784), .D(N263), .Q(
        \REGISTERS[28][19] ) );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(N278), .D(N262), .Q(\REGISTERS[28][18] )
         );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n37784), .D(N261), .Q(
        \REGISTERS[28][17] ) );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(N278), .D(N260), .Q(\REGISTERS[28][16] )
         );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(n37784), .D(N259), .Q(
        \REGISTERS[28][15] ) );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(N278), .D(N258), .Q(\REGISTERS[28][14] )
         );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(N278), .D(N257), .Q(\REGISTERS[28][13] )
         );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(N278), .D(N256), .Q(\REGISTERS[28][12] )
         );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(N278), .D(N255), .Q(\REGISTERS[28][11] )
         );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n37784), .D(N254), .Q(
        \REGISTERS[28][10] ) );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(N278), .D(N253), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(N278), .D(N252), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n37784), .D(N251), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(n37784), .D(N250), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(N278), .D(N249), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(N278), .D(N248), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(N278), .D(N247), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(N278), .D(N246), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(n37784), .D(N245), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(N278), .D(N244), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(n37785), .D(N275), .Q(
        \REGISTERS[29][31] ) );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(n37785), .D(N274), .Q(
        \REGISTERS[29][30] ) );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(n37785), .D(N273), .Q(
        \REGISTERS[29][29] ) );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(n37785), .D(N272), .Q(
        \REGISTERS[29][28] ) );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(n37785), .D(N271), .Q(
        \REGISTERS[29][27] ) );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(n37785), .D(N270), .Q(
        \REGISTERS[29][26] ) );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(N277), .D(N269), .Q(\REGISTERS[29][25] )
         );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(N277), .D(N268), .Q(\REGISTERS[29][24] )
         );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n37785), .D(N267), .Q(
        \REGISTERS[29][23] ) );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n37785), .D(N266), .Q(
        \REGISTERS[29][22] ) );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(n37785), .D(N265), .Q(
        \REGISTERS[29][21] ) );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(n37785), .D(N264), .Q(
        \REGISTERS[29][20] ) );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n37785), .D(N263), .Q(
        \REGISTERS[29][19] ) );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(N277), .D(N262), .Q(\REGISTERS[29][18] )
         );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n37785), .D(N261), .Q(
        \REGISTERS[29][17] ) );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(N277), .D(N260), .Q(\REGISTERS[29][16] )
         );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(n37785), .D(N259), .Q(
        \REGISTERS[29][15] ) );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(N277), .D(N258), .Q(\REGISTERS[29][14] )
         );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(N277), .D(N257), .Q(\REGISTERS[29][13] )
         );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(N277), .D(N256), .Q(\REGISTERS[29][12] )
         );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(N277), .D(N255), .Q(\REGISTERS[29][11] )
         );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n37785), .D(N254), .Q(
        \REGISTERS[29][10] ) );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(N277), .D(N253), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(N277), .D(N252), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n37785), .D(N251), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(n37785), .D(N250), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(N277), .D(N249), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(N277), .D(N248), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(N277), .D(N247), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(N277), .D(N246), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(n37785), .D(N245), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(N277), .D(N244), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(n37786), .D(N275), .Q(
        \REGISTERS[30][31] ) );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(n37786), .D(N274), .Q(
        \REGISTERS[30][30] ) );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(n37786), .D(N273), .Q(
        \REGISTERS[30][29] ) );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(n37786), .D(N272), .Q(
        \REGISTERS[30][28] ) );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(n37786), .D(N271), .Q(
        \REGISTERS[30][27] ) );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(n37786), .D(N270), .Q(
        \REGISTERS[30][26] ) );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(N276), .D(N269), .Q(\REGISTERS[30][25] )
         );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(N276), .D(N268), .Q(\REGISTERS[30][24] )
         );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n37786), .D(N267), .Q(
        \REGISTERS[30][23] ) );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n37786), .D(N266), .Q(
        \REGISTERS[30][22] ) );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(n37786), .D(N265), .Q(
        \REGISTERS[30][21] ) );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(n37786), .D(N264), .Q(
        \REGISTERS[30][20] ) );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n37786), .D(N263), .Q(
        \REGISTERS[30][19] ) );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(N276), .D(N262), .Q(\REGISTERS[30][18] )
         );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n37786), .D(N261), .Q(
        \REGISTERS[30][17] ) );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(N276), .D(N260), .Q(\REGISTERS[30][16] )
         );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(n37786), .D(N259), .Q(
        \REGISTERS[30][15] ) );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(N276), .D(N258), .Q(\REGISTERS[30][14] )
         );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(N276), .D(N257), .Q(\REGISTERS[30][13] )
         );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(N276), .D(N256), .Q(\REGISTERS[30][12] )
         );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(N276), .D(N255), .Q(\REGISTERS[30][11] )
         );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n37786), .D(N254), .Q(
        \REGISTERS[30][10] ) );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(N276), .D(N253), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(N276), .D(N252), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n37786), .D(N251), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(n37786), .D(N250), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(N276), .D(N249), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(N276), .D(N248), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(N276), .D(N247), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(N276), .D(N246), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(n37786), .D(N245), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(N276), .D(N244), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(n37787), .D(N275), .Q(
        \REGISTERS[31][31] ) );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(n37787), .D(N274), .Q(
        \REGISTERS[31][30] ) );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(n37787), .D(N273), .Q(
        \REGISTERS[31][29] ) );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(n37787), .D(N272), .Q(
        \REGISTERS[31][28] ) );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(n37787), .D(N271), .Q(
        \REGISTERS[31][27] ) );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(n37787), .D(N270), .Q(
        \REGISTERS[31][26] ) );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(n37787), .D(N269), .Q(
        \REGISTERS[31][25] ) );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(n37787), .D(N268), .Q(
        \REGISTERS[31][24] ) );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(n37787), .D(N267), .Q(
        \REGISTERS[31][23] ) );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(n37787), .D(N266), .Q(
        \REGISTERS[31][22] ) );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n37787), .D(N265), .Q(
        \REGISTERS[31][21] ) );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(N243), .D(N264), .Q(\REGISTERS[31][20] )
         );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n37787), .D(N263), .Q(
        \REGISTERS[31][19] ) );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(N243), .D(N262), .Q(\REGISTERS[31][18] )
         );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n37787), .D(N261), .Q(
        \REGISTERS[31][17] ) );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(N243), .D(N260), .Q(\REGISTERS[31][16] )
         );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(n37787), .D(N259), .Q(
        \REGISTERS[31][15] ) );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(N243), .D(N258), .Q(\REGISTERS[31][14] )
         );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(N243), .D(N257), .Q(\REGISTERS[31][13] )
         );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(N243), .D(N256), .Q(\REGISTERS[31][12] )
         );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n37787), .D(N255), .Q(
        \REGISTERS[31][11] ) );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n37787), .D(N254), .Q(
        \REGISTERS[31][10] ) );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(N243), .D(N253), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(N243), .D(N252), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(N243), .D(N251), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(N243), .D(N250), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(N243), .D(N249), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(N243), .D(N248), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(N243), .D(N247), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(N243), .D(N246), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(N243), .D(N245), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n37787), .D(N244), .Q(\REGISTERS[31][0] )
         );
  AOI22_X1 U3 ( .A1(\REGISTERS[29][17] ), .A2(n37741), .B1(\REGISTERS[30][17] ), .B2(n37742), .ZN(n36859) );
  AOI22_X1 U4 ( .A1(\REGISTERS[4][17] ), .A2(n37743), .B1(\REGISTERS[27][17] ), 
        .B2(n37744), .ZN(n36860) );
  AOI22_X1 U5 ( .A1(\REGISTERS[28][17] ), .A2(n37745), .B1(\REGISTERS[10][17] ), .B2(n37746), .ZN(n36861) );
  AOI22_X1 U6 ( .A1(\REGISTERS[7][17] ), .A2(n37747), .B1(\REGISTERS[6][17] ), 
        .B2(n37748), .ZN(n36862) );
  NAND4_X1 U7 ( .A1(n36859), .A2(n36860), .A3(n36861), .A4(n36862), .ZN(n36863) );
  AOI22_X1 U8 ( .A1(\REGISTERS[5][17] ), .A2(n37749), .B1(\REGISTERS[26][17] ), 
        .B2(n37750), .ZN(n36864) );
  AOI22_X1 U9 ( .A1(\REGISTERS[25][17] ), .A2(n37751), .B1(\REGISTERS[21][17] ), .B2(n37752), .ZN(n36865) );
  AOI22_X1 U10 ( .A1(\REGISTERS[17][17] ), .A2(n37753), .B1(
        \REGISTERS[23][17] ), .B2(n37754), .ZN(n36866) );
  AOI22_X1 U11 ( .A1(\REGISTERS[19][17] ), .A2(n37755), .B1(
        \REGISTERS[14][17] ), .B2(n37756), .ZN(n36867) );
  NAND4_X1 U12 ( .A1(n36864), .A2(n36865), .A3(n36866), .A4(n36867), .ZN(
        n36868) );
  AOI22_X1 U13 ( .A1(\REGISTERS[16][17] ), .A2(n37726), .B1(
        \REGISTERS[11][17] ), .B2(n37727), .ZN(n36869) );
  AOI22_X1 U14 ( .A1(\REGISTERS[24][17] ), .A2(n37728), .B1(\REGISTERS[1][17] ), .B2(n37729), .ZN(n36870) );
  AOI222_X1 U15 ( .A1(\REGISTERS[15][17] ), .A2(n37730), .B1(
        \REGISTERS[12][17] ), .B2(n37731), .C1(\REGISTERS[13][17] ), .C2(
        n37732), .ZN(n36871) );
  NAND3_X1 U16 ( .A1(n36869), .A2(n36870), .A3(n36871), .ZN(n36872) );
  AOI22_X1 U17 ( .A1(\REGISTERS[22][17] ), .A2(n37733), .B1(
        \REGISTERS[20][17] ), .B2(n37734), .ZN(n36873) );
  AOI22_X1 U18 ( .A1(\REGISTERS[9][17] ), .A2(n37735), .B1(\REGISTERS[18][17] ), .B2(n37736), .ZN(n36874) );
  AOI22_X1 U19 ( .A1(\REGISTERS[31][17] ), .A2(n37737), .B1(\REGISTERS[2][17] ), .B2(n37738), .ZN(n36875) );
  AOI22_X1 U20 ( .A1(\REGISTERS[8][17] ), .A2(n37739), .B1(\REGISTERS[3][17] ), 
        .B2(n37740), .ZN(n36876) );
  NAND4_X1 U21 ( .A1(n36873), .A2(n36874), .A3(n36875), .A4(n36876), .ZN(
        n36877) );
  OR4_X1 U22 ( .A1(n36863), .A2(n36868), .A3(n36872), .A4(n36877), .ZN(
        OUTA[17]) );
  AOI22_X1 U23 ( .A1(\REGISTERS[29][16] ), .A2(n37741), .B1(
        \REGISTERS[30][16] ), .B2(n37742), .ZN(n36878) );
  AOI22_X1 U24 ( .A1(\REGISTERS[4][16] ), .A2(n37743), .B1(\REGISTERS[27][16] ), .B2(n37744), .ZN(n36879) );
  AOI22_X1 U25 ( .A1(\REGISTERS[28][16] ), .A2(n37745), .B1(
        \REGISTERS[10][16] ), .B2(n37746), .ZN(n36880) );
  AOI22_X1 U26 ( .A1(\REGISTERS[7][16] ), .A2(n37747), .B1(\REGISTERS[6][16] ), 
        .B2(n37748), .ZN(n36881) );
  NAND4_X1 U27 ( .A1(n36878), .A2(n36879), .A3(n36880), .A4(n36881), .ZN(
        n36882) );
  AOI22_X1 U28 ( .A1(\REGISTERS[5][16] ), .A2(n37749), .B1(\REGISTERS[26][16] ), .B2(n37750), .ZN(n36883) );
  AOI22_X1 U29 ( .A1(\REGISTERS[25][16] ), .A2(n37751), .B1(
        \REGISTERS[21][16] ), .B2(n37752), .ZN(n36884) );
  AOI22_X1 U30 ( .A1(\REGISTERS[17][16] ), .A2(n37753), .B1(
        \REGISTERS[23][16] ), .B2(n37754), .ZN(n36885) );
  AOI22_X1 U31 ( .A1(\REGISTERS[19][16] ), .A2(n37755), .B1(
        \REGISTERS[14][16] ), .B2(n37756), .ZN(n36886) );
  NAND4_X1 U32 ( .A1(n36883), .A2(n36884), .A3(n36885), .A4(n36886), .ZN(
        n36887) );
  AOI22_X1 U33 ( .A1(\REGISTERS[16][16] ), .A2(n37726), .B1(
        \REGISTERS[11][16] ), .B2(n37727), .ZN(n36888) );
  AOI22_X1 U34 ( .A1(\REGISTERS[24][16] ), .A2(n37728), .B1(\REGISTERS[1][16] ), .B2(n37729), .ZN(n36889) );
  AOI222_X1 U35 ( .A1(\REGISTERS[15][16] ), .A2(n37730), .B1(
        \REGISTERS[12][16] ), .B2(n37731), .C1(\REGISTERS[13][16] ), .C2(
        n37732), .ZN(n36890) );
  NAND3_X1 U36 ( .A1(n36888), .A2(n36889), .A3(n36890), .ZN(n36891) );
  AOI22_X1 U37 ( .A1(\REGISTERS[22][16] ), .A2(n37733), .B1(
        \REGISTERS[20][16] ), .B2(n37734), .ZN(n36892) );
  AOI22_X1 U38 ( .A1(\REGISTERS[9][16] ), .A2(n37735), .B1(\REGISTERS[18][16] ), .B2(n37736), .ZN(n36893) );
  AOI22_X1 U39 ( .A1(\REGISTERS[31][16] ), .A2(n37737), .B1(\REGISTERS[2][16] ), .B2(n37738), .ZN(n36894) );
  AOI22_X1 U40 ( .A1(\REGISTERS[8][16] ), .A2(n37739), .B1(\REGISTERS[3][16] ), 
        .B2(n37740), .ZN(n36895) );
  NAND4_X1 U41 ( .A1(n36892), .A2(n36893), .A3(n36894), .A4(n36895), .ZN(
        n36896) );
  OR4_X1 U42 ( .A1(n36882), .A2(n36887), .A3(n36891), .A4(n36896), .ZN(
        OUTA[16]) );
  AOI22_X1 U43 ( .A1(\REGISTERS[29][15] ), .A2(n37741), .B1(
        \REGISTERS[30][15] ), .B2(n37742), .ZN(n36897) );
  AOI22_X1 U44 ( .A1(\REGISTERS[4][15] ), .A2(n37743), .B1(\REGISTERS[27][15] ), .B2(n37744), .ZN(n36898) );
  AOI22_X1 U45 ( .A1(\REGISTERS[28][15] ), .A2(n37745), .B1(
        \REGISTERS[10][15] ), .B2(n37746), .ZN(n36899) );
  AOI22_X1 U46 ( .A1(\REGISTERS[7][15] ), .A2(n37747), .B1(\REGISTERS[6][15] ), 
        .B2(n37748), .ZN(n36900) );
  NAND4_X1 U47 ( .A1(n36897), .A2(n36898), .A3(n36899), .A4(n36900), .ZN(
        n36901) );
  AOI22_X1 U48 ( .A1(\REGISTERS[5][15] ), .A2(n37749), .B1(\REGISTERS[26][15] ), .B2(n37750), .ZN(n36902) );
  AOI22_X1 U49 ( .A1(\REGISTERS[25][15] ), .A2(n37751), .B1(
        \REGISTERS[21][15] ), .B2(n37752), .ZN(n36903) );
  AOI22_X1 U50 ( .A1(\REGISTERS[17][15] ), .A2(n37753), .B1(
        \REGISTERS[23][15] ), .B2(n37754), .ZN(n36904) );
  AOI22_X1 U51 ( .A1(\REGISTERS[19][15] ), .A2(n37755), .B1(
        \REGISTERS[14][15] ), .B2(n37756), .ZN(n36905) );
  NAND4_X1 U52 ( .A1(n36902), .A2(n36903), .A3(n36904), .A4(n36905), .ZN(
        n36906) );
  AOI22_X1 U53 ( .A1(\REGISTERS[16][15] ), .A2(n37726), .B1(
        \REGISTERS[11][15] ), .B2(n37727), .ZN(n36907) );
  AOI22_X1 U54 ( .A1(\REGISTERS[24][15] ), .A2(n37728), .B1(\REGISTERS[1][15] ), .B2(n37729), .ZN(n36908) );
  AOI222_X1 U55 ( .A1(\REGISTERS[15][15] ), .A2(n37730), .B1(
        \REGISTERS[12][15] ), .B2(n37731), .C1(\REGISTERS[13][15] ), .C2(
        n37732), .ZN(n36909) );
  NAND3_X1 U56 ( .A1(n36907), .A2(n36908), .A3(n36909), .ZN(n36910) );
  AOI22_X1 U57 ( .A1(\REGISTERS[22][15] ), .A2(n37733), .B1(
        \REGISTERS[20][15] ), .B2(n37734), .ZN(n36911) );
  AOI22_X1 U58 ( .A1(\REGISTERS[9][15] ), .A2(n37735), .B1(\REGISTERS[18][15] ), .B2(n37736), .ZN(n36912) );
  AOI22_X1 U59 ( .A1(\REGISTERS[31][15] ), .A2(n37737), .B1(\REGISTERS[2][15] ), .B2(n37738), .ZN(n36913) );
  AOI22_X1 U60 ( .A1(\REGISTERS[8][15] ), .A2(n37739), .B1(\REGISTERS[3][15] ), 
        .B2(n37740), .ZN(n36914) );
  NAND4_X1 U61 ( .A1(n36911), .A2(n36912), .A3(n36913), .A4(n36914), .ZN(
        n36915) );
  OR4_X1 U62 ( .A1(n36901), .A2(n36906), .A3(n36910), .A4(n36915), .ZN(
        OUTA[15]) );
  AOI22_X1 U63 ( .A1(\REGISTERS[29][14] ), .A2(n37741), .B1(
        \REGISTERS[30][14] ), .B2(n37742), .ZN(n36916) );
  AOI22_X1 U64 ( .A1(\REGISTERS[4][14] ), .A2(n37743), .B1(\REGISTERS[27][14] ), .B2(n37744), .ZN(n36917) );
  AOI22_X1 U65 ( .A1(\REGISTERS[28][14] ), .A2(n37745), .B1(
        \REGISTERS[10][14] ), .B2(n37746), .ZN(n36918) );
  AOI22_X1 U66 ( .A1(\REGISTERS[7][14] ), .A2(n37747), .B1(\REGISTERS[6][14] ), 
        .B2(n37748), .ZN(n36919) );
  NAND4_X1 U67 ( .A1(n36916), .A2(n36917), .A3(n36918), .A4(n36919), .ZN(
        n36920) );
  AOI22_X1 U68 ( .A1(\REGISTERS[5][14] ), .A2(n37749), .B1(\REGISTERS[26][14] ), .B2(n37750), .ZN(n36921) );
  AOI22_X1 U69 ( .A1(\REGISTERS[25][14] ), .A2(n37751), .B1(
        \REGISTERS[21][14] ), .B2(n37752), .ZN(n36922) );
  AOI22_X1 U70 ( .A1(\REGISTERS[17][14] ), .A2(n37753), .B1(
        \REGISTERS[23][14] ), .B2(n37754), .ZN(n36923) );
  AOI22_X1 U71 ( .A1(\REGISTERS[19][14] ), .A2(n37755), .B1(
        \REGISTERS[14][14] ), .B2(n37756), .ZN(n36924) );
  NAND4_X1 U72 ( .A1(n36921), .A2(n36922), .A3(n36923), .A4(n36924), .ZN(
        n36925) );
  AOI22_X1 U73 ( .A1(\REGISTERS[16][14] ), .A2(n37726), .B1(
        \REGISTERS[11][14] ), .B2(n37727), .ZN(n36926) );
  AOI22_X1 U74 ( .A1(\REGISTERS[24][14] ), .A2(n37728), .B1(\REGISTERS[1][14] ), .B2(n37729), .ZN(n36927) );
  AOI222_X1 U75 ( .A1(\REGISTERS[15][14] ), .A2(n37730), .B1(
        \REGISTERS[12][14] ), .B2(n37731), .C1(\REGISTERS[13][14] ), .C2(
        n37732), .ZN(n36928) );
  NAND3_X1 U76 ( .A1(n36926), .A2(n36927), .A3(n36928), .ZN(n36929) );
  AOI22_X1 U77 ( .A1(\REGISTERS[22][14] ), .A2(n37733), .B1(
        \REGISTERS[20][14] ), .B2(n37734), .ZN(n36930) );
  AOI22_X1 U78 ( .A1(\REGISTERS[9][14] ), .A2(n37735), .B1(\REGISTERS[18][14] ), .B2(n37736), .ZN(n36931) );
  AOI22_X1 U79 ( .A1(\REGISTERS[31][14] ), .A2(n37737), .B1(\REGISTERS[2][14] ), .B2(n37738), .ZN(n36932) );
  AOI22_X1 U80 ( .A1(\REGISTERS[8][14] ), .A2(n37739), .B1(\REGISTERS[3][14] ), 
        .B2(n37740), .ZN(n36933) );
  NAND4_X1 U81 ( .A1(n36930), .A2(n36931), .A3(n36932), .A4(n36933), .ZN(
        n36934) );
  OR4_X1 U82 ( .A1(n36920), .A2(n36925), .A3(n36929), .A4(n36934), .ZN(
        OUTA[14]) );
  AOI22_X1 U83 ( .A1(\REGISTERS[29][13] ), .A2(n37741), .B1(
        \REGISTERS[30][13] ), .B2(n37742), .ZN(n36935) );
  AOI22_X1 U84 ( .A1(\REGISTERS[4][13] ), .A2(n37743), .B1(\REGISTERS[27][13] ), .B2(n37744), .ZN(n36936) );
  AOI22_X1 U85 ( .A1(\REGISTERS[28][13] ), .A2(n37745), .B1(
        \REGISTERS[10][13] ), .B2(n37746), .ZN(n36937) );
  AOI22_X1 U86 ( .A1(\REGISTERS[7][13] ), .A2(n37747), .B1(\REGISTERS[6][13] ), 
        .B2(n37748), .ZN(n36938) );
  NAND4_X1 U87 ( .A1(n36935), .A2(n36936), .A3(n36937), .A4(n36938), .ZN(
        n36939) );
  AOI22_X1 U88 ( .A1(\REGISTERS[5][13] ), .A2(n37749), .B1(\REGISTERS[26][13] ), .B2(n37750), .ZN(n36940) );
  AOI22_X1 U89 ( .A1(\REGISTERS[25][13] ), .A2(n37751), .B1(
        \REGISTERS[21][13] ), .B2(n37752), .ZN(n36941) );
  AOI22_X1 U90 ( .A1(\REGISTERS[17][13] ), .A2(n37753), .B1(
        \REGISTERS[23][13] ), .B2(n37754), .ZN(n36942) );
  AOI22_X1 U91 ( .A1(\REGISTERS[19][13] ), .A2(n37755), .B1(
        \REGISTERS[14][13] ), .B2(n37756), .ZN(n36943) );
  NAND4_X1 U92 ( .A1(n36940), .A2(n36941), .A3(n36942), .A4(n36943), .ZN(
        n36944) );
  AOI22_X1 U93 ( .A1(\REGISTERS[16][13] ), .A2(n37726), .B1(
        \REGISTERS[11][13] ), .B2(n37727), .ZN(n36945) );
  AOI22_X1 U94 ( .A1(\REGISTERS[24][13] ), .A2(n37728), .B1(\REGISTERS[1][13] ), .B2(n37729), .ZN(n36946) );
  AOI222_X1 U95 ( .A1(\REGISTERS[15][13] ), .A2(n37730), .B1(
        \REGISTERS[12][13] ), .B2(n37731), .C1(\REGISTERS[13][13] ), .C2(
        n37732), .ZN(n36947) );
  NAND3_X1 U96 ( .A1(n36945), .A2(n36946), .A3(n36947), .ZN(n36948) );
  AOI22_X1 U97 ( .A1(\REGISTERS[22][13] ), .A2(n37733), .B1(
        \REGISTERS[20][13] ), .B2(n37734), .ZN(n36949) );
  AOI22_X1 U98 ( .A1(\REGISTERS[9][13] ), .A2(n37735), .B1(\REGISTERS[18][13] ), .B2(n37736), .ZN(n36950) );
  AOI22_X1 U99 ( .A1(\REGISTERS[31][13] ), .A2(n37737), .B1(\REGISTERS[2][13] ), .B2(n37738), .ZN(n36951) );
  AOI22_X1 U100 ( .A1(\REGISTERS[8][13] ), .A2(n37739), .B1(\REGISTERS[3][13] ), .B2(n37740), .ZN(n36952) );
  NAND4_X1 U101 ( .A1(n36949), .A2(n36950), .A3(n36951), .A4(n36952), .ZN(
        n36953) );
  OR4_X1 U102 ( .A1(n36939), .A2(n36944), .A3(n36948), .A4(n36953), .ZN(
        OUTA[13]) );
  AOI22_X1 U103 ( .A1(\REGISTERS[29][12] ), .A2(n37741), .B1(
        \REGISTERS[30][12] ), .B2(n37742), .ZN(n36954) );
  AOI22_X1 U104 ( .A1(\REGISTERS[4][12] ), .A2(n37743), .B1(
        \REGISTERS[27][12] ), .B2(n37744), .ZN(n36955) );
  AOI22_X1 U105 ( .A1(\REGISTERS[28][12] ), .A2(n37745), .B1(
        \REGISTERS[10][12] ), .B2(n37746), .ZN(n36956) );
  AOI22_X1 U106 ( .A1(\REGISTERS[7][12] ), .A2(n37747), .B1(\REGISTERS[6][12] ), .B2(n37748), .ZN(n36957) );
  NAND4_X1 U107 ( .A1(n36954), .A2(n36955), .A3(n36956), .A4(n36957), .ZN(
        n36958) );
  AOI22_X1 U108 ( .A1(\REGISTERS[5][12] ), .A2(n37749), .B1(
        \REGISTERS[26][12] ), .B2(n37750), .ZN(n36959) );
  AOI22_X1 U109 ( .A1(\REGISTERS[25][12] ), .A2(n37751), .B1(
        \REGISTERS[21][12] ), .B2(n37752), .ZN(n36960) );
  AOI22_X1 U110 ( .A1(\REGISTERS[17][12] ), .A2(n37753), .B1(
        \REGISTERS[23][12] ), .B2(n37754), .ZN(n36961) );
  AOI22_X1 U111 ( .A1(\REGISTERS[19][12] ), .A2(n37755), .B1(
        \REGISTERS[14][12] ), .B2(n37756), .ZN(n36962) );
  NAND4_X1 U112 ( .A1(n36959), .A2(n36960), .A3(n36961), .A4(n36962), .ZN(
        n36963) );
  AOI22_X1 U113 ( .A1(\REGISTERS[16][12] ), .A2(n37726), .B1(
        \REGISTERS[11][12] ), .B2(n37727), .ZN(n36964) );
  AOI22_X1 U114 ( .A1(\REGISTERS[24][12] ), .A2(n37728), .B1(
        \REGISTERS[1][12] ), .B2(n37729), .ZN(n36965) );
  AOI222_X1 U115 ( .A1(\REGISTERS[15][12] ), .A2(n37730), .B1(
        \REGISTERS[12][12] ), .B2(n37731), .C1(\REGISTERS[13][12] ), .C2(
        n37732), .ZN(n36966) );
  NAND3_X1 U116 ( .A1(n36964), .A2(n36965), .A3(n36966), .ZN(n36967) );
  AOI22_X1 U117 ( .A1(\REGISTERS[22][12] ), .A2(n37733), .B1(
        \REGISTERS[20][12] ), .B2(n37734), .ZN(n36968) );
  AOI22_X1 U118 ( .A1(\REGISTERS[9][12] ), .A2(n37735), .B1(
        \REGISTERS[18][12] ), .B2(n37736), .ZN(n36969) );
  AOI22_X1 U119 ( .A1(\REGISTERS[31][12] ), .A2(n37737), .B1(
        \REGISTERS[2][12] ), .B2(n37738), .ZN(n36970) );
  AOI22_X1 U120 ( .A1(\REGISTERS[8][12] ), .A2(n37739), .B1(\REGISTERS[3][12] ), .B2(n37740), .ZN(n36971) );
  NAND4_X1 U121 ( .A1(n36968), .A2(n36969), .A3(n36970), .A4(n36971), .ZN(
        n36972) );
  OR4_X1 U122 ( .A1(n36958), .A2(n36963), .A3(n36967), .A4(n36972), .ZN(
        OUTA[12]) );
  AOI22_X1 U123 ( .A1(\REGISTERS[29][11] ), .A2(n37741), .B1(
        \REGISTERS[30][11] ), .B2(n37742), .ZN(n36973) );
  AOI22_X1 U124 ( .A1(\REGISTERS[4][11] ), .A2(n37743), .B1(
        \REGISTERS[27][11] ), .B2(n37744), .ZN(n36974) );
  AOI22_X1 U125 ( .A1(\REGISTERS[28][11] ), .A2(n37745), .B1(
        \REGISTERS[10][11] ), .B2(n37746), .ZN(n36975) );
  AOI22_X1 U126 ( .A1(\REGISTERS[7][11] ), .A2(n37747), .B1(\REGISTERS[6][11] ), .B2(n37748), .ZN(n36976) );
  NAND4_X1 U127 ( .A1(n36973), .A2(n36974), .A3(n36975), .A4(n36976), .ZN(
        n36977) );
  AOI22_X1 U128 ( .A1(\REGISTERS[5][11] ), .A2(n37749), .B1(
        \REGISTERS[26][11] ), .B2(n37750), .ZN(n36978) );
  AOI22_X1 U129 ( .A1(\REGISTERS[25][11] ), .A2(n37751), .B1(
        \REGISTERS[21][11] ), .B2(n37752), .ZN(n36979) );
  AOI22_X1 U130 ( .A1(\REGISTERS[17][11] ), .A2(n37753), .B1(
        \REGISTERS[23][11] ), .B2(n37754), .ZN(n36980) );
  AOI22_X1 U131 ( .A1(\REGISTERS[19][11] ), .A2(n37755), .B1(
        \REGISTERS[14][11] ), .B2(n37756), .ZN(n36981) );
  NAND4_X1 U132 ( .A1(n36978), .A2(n36979), .A3(n36980), .A4(n36981), .ZN(
        n36982) );
  AOI22_X1 U133 ( .A1(\REGISTERS[16][11] ), .A2(n37726), .B1(
        \REGISTERS[11][11] ), .B2(n37727), .ZN(n36983) );
  AOI22_X1 U134 ( .A1(\REGISTERS[24][11] ), .A2(n37728), .B1(
        \REGISTERS[1][11] ), .B2(n37729), .ZN(n36984) );
  AOI222_X1 U135 ( .A1(\REGISTERS[15][11] ), .A2(n37730), .B1(
        \REGISTERS[12][11] ), .B2(n37731), .C1(\REGISTERS[13][11] ), .C2(
        n37732), .ZN(n36985) );
  NAND3_X1 U136 ( .A1(n36983), .A2(n36984), .A3(n36985), .ZN(n36986) );
  AOI22_X1 U137 ( .A1(\REGISTERS[22][11] ), .A2(n37733), .B1(
        \REGISTERS[20][11] ), .B2(n37734), .ZN(n36987) );
  AOI22_X1 U138 ( .A1(\REGISTERS[9][11] ), .A2(n37735), .B1(
        \REGISTERS[18][11] ), .B2(n37736), .ZN(n36988) );
  AOI22_X1 U139 ( .A1(\REGISTERS[31][11] ), .A2(n37737), .B1(
        \REGISTERS[2][11] ), .B2(n37738), .ZN(n36989) );
  AOI22_X1 U140 ( .A1(\REGISTERS[8][11] ), .A2(n37739), .B1(\REGISTERS[3][11] ), .B2(n37740), .ZN(n36990) );
  NAND4_X1 U141 ( .A1(n36987), .A2(n36988), .A3(n36989), .A4(n36990), .ZN(
        n36991) );
  OR4_X1 U142 ( .A1(n36977), .A2(n36982), .A3(n36986), .A4(n36991), .ZN(
        OUTA[11]) );
  AOI22_X1 U143 ( .A1(\REGISTERS[29][10] ), .A2(n37741), .B1(
        \REGISTERS[30][10] ), .B2(n37742), .ZN(n36992) );
  AOI22_X1 U144 ( .A1(\REGISTERS[4][10] ), .A2(n37743), .B1(
        \REGISTERS[27][10] ), .B2(n37744), .ZN(n36993) );
  AOI22_X1 U145 ( .A1(\REGISTERS[28][10] ), .A2(n37745), .B1(
        \REGISTERS[10][10] ), .B2(n37746), .ZN(n36994) );
  AOI22_X1 U146 ( .A1(\REGISTERS[7][10] ), .A2(n37747), .B1(\REGISTERS[6][10] ), .B2(n37748), .ZN(n36995) );
  NAND4_X1 U147 ( .A1(n36992), .A2(n36993), .A3(n36994), .A4(n36995), .ZN(
        n36996) );
  AOI22_X1 U148 ( .A1(\REGISTERS[5][10] ), .A2(n37749), .B1(
        \REGISTERS[26][10] ), .B2(n37750), .ZN(n36997) );
  AOI22_X1 U149 ( .A1(\REGISTERS[25][10] ), .A2(n37751), .B1(
        \REGISTERS[21][10] ), .B2(n37752), .ZN(n36998) );
  AOI22_X1 U150 ( .A1(\REGISTERS[17][10] ), .A2(n37753), .B1(
        \REGISTERS[23][10] ), .B2(n37754), .ZN(n36999) );
  AOI22_X1 U151 ( .A1(\REGISTERS[19][10] ), .A2(n37755), .B1(
        \REGISTERS[14][10] ), .B2(n37756), .ZN(n37000) );
  NAND4_X1 U152 ( .A1(n36997), .A2(n36998), .A3(n36999), .A4(n37000), .ZN(
        n37001) );
  AOI22_X1 U153 ( .A1(\REGISTERS[16][10] ), .A2(n37726), .B1(
        \REGISTERS[11][10] ), .B2(n37727), .ZN(n37002) );
  AOI22_X1 U154 ( .A1(\REGISTERS[24][10] ), .A2(n37728), .B1(
        \REGISTERS[1][10] ), .B2(n37729), .ZN(n37003) );
  AOI222_X1 U155 ( .A1(\REGISTERS[15][10] ), .A2(n37730), .B1(
        \REGISTERS[12][10] ), .B2(n37731), .C1(\REGISTERS[13][10] ), .C2(
        n37732), .ZN(n37004) );
  NAND3_X1 U156 ( .A1(n37002), .A2(n37003), .A3(n37004), .ZN(n37005) );
  AOI22_X1 U157 ( .A1(\REGISTERS[22][10] ), .A2(n37733), .B1(
        \REGISTERS[20][10] ), .B2(n37734), .ZN(n37006) );
  AOI22_X1 U158 ( .A1(\REGISTERS[9][10] ), .A2(n37735), .B1(
        \REGISTERS[18][10] ), .B2(n37736), .ZN(n37007) );
  AOI22_X1 U159 ( .A1(\REGISTERS[31][10] ), .A2(n37737), .B1(
        \REGISTERS[2][10] ), .B2(n37738), .ZN(n37008) );
  AOI22_X1 U160 ( .A1(\REGISTERS[8][10] ), .A2(n37739), .B1(\REGISTERS[3][10] ), .B2(n37740), .ZN(n37009) );
  NAND4_X1 U161 ( .A1(n37006), .A2(n37007), .A3(n37008), .A4(n37009), .ZN(
        n37010) );
  OR4_X1 U162 ( .A1(n36996), .A2(n37001), .A3(n37005), .A4(n37010), .ZN(
        OUTA[10]) );
  AOI22_X1 U163 ( .A1(n37702), .A2(\REGISTERS[9][7] ), .B1(n37701), .B2(
        \REGISTERS[16][7] ), .ZN(n37011) );
  AOI22_X1 U164 ( .A1(n37708), .A2(\REGISTERS[23][7] ), .B1(n37710), .B2(
        \REGISTERS[6][7] ), .ZN(n37012) );
  AOI22_X1 U165 ( .A1(n37706), .A2(\REGISTERS[14][7] ), .B1(n37707), .B2(
        \REGISTERS[24][7] ), .ZN(n37013) );
  AOI22_X1 U166 ( .A1(n37704), .A2(\REGISTERS[10][7] ), .B1(n37705), .B2(
        \REGISTERS[12][7] ), .ZN(n37014) );
  NAND4_X1 U167 ( .A1(n37011), .A2(n37012), .A3(n37013), .A4(n37014), .ZN(
        n37015) );
  AOI22_X1 U168 ( .A1(n37723), .A2(\REGISTERS[27][7] ), .B1(n37703), .B2(
        \REGISTERS[1][7] ), .ZN(n37016) );
  AOI22_X1 U169 ( .A1(n37695), .A2(\REGISTERS[21][7] ), .B1(n37699), .B2(
        \REGISTERS[20][7] ), .ZN(n37017) );
  AOI22_X1 U170 ( .A1(n37698), .A2(\REGISTERS[7][7] ), .B1(n37700), .B2(
        \REGISTERS[18][7] ), .ZN(n37018) );
  AOI22_X1 U171 ( .A1(n37716), .A2(\REGISTERS[5][7] ), .B1(n37718), .B2(
        \REGISTERS[28][7] ), .ZN(n37019) );
  NAND4_X1 U172 ( .A1(n37016), .A2(n37017), .A3(n37018), .A4(n37019), .ZN(
        n37020) );
  AOI22_X1 U173 ( .A1(n37709), .A2(\REGISTERS[25][7] ), .B1(n37720), .B2(
        \REGISTERS[11][7] ), .ZN(n37021) );
  AOI22_X1 U174 ( .A1(n37725), .A2(\REGISTERS[31][7] ), .B1(n38278), .B2(
        \REGISTERS[2][7] ), .ZN(n37022) );
  AOI222_X1 U175 ( .A1(n37696), .A2(\REGISTERS[29][7] ), .B1(n37697), .B2(
        \REGISTERS[13][7] ), .C1(n37722), .C2(\REGISTERS[19][7] ), .ZN(n37023)
         );
  NAND3_X1 U176 ( .A1(n37021), .A2(n37022), .A3(n37023), .ZN(n37024) );
  AOI22_X1 U177 ( .A1(n37712), .A2(\REGISTERS[26][7] ), .B1(n37715), .B2(
        \REGISTERS[8][7] ), .ZN(n37025) );
  AOI22_X1 U178 ( .A1(n37714), .A2(\REGISTERS[30][7] ), .B1(n37711), .B2(
        \REGISTERS[3][7] ), .ZN(n37026) );
  AOI22_X1 U179 ( .A1(n37719), .A2(\REGISTERS[17][7] ), .B1(n37717), .B2(
        \REGISTERS[4][7] ), .ZN(n37027) );
  AOI22_X1 U180 ( .A1(n37713), .A2(\REGISTERS[22][7] ), .B1(n37724), .B2(
        \REGISTERS[15][7] ), .ZN(n37028) );
  NAND4_X1 U181 ( .A1(n37025), .A2(n37026), .A3(n37027), .A4(n37028), .ZN(
        n37029) );
  OR4_X1 U182 ( .A1(n37015), .A2(n37020), .A3(n37024), .A4(n37029), .ZN(
        OUTB[7]) );
  AOI22_X1 U183 ( .A1(\REGISTERS[29][7] ), .A2(n37741), .B1(\REGISTERS[30][7] ), .B2(n37742), .ZN(n37030) );
  AOI22_X1 U184 ( .A1(\REGISTERS[4][7] ), .A2(n37743), .B1(\REGISTERS[27][7] ), 
        .B2(n37744), .ZN(n37031) );
  AOI22_X1 U185 ( .A1(\REGISTERS[28][7] ), .A2(n37745), .B1(\REGISTERS[10][7] ), .B2(n37746), .ZN(n37032) );
  AOI22_X1 U186 ( .A1(\REGISTERS[7][7] ), .A2(n37747), .B1(\REGISTERS[6][7] ), 
        .B2(n37748), .ZN(n37033) );
  NAND4_X1 U187 ( .A1(n37030), .A2(n37031), .A3(n37032), .A4(n37033), .ZN(
        n37034) );
  AOI22_X1 U188 ( .A1(\REGISTERS[5][7] ), .A2(n37749), .B1(\REGISTERS[26][7] ), 
        .B2(n37750), .ZN(n37035) );
  AOI22_X1 U189 ( .A1(\REGISTERS[25][7] ), .A2(n37751), .B1(\REGISTERS[21][7] ), .B2(n37752), .ZN(n37036) );
  AOI22_X1 U190 ( .A1(\REGISTERS[17][7] ), .A2(n37753), .B1(\REGISTERS[23][7] ), .B2(n37754), .ZN(n37037) );
  AOI22_X1 U191 ( .A1(\REGISTERS[19][7] ), .A2(n37755), .B1(\REGISTERS[14][7] ), .B2(n37756), .ZN(n37038) );
  NAND4_X1 U192 ( .A1(n37035), .A2(n37036), .A3(n37037), .A4(n37038), .ZN(
        n37039) );
  AOI22_X1 U193 ( .A1(\REGISTERS[16][7] ), .A2(n37726), .B1(\REGISTERS[11][7] ), .B2(n37727), .ZN(n37040) );
  AOI22_X1 U194 ( .A1(\REGISTERS[24][7] ), .A2(n37728), .B1(\REGISTERS[1][7] ), 
        .B2(n37729), .ZN(n37041) );
  AOI222_X1 U195 ( .A1(\REGISTERS[15][7] ), .A2(n37730), .B1(
        \REGISTERS[12][7] ), .B2(n37731), .C1(\REGISTERS[13][7] ), .C2(n38211), 
        .ZN(n37042) );
  NAND3_X1 U196 ( .A1(n37040), .A2(n37041), .A3(n37042), .ZN(n37043) );
  AOI22_X1 U197 ( .A1(\REGISTERS[22][7] ), .A2(n37733), .B1(\REGISTERS[20][7] ), .B2(n37734), .ZN(n37044) );
  AOI22_X1 U198 ( .A1(\REGISTERS[9][7] ), .A2(n37735), .B1(\REGISTERS[18][7] ), 
        .B2(n37736), .ZN(n37045) );
  AOI22_X1 U199 ( .A1(\REGISTERS[31][7] ), .A2(n37737), .B1(\REGISTERS[2][7] ), 
        .B2(n37738), .ZN(n37046) );
  AOI22_X1 U200 ( .A1(\REGISTERS[8][7] ), .A2(n37739), .B1(\REGISTERS[3][7] ), 
        .B2(n37740), .ZN(n37047) );
  NAND4_X1 U201 ( .A1(n37044), .A2(n37045), .A3(n37046), .A4(n37047), .ZN(
        n37048) );
  OR4_X1 U202 ( .A1(n37034), .A2(n37039), .A3(n37043), .A4(n37048), .ZN(
        OUTA[7]) );
  AOI22_X1 U203 ( .A1(n37702), .A2(\REGISTERS[9][6] ), .B1(n37701), .B2(
        \REGISTERS[16][6] ), .ZN(n37049) );
  AOI22_X1 U204 ( .A1(n37708), .A2(\REGISTERS[23][6] ), .B1(n37710), .B2(
        \REGISTERS[6][6] ), .ZN(n37050) );
  AOI22_X1 U205 ( .A1(n37706), .A2(\REGISTERS[14][6] ), .B1(n37707), .B2(
        \REGISTERS[24][6] ), .ZN(n37051) );
  AOI22_X1 U206 ( .A1(n37704), .A2(\REGISTERS[10][6] ), .B1(n37705), .B2(
        \REGISTERS[12][6] ), .ZN(n37052) );
  NAND4_X1 U207 ( .A1(n37049), .A2(n37050), .A3(n37051), .A4(n37052), .ZN(
        n37053) );
  AOI22_X1 U208 ( .A1(n37723), .A2(\REGISTERS[27][6] ), .B1(n37703), .B2(
        \REGISTERS[1][6] ), .ZN(n37054) );
  AOI22_X1 U209 ( .A1(n37695), .A2(\REGISTERS[21][6] ), .B1(n37699), .B2(
        \REGISTERS[20][6] ), .ZN(n37055) );
  AOI22_X1 U210 ( .A1(n37698), .A2(\REGISTERS[7][6] ), .B1(n37700), .B2(
        \REGISTERS[18][6] ), .ZN(n37056) );
  AOI22_X1 U211 ( .A1(n37716), .A2(\REGISTERS[5][6] ), .B1(n37718), .B2(
        \REGISTERS[28][6] ), .ZN(n37057) );
  NAND4_X1 U212 ( .A1(n37054), .A2(n37055), .A3(n37056), .A4(n37057), .ZN(
        n37058) );
  AOI22_X1 U213 ( .A1(n37709), .A2(\REGISTERS[25][6] ), .B1(n37720), .B2(
        \REGISTERS[11][6] ), .ZN(n37059) );
  AOI22_X1 U214 ( .A1(n37725), .A2(\REGISTERS[31][6] ), .B1(n38278), .B2(
        \REGISTERS[2][6] ), .ZN(n37060) );
  AOI222_X1 U215 ( .A1(n37696), .A2(\REGISTERS[29][6] ), .B1(n37697), .B2(
        \REGISTERS[13][6] ), .C1(n37722), .C2(\REGISTERS[19][6] ), .ZN(n37061)
         );
  NAND3_X1 U216 ( .A1(n37059), .A2(n37060), .A3(n37061), .ZN(n37062) );
  AOI22_X1 U217 ( .A1(n37712), .A2(\REGISTERS[26][6] ), .B1(n37715), .B2(
        \REGISTERS[8][6] ), .ZN(n37063) );
  AOI22_X1 U218 ( .A1(n37714), .A2(\REGISTERS[30][6] ), .B1(n37711), .B2(
        \REGISTERS[3][6] ), .ZN(n37064) );
  AOI22_X1 U219 ( .A1(n37719), .A2(\REGISTERS[17][6] ), .B1(n37717), .B2(
        \REGISTERS[4][6] ), .ZN(n37065) );
  AOI22_X1 U220 ( .A1(n37713), .A2(\REGISTERS[22][6] ), .B1(n37724), .B2(
        \REGISTERS[15][6] ), .ZN(n37066) );
  NAND4_X1 U221 ( .A1(n37063), .A2(n37064), .A3(n37065), .A4(n37066), .ZN(
        n37067) );
  OR4_X1 U222 ( .A1(n37053), .A2(n37058), .A3(n37062), .A4(n37067), .ZN(
        OUTB[6]) );
  AOI22_X1 U223 ( .A1(\REGISTERS[29][1] ), .A2(n37741), .B1(\REGISTERS[30][1] ), .B2(n37742), .ZN(n37068) );
  AOI22_X1 U224 ( .A1(\REGISTERS[4][1] ), .A2(n37743), .B1(\REGISTERS[27][1] ), 
        .B2(n37744), .ZN(n37069) );
  AOI22_X1 U225 ( .A1(\REGISTERS[28][1] ), .A2(n37745), .B1(\REGISTERS[10][1] ), .B2(n37746), .ZN(n37070) );
  AOI22_X1 U226 ( .A1(\REGISTERS[7][1] ), .A2(n37747), .B1(\REGISTERS[6][1] ), 
        .B2(n37748), .ZN(n37071) );
  NAND4_X1 U227 ( .A1(n37068), .A2(n37069), .A3(n37070), .A4(n37071), .ZN(
        n37072) );
  AOI22_X1 U228 ( .A1(\REGISTERS[5][1] ), .A2(n37749), .B1(\REGISTERS[26][1] ), 
        .B2(n37750), .ZN(n37073) );
  AOI22_X1 U229 ( .A1(\REGISTERS[25][1] ), .A2(n37751), .B1(\REGISTERS[21][1] ), .B2(n37752), .ZN(n37074) );
  AOI22_X1 U230 ( .A1(\REGISTERS[17][1] ), .A2(n37753), .B1(\REGISTERS[23][1] ), .B2(n37754), .ZN(n37075) );
  AOI22_X1 U231 ( .A1(\REGISTERS[19][1] ), .A2(n37755), .B1(\REGISTERS[14][1] ), .B2(n37756), .ZN(n37076) );
  NAND4_X1 U232 ( .A1(n37073), .A2(n37074), .A3(n37075), .A4(n37076), .ZN(
        n37077) );
  AOI22_X1 U233 ( .A1(\REGISTERS[16][1] ), .A2(n37726), .B1(\REGISTERS[11][1] ), .B2(n37727), .ZN(n37078) );
  AOI22_X1 U234 ( .A1(\REGISTERS[24][1] ), .A2(n37728), .B1(\REGISTERS[1][1] ), 
        .B2(n37729), .ZN(n37079) );
  AOI222_X1 U235 ( .A1(\REGISTERS[15][1] ), .A2(n37730), .B1(
        \REGISTERS[12][1] ), .B2(n37731), .C1(\REGISTERS[13][1] ), .C2(n37732), 
        .ZN(n37080) );
  NAND3_X1 U236 ( .A1(n37078), .A2(n37079), .A3(n37080), .ZN(n37081) );
  AOI22_X1 U237 ( .A1(\REGISTERS[22][1] ), .A2(n37733), .B1(\REGISTERS[20][1] ), .B2(n37734), .ZN(n37082) );
  AOI22_X1 U238 ( .A1(\REGISTERS[9][1] ), .A2(n37735), .B1(\REGISTERS[18][1] ), 
        .B2(n37736), .ZN(n37083) );
  AOI22_X1 U239 ( .A1(\REGISTERS[31][1] ), .A2(n37737), .B1(\REGISTERS[2][1] ), 
        .B2(n37738), .ZN(n37084) );
  AOI22_X1 U240 ( .A1(\REGISTERS[8][1] ), .A2(n37739), .B1(\REGISTERS[3][1] ), 
        .B2(n37740), .ZN(n37085) );
  NAND4_X1 U241 ( .A1(n37082), .A2(n37083), .A3(n37084), .A4(n37085), .ZN(
        n37086) );
  OR4_X1 U242 ( .A1(n37072), .A2(n37077), .A3(n37081), .A4(n37086), .ZN(
        OUTA[1]) );
  AOI22_X1 U243 ( .A1(n37702), .A2(\REGISTERS[9][5] ), .B1(n37701), .B2(
        \REGISTERS[16][5] ), .ZN(n37087) );
  AOI22_X1 U244 ( .A1(n37708), .A2(\REGISTERS[23][5] ), .B1(n37710), .B2(
        \REGISTERS[6][5] ), .ZN(n37088) );
  AOI22_X1 U245 ( .A1(n37706), .A2(\REGISTERS[14][5] ), .B1(n37707), .B2(
        \REGISTERS[24][5] ), .ZN(n37089) );
  AOI22_X1 U246 ( .A1(n37704), .A2(\REGISTERS[10][5] ), .B1(n37705), .B2(
        \REGISTERS[12][5] ), .ZN(n37090) );
  NAND4_X1 U247 ( .A1(n37087), .A2(n37088), .A3(n37089), .A4(n37090), .ZN(
        n37091) );
  AOI22_X1 U248 ( .A1(n37723), .A2(\REGISTERS[27][5] ), .B1(n37703), .B2(
        \REGISTERS[1][5] ), .ZN(n37092) );
  AOI22_X1 U249 ( .A1(n37695), .A2(\REGISTERS[21][5] ), .B1(n37699), .B2(
        \REGISTERS[20][5] ), .ZN(n37093) );
  AOI22_X1 U250 ( .A1(n37698), .A2(\REGISTERS[7][5] ), .B1(n37700), .B2(
        \REGISTERS[18][5] ), .ZN(n37094) );
  AOI22_X1 U251 ( .A1(n37716), .A2(\REGISTERS[5][5] ), .B1(n37718), .B2(
        \REGISTERS[28][5] ), .ZN(n37095) );
  NAND4_X1 U252 ( .A1(n37092), .A2(n37093), .A3(n37094), .A4(n37095), .ZN(
        n37096) );
  AOI22_X1 U253 ( .A1(n37709), .A2(\REGISTERS[25][5] ), .B1(n37720), .B2(
        \REGISTERS[11][5] ), .ZN(n37097) );
  AOI22_X1 U254 ( .A1(n37725), .A2(\REGISTERS[31][5] ), .B1(n38278), .B2(
        \REGISTERS[2][5] ), .ZN(n37098) );
  AOI222_X1 U255 ( .A1(n37696), .A2(\REGISTERS[29][5] ), .B1(n37697), .B2(
        \REGISTERS[13][5] ), .C1(n37722), .C2(\REGISTERS[19][5] ), .ZN(n37099)
         );
  NAND3_X1 U256 ( .A1(n37097), .A2(n37098), .A3(n37099), .ZN(n37100) );
  AOI22_X1 U257 ( .A1(n37712), .A2(\REGISTERS[26][5] ), .B1(n37715), .B2(
        \REGISTERS[8][5] ), .ZN(n37101) );
  AOI22_X1 U258 ( .A1(n37714), .A2(\REGISTERS[30][5] ), .B1(n37711), .B2(
        \REGISTERS[3][5] ), .ZN(n37102) );
  AOI22_X1 U259 ( .A1(n37719), .A2(\REGISTERS[17][5] ), .B1(n37717), .B2(
        \REGISTERS[4][5] ), .ZN(n37103) );
  AOI22_X1 U260 ( .A1(n37713), .A2(\REGISTERS[22][5] ), .B1(n37724), .B2(
        \REGISTERS[15][5] ), .ZN(n37104) );
  NAND4_X1 U261 ( .A1(n37101), .A2(n37102), .A3(n37103), .A4(n37104), .ZN(
        n37105) );
  OR4_X1 U262 ( .A1(n37091), .A2(n37096), .A3(n37100), .A4(n37105), .ZN(
        OUTB[5]) );
  AOI22_X1 U263 ( .A1(n37741), .A2(\REGISTERS[29][0] ), .B1(n37742), .B2(
        \REGISTERS[30][0] ), .ZN(n37106) );
  AOI22_X1 U264 ( .A1(n37743), .A2(\REGISTERS[4][0] ), .B1(n37744), .B2(
        \REGISTERS[27][0] ), .ZN(n37107) );
  AOI22_X1 U265 ( .A1(n37745), .A2(\REGISTERS[28][0] ), .B1(n37746), .B2(
        \REGISTERS[10][0] ), .ZN(n37108) );
  AOI22_X1 U266 ( .A1(n37747), .A2(\REGISTERS[7][0] ), .B1(n37748), .B2(
        \REGISTERS[6][0] ), .ZN(n37109) );
  NAND4_X1 U267 ( .A1(n37106), .A2(n37107), .A3(n37108), .A4(n37109), .ZN(
        n37110) );
  AOI22_X1 U268 ( .A1(n37749), .A2(\REGISTERS[5][0] ), .B1(n37750), .B2(
        \REGISTERS[26][0] ), .ZN(n37111) );
  AOI22_X1 U269 ( .A1(n37751), .A2(\REGISTERS[25][0] ), .B1(n37752), .B2(
        \REGISTERS[21][0] ), .ZN(n37112) );
  AOI22_X1 U270 ( .A1(n37753), .A2(\REGISTERS[17][0] ), .B1(n37754), .B2(
        \REGISTERS[23][0] ), .ZN(n37113) );
  AOI22_X1 U271 ( .A1(n37755), .A2(\REGISTERS[19][0] ), .B1(n37756), .B2(
        \REGISTERS[14][0] ), .ZN(n37114) );
  NAND4_X1 U272 ( .A1(n37111), .A2(n37112), .A3(n37113), .A4(n37114), .ZN(
        n37115) );
  AOI22_X1 U273 ( .A1(n37726), .A2(\REGISTERS[16][0] ), .B1(n37727), .B2(
        \REGISTERS[11][0] ), .ZN(n37116) );
  AOI22_X1 U274 ( .A1(n37728), .A2(\REGISTERS[24][0] ), .B1(n37729), .B2(
        \REGISTERS[1][0] ), .ZN(n37117) );
  AOI222_X1 U275 ( .A1(n37730), .A2(\REGISTERS[15][0] ), .B1(n37731), .B2(
        \REGISTERS[12][0] ), .C1(n37732), .C2(\REGISTERS[13][0] ), .ZN(n37118)
         );
  NAND3_X1 U276 ( .A1(n37116), .A2(n37117), .A3(n37118), .ZN(n37119) );
  AOI22_X1 U277 ( .A1(n37733), .A2(\REGISTERS[22][0] ), .B1(n37734), .B2(
        \REGISTERS[20][0] ), .ZN(n37120) );
  AOI22_X1 U278 ( .A1(n37735), .A2(\REGISTERS[9][0] ), .B1(n37736), .B2(
        \REGISTERS[18][0] ), .ZN(n37121) );
  AOI22_X1 U279 ( .A1(n37737), .A2(\REGISTERS[31][0] ), .B1(n37738), .B2(
        \REGISTERS[2][0] ), .ZN(n37122) );
  AOI22_X1 U280 ( .A1(n37739), .A2(\REGISTERS[8][0] ), .B1(n37740), .B2(
        \REGISTERS[3][0] ), .ZN(n37123) );
  NAND4_X1 U281 ( .A1(n37120), .A2(n37121), .A3(n37122), .A4(n37123), .ZN(
        n37124) );
  OR4_X1 U282 ( .A1(n37110), .A2(n37115), .A3(n37119), .A4(n37124), .ZN(
        OUTA[0]) );
  AOI22_X1 U283 ( .A1(n37702), .A2(\REGISTERS[9][31] ), .B1(n37701), .B2(
        \REGISTERS[16][31] ), .ZN(n37125) );
  AOI22_X1 U284 ( .A1(n37708), .A2(\REGISTERS[23][31] ), .B1(n37710), .B2(
        \REGISTERS[6][31] ), .ZN(n37126) );
  AOI22_X1 U285 ( .A1(n37706), .A2(\REGISTERS[14][31] ), .B1(n37707), .B2(
        \REGISTERS[24][31] ), .ZN(n37127) );
  AOI22_X1 U286 ( .A1(n37704), .A2(\REGISTERS[10][31] ), .B1(n37705), .B2(
        \REGISTERS[12][31] ), .ZN(n37128) );
  NAND4_X1 U287 ( .A1(n37125), .A2(n37126), .A3(n37127), .A4(n37128), .ZN(
        n37129) );
  AOI22_X1 U288 ( .A1(n37723), .A2(\REGISTERS[27][31] ), .B1(n37703), .B2(
        \REGISTERS[1][31] ), .ZN(n37130) );
  AOI22_X1 U289 ( .A1(n37695), .A2(\REGISTERS[21][31] ), .B1(n37699), .B2(
        \REGISTERS[20][31] ), .ZN(n37131) );
  AOI22_X1 U290 ( .A1(n37698), .A2(\REGISTERS[7][31] ), .B1(n37700), .B2(
        \REGISTERS[18][31] ), .ZN(n37132) );
  AOI22_X1 U291 ( .A1(n37716), .A2(\REGISTERS[5][31] ), .B1(n37718), .B2(
        \REGISTERS[28][31] ), .ZN(n37133) );
  NAND4_X1 U292 ( .A1(n37130), .A2(n37131), .A3(n37132), .A4(n37133), .ZN(
        n37134) );
  AOI22_X1 U293 ( .A1(n37709), .A2(\REGISTERS[25][31] ), .B1(n37720), .B2(
        \REGISTERS[11][31] ), .ZN(n37135) );
  AOI22_X1 U294 ( .A1(n38277), .A2(\REGISTERS[31][31] ), .B1(n37721), .B2(
        \REGISTERS[2][31] ), .ZN(n37136) );
  AOI222_X1 U295 ( .A1(n37696), .A2(\REGISTERS[29][31] ), .B1(n37697), .B2(
        \REGISTERS[13][31] ), .C1(n37722), .C2(\REGISTERS[19][31] ), .ZN(
        n37137) );
  NAND3_X1 U296 ( .A1(n37135), .A2(n37136), .A3(n37137), .ZN(n37138) );
  AOI22_X1 U297 ( .A1(n37712), .A2(\REGISTERS[26][31] ), .B1(n37715), .B2(
        \REGISTERS[8][31] ), .ZN(n37139) );
  AOI22_X1 U298 ( .A1(n37714), .A2(\REGISTERS[30][31] ), .B1(n37711), .B2(
        \REGISTERS[3][31] ), .ZN(n37140) );
  AOI22_X1 U299 ( .A1(n37719), .A2(\REGISTERS[17][31] ), .B1(n37717), .B2(
        \REGISTERS[4][31] ), .ZN(n37141) );
  AOI22_X1 U300 ( .A1(n37713), .A2(\REGISTERS[22][31] ), .B1(n38289), .B2(
        \REGISTERS[15][31] ), .ZN(n37142) );
  NAND4_X1 U301 ( .A1(n37139), .A2(n37140), .A3(n37141), .A4(n37142), .ZN(
        n37143) );
  OR4_X1 U302 ( .A1(n37129), .A2(n37134), .A3(n37138), .A4(n37143), .ZN(
        OUTB[31]) );
  AOI22_X1 U303 ( .A1(n37702), .A2(\REGISTERS[9][4] ), .B1(n37701), .B2(
        \REGISTERS[16][4] ), .ZN(n37144) );
  AOI22_X1 U304 ( .A1(n37708), .A2(\REGISTERS[23][4] ), .B1(n37710), .B2(
        \REGISTERS[6][4] ), .ZN(n37145) );
  AOI22_X1 U305 ( .A1(n37706), .A2(\REGISTERS[14][4] ), .B1(n37707), .B2(
        \REGISTERS[24][4] ), .ZN(n37146) );
  AOI22_X1 U306 ( .A1(n37704), .A2(\REGISTERS[10][4] ), .B1(n37705), .B2(
        \REGISTERS[12][4] ), .ZN(n37147) );
  NAND4_X1 U307 ( .A1(n37144), .A2(n37145), .A3(n37146), .A4(n37147), .ZN(
        n37148) );
  AOI22_X1 U308 ( .A1(n37723), .A2(\REGISTERS[27][4] ), .B1(n37703), .B2(
        \REGISTERS[1][4] ), .ZN(n37149) );
  AOI22_X1 U309 ( .A1(n37695), .A2(\REGISTERS[21][4] ), .B1(n37699), .B2(
        \REGISTERS[20][4] ), .ZN(n37150) );
  AOI22_X1 U310 ( .A1(n37698), .A2(\REGISTERS[7][4] ), .B1(n37700), .B2(
        \REGISTERS[18][4] ), .ZN(n37151) );
  AOI22_X1 U311 ( .A1(n37716), .A2(\REGISTERS[5][4] ), .B1(n37718), .B2(
        \REGISTERS[28][4] ), .ZN(n37152) );
  NAND4_X1 U312 ( .A1(n37149), .A2(n37150), .A3(n37151), .A4(n37152), .ZN(
        n37153) );
  AOI22_X1 U313 ( .A1(n37709), .A2(\REGISTERS[25][4] ), .B1(n37720), .B2(
        \REGISTERS[11][4] ), .ZN(n37154) );
  AOI22_X1 U314 ( .A1(n37725), .A2(\REGISTERS[31][4] ), .B1(n38278), .B2(
        \REGISTERS[2][4] ), .ZN(n37155) );
  AOI222_X1 U315 ( .A1(n37696), .A2(\REGISTERS[29][4] ), .B1(n37697), .B2(
        \REGISTERS[13][4] ), .C1(n37722), .C2(\REGISTERS[19][4] ), .ZN(n37156)
         );
  NAND3_X1 U316 ( .A1(n37154), .A2(n37155), .A3(n37156), .ZN(n37157) );
  AOI22_X1 U317 ( .A1(n37712), .A2(\REGISTERS[26][4] ), .B1(n37715), .B2(
        \REGISTERS[8][4] ), .ZN(n37158) );
  AOI22_X1 U318 ( .A1(n37714), .A2(\REGISTERS[30][4] ), .B1(n37711), .B2(
        \REGISTERS[3][4] ), .ZN(n37159) );
  AOI22_X1 U319 ( .A1(n37719), .A2(\REGISTERS[17][4] ), .B1(n37717), .B2(
        \REGISTERS[4][4] ), .ZN(n37160) );
  AOI22_X1 U320 ( .A1(n37713), .A2(\REGISTERS[22][4] ), .B1(n37724), .B2(
        \REGISTERS[15][4] ), .ZN(n37161) );
  NAND4_X1 U321 ( .A1(n37158), .A2(n37159), .A3(n37160), .A4(n37161), .ZN(
        n37162) );
  OR4_X1 U322 ( .A1(n37148), .A2(n37153), .A3(n37157), .A4(n37162), .ZN(
        OUTB[4]) );
  AOI22_X1 U323 ( .A1(\REGISTERS[29][4] ), .A2(n38228), .B1(\REGISTERS[30][4] ), .B2(n38229), .ZN(n37163) );
  AOI22_X1 U324 ( .A1(\REGISTERS[4][4] ), .A2(n38230), .B1(\REGISTERS[27][4] ), 
        .B2(n38231), .ZN(n37164) );
  AOI22_X1 U325 ( .A1(\REGISTERS[28][4] ), .A2(n38232), .B1(\REGISTERS[10][4] ), .B2(n38233), .ZN(n37165) );
  AOI22_X1 U326 ( .A1(\REGISTERS[7][4] ), .A2(n38234), .B1(\REGISTERS[6][4] ), 
        .B2(n38235), .ZN(n37166) );
  NAND4_X1 U327 ( .A1(n37163), .A2(n37164), .A3(n37165), .A4(n37166), .ZN(
        n37167) );
  AOI22_X1 U328 ( .A1(\REGISTERS[5][4] ), .A2(n38240), .B1(\REGISTERS[26][4] ), 
        .B2(n38241), .ZN(n37168) );
  AOI22_X1 U329 ( .A1(\REGISTERS[25][4] ), .A2(n38242), .B1(\REGISTERS[21][4] ), .B2(n38243), .ZN(n37169) );
  AOI22_X1 U330 ( .A1(\REGISTERS[17][4] ), .A2(n38244), .B1(\REGISTERS[23][4] ), .B2(n38245), .ZN(n37170) );
  AOI22_X1 U331 ( .A1(\REGISTERS[19][4] ), .A2(n38246), .B1(\REGISTERS[14][4] ), .B2(n38247), .ZN(n37171) );
  NAND4_X1 U332 ( .A1(n37168), .A2(n37169), .A3(n37170), .A4(n37171), .ZN(
        n37172) );
  AOI22_X1 U333 ( .A1(\REGISTERS[16][4] ), .A2(n38205), .B1(\REGISTERS[11][4] ), .B2(n38206), .ZN(n37173) );
  AOI22_X1 U334 ( .A1(\REGISTERS[24][4] ), .A2(n38207), .B1(\REGISTERS[1][4] ), 
        .B2(n38208), .ZN(n37174) );
  AOI222_X1 U335 ( .A1(\REGISTERS[15][4] ), .A2(n38209), .B1(
        \REGISTERS[12][4] ), .B2(n38210), .C1(\REGISTERS[13][4] ), .C2(n38211), 
        .ZN(n37175) );
  NAND3_X1 U336 ( .A1(n37173), .A2(n37174), .A3(n37175), .ZN(n37176) );
  AOI22_X1 U337 ( .A1(\REGISTERS[22][4] ), .A2(n38216), .B1(\REGISTERS[20][4] ), .B2(n38217), .ZN(n37177) );
  AOI22_X1 U338 ( .A1(\REGISTERS[9][4] ), .A2(n38218), .B1(\REGISTERS[18][4] ), 
        .B2(n38219), .ZN(n37178) );
  AOI22_X1 U339 ( .A1(\REGISTERS[31][4] ), .A2(n38220), .B1(\REGISTERS[2][4] ), 
        .B2(n38221), .ZN(n37179) );
  AOI22_X1 U340 ( .A1(\REGISTERS[8][4] ), .A2(n38222), .B1(\REGISTERS[3][4] ), 
        .B2(n38223), .ZN(n37180) );
  NAND4_X1 U341 ( .A1(n37177), .A2(n37178), .A3(n37179), .A4(n37180), .ZN(
        n37181) );
  OR4_X1 U342 ( .A1(n37167), .A2(n37172), .A3(n37176), .A4(n37181), .ZN(
        OUTA[4]) );
  AOI22_X1 U343 ( .A1(n37702), .A2(\REGISTERS[9][30] ), .B1(n37701), .B2(
        \REGISTERS[16][30] ), .ZN(n37182) );
  AOI22_X1 U344 ( .A1(n37708), .A2(\REGISTERS[23][30] ), .B1(n37710), .B2(
        \REGISTERS[6][30] ), .ZN(n37183) );
  AOI22_X1 U345 ( .A1(n37706), .A2(\REGISTERS[14][30] ), .B1(n37707), .B2(
        \REGISTERS[24][30] ), .ZN(n37184) );
  AOI22_X1 U346 ( .A1(n37704), .A2(\REGISTERS[10][30] ), .B1(n37705), .B2(
        \REGISTERS[12][30] ), .ZN(n37185) );
  NAND4_X1 U347 ( .A1(n37182), .A2(n37183), .A3(n37184), .A4(n37185), .ZN(
        n37186) );
  AOI22_X1 U348 ( .A1(n37723), .A2(\REGISTERS[27][30] ), .B1(n37703), .B2(
        \REGISTERS[1][30] ), .ZN(n37187) );
  AOI22_X1 U349 ( .A1(n37695), .A2(\REGISTERS[21][30] ), .B1(n37699), .B2(
        \REGISTERS[20][30] ), .ZN(n37188) );
  AOI22_X1 U350 ( .A1(n37698), .A2(\REGISTERS[7][30] ), .B1(n37700), .B2(
        \REGISTERS[18][30] ), .ZN(n37189) );
  AOI22_X1 U351 ( .A1(n37716), .A2(\REGISTERS[5][30] ), .B1(n37718), .B2(
        \REGISTERS[28][30] ), .ZN(n37190) );
  NAND4_X1 U352 ( .A1(n37187), .A2(n37188), .A3(n37189), .A4(n37190), .ZN(
        n37191) );
  AOI22_X1 U353 ( .A1(n37709), .A2(\REGISTERS[25][30] ), .B1(n37720), .B2(
        \REGISTERS[11][30] ), .ZN(n37192) );
  AOI22_X1 U354 ( .A1(n37725), .A2(\REGISTERS[31][30] ), .B1(n37721), .B2(
        \REGISTERS[2][30] ), .ZN(n37193) );
  AOI222_X1 U355 ( .A1(n37696), .A2(\REGISTERS[29][30] ), .B1(n37697), .B2(
        \REGISTERS[13][30] ), .C1(n37722), .C2(\REGISTERS[19][30] ), .ZN(
        n37194) );
  NAND3_X1 U356 ( .A1(n37192), .A2(n37193), .A3(n37194), .ZN(n37195) );
  AOI22_X1 U357 ( .A1(n37712), .A2(\REGISTERS[26][30] ), .B1(n37715), .B2(
        \REGISTERS[8][30] ), .ZN(n37196) );
  AOI22_X1 U358 ( .A1(n37714), .A2(\REGISTERS[30][30] ), .B1(n37711), .B2(
        \REGISTERS[3][30] ), .ZN(n37197) );
  AOI22_X1 U359 ( .A1(n37719), .A2(\REGISTERS[17][30] ), .B1(n37717), .B2(
        \REGISTERS[4][30] ), .ZN(n37198) );
  AOI22_X1 U360 ( .A1(n37713), .A2(\REGISTERS[22][30] ), .B1(n37724), .B2(
        \REGISTERS[15][30] ), .ZN(n37199) );
  NAND4_X1 U361 ( .A1(n37196), .A2(n37197), .A3(n37198), .A4(n37199), .ZN(
        n37200) );
  OR4_X1 U362 ( .A1(n37186), .A2(n37191), .A3(n37195), .A4(n37200), .ZN(
        OUTB[30]) );
  AOI22_X1 U363 ( .A1(n37702), .A2(\REGISTERS[9][29] ), .B1(n37701), .B2(
        \REGISTERS[16][29] ), .ZN(n37201) );
  AOI22_X1 U364 ( .A1(n37708), .A2(\REGISTERS[23][29] ), .B1(n37710), .B2(
        \REGISTERS[6][29] ), .ZN(n37202) );
  AOI22_X1 U365 ( .A1(n37706), .A2(\REGISTERS[14][29] ), .B1(n37707), .B2(
        \REGISTERS[24][29] ), .ZN(n37203) );
  AOI22_X1 U366 ( .A1(n37704), .A2(\REGISTERS[10][29] ), .B1(n37705), .B2(
        \REGISTERS[12][29] ), .ZN(n37204) );
  NAND4_X1 U367 ( .A1(n37201), .A2(n37202), .A3(n37203), .A4(n37204), .ZN(
        n37205) );
  AOI22_X1 U368 ( .A1(n37723), .A2(\REGISTERS[27][29] ), .B1(n37703), .B2(
        \REGISTERS[1][29] ), .ZN(n37206) );
  AOI22_X1 U369 ( .A1(n37695), .A2(\REGISTERS[21][29] ), .B1(n37699), .B2(
        \REGISTERS[20][29] ), .ZN(n37207) );
  AOI22_X1 U370 ( .A1(n37698), .A2(\REGISTERS[7][29] ), .B1(n37700), .B2(
        \REGISTERS[18][29] ), .ZN(n37208) );
  AOI22_X1 U371 ( .A1(n37716), .A2(\REGISTERS[5][29] ), .B1(n37718), .B2(
        \REGISTERS[28][29] ), .ZN(n37209) );
  NAND4_X1 U372 ( .A1(n37206), .A2(n37207), .A3(n37208), .A4(n37209), .ZN(
        n37210) );
  AOI22_X1 U373 ( .A1(n37709), .A2(\REGISTERS[25][29] ), .B1(n37720), .B2(
        \REGISTERS[11][29] ), .ZN(n37211) );
  AOI22_X1 U374 ( .A1(n37725), .A2(\REGISTERS[31][29] ), .B1(n37721), .B2(
        \REGISTERS[2][29] ), .ZN(n37212) );
  AOI222_X1 U375 ( .A1(n37696), .A2(\REGISTERS[29][29] ), .B1(n37697), .B2(
        \REGISTERS[13][29] ), .C1(n37722), .C2(\REGISTERS[19][29] ), .ZN(
        n37213) );
  NAND3_X1 U376 ( .A1(n37211), .A2(n37212), .A3(n37213), .ZN(n37214) );
  AOI22_X1 U377 ( .A1(n37712), .A2(\REGISTERS[26][29] ), .B1(n37715), .B2(
        \REGISTERS[8][29] ), .ZN(n37215) );
  AOI22_X1 U378 ( .A1(n37714), .A2(\REGISTERS[30][29] ), .B1(n37711), .B2(
        \REGISTERS[3][29] ), .ZN(n37216) );
  AOI22_X1 U379 ( .A1(n37719), .A2(\REGISTERS[17][29] ), .B1(n37717), .B2(
        \REGISTERS[4][29] ), .ZN(n37217) );
  AOI22_X1 U380 ( .A1(n37713), .A2(\REGISTERS[22][29] ), .B1(n37724), .B2(
        \REGISTERS[15][29] ), .ZN(n37218) );
  NAND4_X1 U381 ( .A1(n37215), .A2(n37216), .A3(n37217), .A4(n37218), .ZN(
        n37219) );
  OR4_X1 U382 ( .A1(n37205), .A2(n37210), .A3(n37214), .A4(n37219), .ZN(
        OUTB[29]) );
  AOI22_X1 U383 ( .A1(n37702), .A2(\REGISTERS[9][28] ), .B1(n37701), .B2(
        \REGISTERS[16][28] ), .ZN(n37220) );
  AOI22_X1 U384 ( .A1(n37708), .A2(\REGISTERS[23][28] ), .B1(n37710), .B2(
        \REGISTERS[6][28] ), .ZN(n37221) );
  AOI22_X1 U385 ( .A1(n37706), .A2(\REGISTERS[14][28] ), .B1(n37707), .B2(
        \REGISTERS[24][28] ), .ZN(n37222) );
  AOI22_X1 U386 ( .A1(n37704), .A2(\REGISTERS[10][28] ), .B1(n37705), .B2(
        \REGISTERS[12][28] ), .ZN(n37223) );
  NAND4_X1 U387 ( .A1(n37220), .A2(n37221), .A3(n37222), .A4(n37223), .ZN(
        n37224) );
  AOI22_X1 U388 ( .A1(n37723), .A2(\REGISTERS[27][28] ), .B1(n37703), .B2(
        \REGISTERS[1][28] ), .ZN(n37225) );
  AOI22_X1 U389 ( .A1(n37695), .A2(\REGISTERS[21][28] ), .B1(n37699), .B2(
        \REGISTERS[20][28] ), .ZN(n37226) );
  AOI22_X1 U390 ( .A1(n37698), .A2(\REGISTERS[7][28] ), .B1(n37700), .B2(
        \REGISTERS[18][28] ), .ZN(n37227) );
  AOI22_X1 U391 ( .A1(n37716), .A2(\REGISTERS[5][28] ), .B1(n37718), .B2(
        \REGISTERS[28][28] ), .ZN(n37228) );
  NAND4_X1 U392 ( .A1(n37225), .A2(n37226), .A3(n37227), .A4(n37228), .ZN(
        n37229) );
  AOI22_X1 U393 ( .A1(n37709), .A2(\REGISTERS[25][28] ), .B1(n37720), .B2(
        \REGISTERS[11][28] ), .ZN(n37230) );
  AOI22_X1 U394 ( .A1(n37725), .A2(\REGISTERS[31][28] ), .B1(n37721), .B2(
        \REGISTERS[2][28] ), .ZN(n37231) );
  AOI222_X1 U395 ( .A1(n37696), .A2(\REGISTERS[29][28] ), .B1(n37697), .B2(
        \REGISTERS[13][28] ), .C1(n37722), .C2(\REGISTERS[19][28] ), .ZN(
        n37232) );
  NAND3_X1 U396 ( .A1(n37230), .A2(n37231), .A3(n37232), .ZN(n37233) );
  AOI22_X1 U397 ( .A1(n37712), .A2(\REGISTERS[26][28] ), .B1(n37715), .B2(
        \REGISTERS[8][28] ), .ZN(n37234) );
  AOI22_X1 U398 ( .A1(n37714), .A2(\REGISTERS[30][28] ), .B1(n37711), .B2(
        \REGISTERS[3][28] ), .ZN(n37235) );
  AOI22_X1 U399 ( .A1(n37719), .A2(\REGISTERS[17][28] ), .B1(n37717), .B2(
        \REGISTERS[4][28] ), .ZN(n37236) );
  AOI22_X1 U400 ( .A1(n37713), .A2(\REGISTERS[22][28] ), .B1(n37724), .B2(
        \REGISTERS[15][28] ), .ZN(n37237) );
  NAND4_X1 U401 ( .A1(n37234), .A2(n37235), .A3(n37236), .A4(n37237), .ZN(
        n37238) );
  OR4_X1 U402 ( .A1(n37224), .A2(n37229), .A3(n37233), .A4(n37238), .ZN(
        OUTB[28]) );
  AOI22_X1 U403 ( .A1(n37702), .A2(\REGISTERS[9][27] ), .B1(n37701), .B2(
        \REGISTERS[16][27] ), .ZN(n37239) );
  AOI22_X1 U404 ( .A1(n37708), .A2(\REGISTERS[23][27] ), .B1(n37710), .B2(
        \REGISTERS[6][27] ), .ZN(n37240) );
  AOI22_X1 U405 ( .A1(n37706), .A2(\REGISTERS[14][27] ), .B1(n37707), .B2(
        \REGISTERS[24][27] ), .ZN(n37241) );
  AOI22_X1 U406 ( .A1(n37704), .A2(\REGISTERS[10][27] ), .B1(n37705), .B2(
        \REGISTERS[12][27] ), .ZN(n37242) );
  NAND4_X1 U407 ( .A1(n37239), .A2(n37240), .A3(n37241), .A4(n37242), .ZN(
        n37243) );
  AOI22_X1 U408 ( .A1(n37723), .A2(\REGISTERS[27][27] ), .B1(n37703), .B2(
        \REGISTERS[1][27] ), .ZN(n37244) );
  AOI22_X1 U409 ( .A1(n37695), .A2(\REGISTERS[21][27] ), .B1(n37699), .B2(
        \REGISTERS[20][27] ), .ZN(n37245) );
  AOI22_X1 U410 ( .A1(n37698), .A2(\REGISTERS[7][27] ), .B1(n37700), .B2(
        \REGISTERS[18][27] ), .ZN(n37246) );
  AOI22_X1 U411 ( .A1(n37716), .A2(\REGISTERS[5][27] ), .B1(n37718), .B2(
        \REGISTERS[28][27] ), .ZN(n37247) );
  NAND4_X1 U412 ( .A1(n37244), .A2(n37245), .A3(n37246), .A4(n37247), .ZN(
        n37248) );
  AOI22_X1 U413 ( .A1(n37709), .A2(\REGISTERS[25][27] ), .B1(n37720), .B2(
        \REGISTERS[11][27] ), .ZN(n37249) );
  AOI22_X1 U414 ( .A1(n37725), .A2(\REGISTERS[31][27] ), .B1(n37721), .B2(
        \REGISTERS[2][27] ), .ZN(n37250) );
  AOI222_X1 U415 ( .A1(n37696), .A2(\REGISTERS[29][27] ), .B1(n37697), .B2(
        \REGISTERS[13][27] ), .C1(n37722), .C2(\REGISTERS[19][27] ), .ZN(
        n37251) );
  NAND3_X1 U416 ( .A1(n37249), .A2(n37250), .A3(n37251), .ZN(n37252) );
  AOI22_X1 U417 ( .A1(n37712), .A2(\REGISTERS[26][27] ), .B1(n37715), .B2(
        \REGISTERS[8][27] ), .ZN(n37253) );
  AOI22_X1 U418 ( .A1(n37714), .A2(\REGISTERS[30][27] ), .B1(n37711), .B2(
        \REGISTERS[3][27] ), .ZN(n37254) );
  AOI22_X1 U419 ( .A1(n37719), .A2(\REGISTERS[17][27] ), .B1(n37717), .B2(
        \REGISTERS[4][27] ), .ZN(n37255) );
  AOI22_X1 U420 ( .A1(n37713), .A2(\REGISTERS[22][27] ), .B1(n37724), .B2(
        \REGISTERS[15][27] ), .ZN(n37256) );
  NAND4_X1 U421 ( .A1(n37253), .A2(n37254), .A3(n37255), .A4(n37256), .ZN(
        n37257) );
  OR4_X1 U422 ( .A1(n37243), .A2(n37248), .A3(n37252), .A4(n37257), .ZN(
        OUTB[27]) );
  AOI22_X1 U423 ( .A1(n37702), .A2(\REGISTERS[9][26] ), .B1(n37701), .B2(
        \REGISTERS[16][26] ), .ZN(n37258) );
  AOI22_X1 U424 ( .A1(n37708), .A2(\REGISTERS[23][26] ), .B1(n37710), .B2(
        \REGISTERS[6][26] ), .ZN(n37259) );
  AOI22_X1 U425 ( .A1(n37706), .A2(\REGISTERS[14][26] ), .B1(n37707), .B2(
        \REGISTERS[24][26] ), .ZN(n37260) );
  AOI22_X1 U426 ( .A1(n37704), .A2(\REGISTERS[10][26] ), .B1(n37705), .B2(
        \REGISTERS[12][26] ), .ZN(n37261) );
  NAND4_X1 U427 ( .A1(n37258), .A2(n37259), .A3(n37260), .A4(n37261), .ZN(
        n37262) );
  AOI22_X1 U428 ( .A1(n37723), .A2(\REGISTERS[27][26] ), .B1(n37703), .B2(
        \REGISTERS[1][26] ), .ZN(n37263) );
  AOI22_X1 U429 ( .A1(n37695), .A2(\REGISTERS[21][26] ), .B1(n37699), .B2(
        \REGISTERS[20][26] ), .ZN(n37264) );
  AOI22_X1 U430 ( .A1(n37698), .A2(\REGISTERS[7][26] ), .B1(n37700), .B2(
        \REGISTERS[18][26] ), .ZN(n37265) );
  AOI22_X1 U431 ( .A1(n37716), .A2(\REGISTERS[5][26] ), .B1(n37718), .B2(
        \REGISTERS[28][26] ), .ZN(n37266) );
  NAND4_X1 U432 ( .A1(n37263), .A2(n37264), .A3(n37265), .A4(n37266), .ZN(
        n37267) );
  AOI22_X1 U433 ( .A1(n37709), .A2(\REGISTERS[25][26] ), .B1(n37720), .B2(
        \REGISTERS[11][26] ), .ZN(n37268) );
  AOI22_X1 U434 ( .A1(n37725), .A2(\REGISTERS[31][26] ), .B1(n37721), .B2(
        \REGISTERS[2][26] ), .ZN(n37269) );
  AOI222_X1 U435 ( .A1(n37696), .A2(\REGISTERS[29][26] ), .B1(n37697), .B2(
        \REGISTERS[13][26] ), .C1(n37722), .C2(\REGISTERS[19][26] ), .ZN(
        n37270) );
  NAND3_X1 U436 ( .A1(n37268), .A2(n37269), .A3(n37270), .ZN(n37271) );
  AOI22_X1 U437 ( .A1(n37712), .A2(\REGISTERS[26][26] ), .B1(n37715), .B2(
        \REGISTERS[8][26] ), .ZN(n37272) );
  AOI22_X1 U438 ( .A1(n37714), .A2(\REGISTERS[30][26] ), .B1(n37711), .B2(
        \REGISTERS[3][26] ), .ZN(n37273) );
  AOI22_X1 U439 ( .A1(n37719), .A2(\REGISTERS[17][26] ), .B1(n37717), .B2(
        \REGISTERS[4][26] ), .ZN(n37274) );
  AOI22_X1 U440 ( .A1(n37713), .A2(\REGISTERS[22][26] ), .B1(n37724), .B2(
        \REGISTERS[15][26] ), .ZN(n37275) );
  NAND4_X1 U441 ( .A1(n37272), .A2(n37273), .A3(n37274), .A4(n37275), .ZN(
        n37276) );
  OR4_X1 U442 ( .A1(n37262), .A2(n37267), .A3(n37271), .A4(n37276), .ZN(
        OUTB[26]) );
  AOI22_X1 U443 ( .A1(n37702), .A2(\REGISTERS[9][25] ), .B1(n37701), .B2(
        \REGISTERS[16][25] ), .ZN(n37277) );
  AOI22_X1 U444 ( .A1(n37708), .A2(\REGISTERS[23][25] ), .B1(n37710), .B2(
        \REGISTERS[6][25] ), .ZN(n37278) );
  AOI22_X1 U445 ( .A1(n37706), .A2(\REGISTERS[14][25] ), .B1(n37707), .B2(
        \REGISTERS[24][25] ), .ZN(n37279) );
  AOI22_X1 U446 ( .A1(n37704), .A2(\REGISTERS[10][25] ), .B1(n37705), .B2(
        \REGISTERS[12][25] ), .ZN(n37280) );
  NAND4_X1 U447 ( .A1(n37277), .A2(n37278), .A3(n37279), .A4(n37280), .ZN(
        n37281) );
  AOI22_X1 U448 ( .A1(n37723), .A2(\REGISTERS[27][25] ), .B1(n37703), .B2(
        \REGISTERS[1][25] ), .ZN(n37282) );
  AOI22_X1 U449 ( .A1(n37695), .A2(\REGISTERS[21][25] ), .B1(n37699), .B2(
        \REGISTERS[20][25] ), .ZN(n37283) );
  AOI22_X1 U450 ( .A1(n37698), .A2(\REGISTERS[7][25] ), .B1(n37700), .B2(
        \REGISTERS[18][25] ), .ZN(n37284) );
  AOI22_X1 U451 ( .A1(n37716), .A2(\REGISTERS[5][25] ), .B1(n37718), .B2(
        \REGISTERS[28][25] ), .ZN(n37285) );
  NAND4_X1 U452 ( .A1(n37282), .A2(n37283), .A3(n37284), .A4(n37285), .ZN(
        n37286) );
  AOI22_X1 U453 ( .A1(n37709), .A2(\REGISTERS[25][25] ), .B1(n37720), .B2(
        \REGISTERS[11][25] ), .ZN(n37287) );
  AOI22_X1 U454 ( .A1(n37725), .A2(\REGISTERS[31][25] ), .B1(n37721), .B2(
        \REGISTERS[2][25] ), .ZN(n37288) );
  AOI222_X1 U455 ( .A1(n37696), .A2(\REGISTERS[29][25] ), .B1(n37697), .B2(
        \REGISTERS[13][25] ), .C1(n37722), .C2(\REGISTERS[19][25] ), .ZN(
        n37289) );
  NAND3_X1 U456 ( .A1(n37287), .A2(n37288), .A3(n37289), .ZN(n37290) );
  AOI22_X1 U457 ( .A1(n37712), .A2(\REGISTERS[26][25] ), .B1(n37715), .B2(
        \REGISTERS[8][25] ), .ZN(n37291) );
  AOI22_X1 U458 ( .A1(n37714), .A2(\REGISTERS[30][25] ), .B1(n37711), .B2(
        \REGISTERS[3][25] ), .ZN(n37292) );
  AOI22_X1 U459 ( .A1(n37719), .A2(\REGISTERS[17][25] ), .B1(n37717), .B2(
        \REGISTERS[4][25] ), .ZN(n37293) );
  AOI22_X1 U460 ( .A1(n37713), .A2(\REGISTERS[22][25] ), .B1(n37724), .B2(
        \REGISTERS[15][25] ), .ZN(n37294) );
  NAND4_X1 U461 ( .A1(n37291), .A2(n37292), .A3(n37293), .A4(n37294), .ZN(
        n37295) );
  OR4_X1 U462 ( .A1(n37281), .A2(n37286), .A3(n37290), .A4(n37295), .ZN(
        OUTB[25]) );
  AOI22_X1 U463 ( .A1(n37702), .A2(\REGISTERS[9][24] ), .B1(n37701), .B2(
        \REGISTERS[16][24] ), .ZN(n37296) );
  AOI22_X1 U464 ( .A1(n37708), .A2(\REGISTERS[23][24] ), .B1(n37710), .B2(
        \REGISTERS[6][24] ), .ZN(n37297) );
  AOI22_X1 U465 ( .A1(n37706), .A2(\REGISTERS[14][24] ), .B1(n37707), .B2(
        \REGISTERS[24][24] ), .ZN(n37298) );
  AOI22_X1 U466 ( .A1(n37704), .A2(\REGISTERS[10][24] ), .B1(n37705), .B2(
        \REGISTERS[12][24] ), .ZN(n37299) );
  NAND4_X1 U467 ( .A1(n37296), .A2(n37297), .A3(n37298), .A4(n37299), .ZN(
        n37300) );
  AOI22_X1 U468 ( .A1(n37723), .A2(\REGISTERS[27][24] ), .B1(n37703), .B2(
        \REGISTERS[1][24] ), .ZN(n37301) );
  AOI22_X1 U469 ( .A1(n37695), .A2(\REGISTERS[21][24] ), .B1(n37699), .B2(
        \REGISTERS[20][24] ), .ZN(n37302) );
  AOI22_X1 U470 ( .A1(n37698), .A2(\REGISTERS[7][24] ), .B1(n37700), .B2(
        \REGISTERS[18][24] ), .ZN(n37303) );
  AOI22_X1 U471 ( .A1(n37716), .A2(\REGISTERS[5][24] ), .B1(n37718), .B2(
        \REGISTERS[28][24] ), .ZN(n37304) );
  NAND4_X1 U472 ( .A1(n37301), .A2(n37302), .A3(n37303), .A4(n37304), .ZN(
        n37305) );
  AOI22_X1 U473 ( .A1(n37709), .A2(\REGISTERS[25][24] ), .B1(n37720), .B2(
        \REGISTERS[11][24] ), .ZN(n37306) );
  AOI22_X1 U474 ( .A1(n37725), .A2(\REGISTERS[31][24] ), .B1(n37721), .B2(
        \REGISTERS[2][24] ), .ZN(n37307) );
  AOI222_X1 U475 ( .A1(n37696), .A2(\REGISTERS[29][24] ), .B1(n37697), .B2(
        \REGISTERS[13][24] ), .C1(n37722), .C2(\REGISTERS[19][24] ), .ZN(
        n37308) );
  NAND3_X1 U476 ( .A1(n37306), .A2(n37307), .A3(n37308), .ZN(n37309) );
  AOI22_X1 U477 ( .A1(n37712), .A2(\REGISTERS[26][24] ), .B1(n37715), .B2(
        \REGISTERS[8][24] ), .ZN(n37310) );
  AOI22_X1 U478 ( .A1(n37714), .A2(\REGISTERS[30][24] ), .B1(n37711), .B2(
        \REGISTERS[3][24] ), .ZN(n37311) );
  AOI22_X1 U479 ( .A1(n37719), .A2(\REGISTERS[17][24] ), .B1(n37717), .B2(
        \REGISTERS[4][24] ), .ZN(n37312) );
  AOI22_X1 U480 ( .A1(n37713), .A2(\REGISTERS[22][24] ), .B1(n37724), .B2(
        \REGISTERS[15][24] ), .ZN(n37313) );
  NAND4_X1 U481 ( .A1(n37310), .A2(n37311), .A3(n37312), .A4(n37313), .ZN(
        n37314) );
  OR4_X1 U482 ( .A1(n37300), .A2(n37305), .A3(n37309), .A4(n37314), .ZN(
        OUTB[24]) );
  AOI22_X1 U483 ( .A1(n37702), .A2(\REGISTERS[9][23] ), .B1(n37701), .B2(
        \REGISTERS[16][23] ), .ZN(n37315) );
  AOI22_X1 U484 ( .A1(n37708), .A2(\REGISTERS[23][23] ), .B1(n37710), .B2(
        \REGISTERS[6][23] ), .ZN(n37316) );
  AOI22_X1 U485 ( .A1(n37706), .A2(\REGISTERS[14][23] ), .B1(n37707), .B2(
        \REGISTERS[24][23] ), .ZN(n37317) );
  AOI22_X1 U486 ( .A1(n37704), .A2(\REGISTERS[10][23] ), .B1(n37705), .B2(
        \REGISTERS[12][23] ), .ZN(n37318) );
  NAND4_X1 U487 ( .A1(n37315), .A2(n37316), .A3(n37317), .A4(n37318), .ZN(
        n37319) );
  AOI22_X1 U488 ( .A1(n37723), .A2(\REGISTERS[27][23] ), .B1(n37703), .B2(
        \REGISTERS[1][23] ), .ZN(n37320) );
  AOI22_X1 U489 ( .A1(n37695), .A2(\REGISTERS[21][23] ), .B1(n37699), .B2(
        \REGISTERS[20][23] ), .ZN(n37321) );
  AOI22_X1 U490 ( .A1(n37698), .A2(\REGISTERS[7][23] ), .B1(n37700), .B2(
        \REGISTERS[18][23] ), .ZN(n37322) );
  AOI22_X1 U491 ( .A1(n37716), .A2(\REGISTERS[5][23] ), .B1(n37718), .B2(
        \REGISTERS[28][23] ), .ZN(n37323) );
  NAND4_X1 U492 ( .A1(n37320), .A2(n37321), .A3(n37322), .A4(n37323), .ZN(
        n37324) );
  AOI22_X1 U493 ( .A1(n37709), .A2(\REGISTERS[25][23] ), .B1(n37720), .B2(
        \REGISTERS[11][23] ), .ZN(n37325) );
  AOI22_X1 U494 ( .A1(n37725), .A2(\REGISTERS[31][23] ), .B1(n37721), .B2(
        \REGISTERS[2][23] ), .ZN(n37326) );
  AOI222_X1 U495 ( .A1(n37696), .A2(\REGISTERS[29][23] ), .B1(n37697), .B2(
        \REGISTERS[13][23] ), .C1(n37722), .C2(\REGISTERS[19][23] ), .ZN(
        n37327) );
  NAND3_X1 U496 ( .A1(n37325), .A2(n37326), .A3(n37327), .ZN(n37328) );
  AOI22_X1 U497 ( .A1(n37712), .A2(\REGISTERS[26][23] ), .B1(n37715), .B2(
        \REGISTERS[8][23] ), .ZN(n37329) );
  AOI22_X1 U498 ( .A1(n37714), .A2(\REGISTERS[30][23] ), .B1(n37711), .B2(
        \REGISTERS[3][23] ), .ZN(n37330) );
  AOI22_X1 U499 ( .A1(n37719), .A2(\REGISTERS[17][23] ), .B1(n37717), .B2(
        \REGISTERS[4][23] ), .ZN(n37331) );
  AOI22_X1 U500 ( .A1(n37713), .A2(\REGISTERS[22][23] ), .B1(n37724), .B2(
        \REGISTERS[15][23] ), .ZN(n37332) );
  NAND4_X1 U501 ( .A1(n37329), .A2(n37330), .A3(n37331), .A4(n37332), .ZN(
        n37333) );
  OR4_X1 U502 ( .A1(n37319), .A2(n37324), .A3(n37328), .A4(n37333), .ZN(
        OUTB[23]) );
  AOI22_X1 U503 ( .A1(n37702), .A2(\REGISTERS[9][22] ), .B1(n37701), .B2(
        \REGISTERS[16][22] ), .ZN(n37334) );
  AOI22_X1 U504 ( .A1(n37708), .A2(\REGISTERS[23][22] ), .B1(n37710), .B2(
        \REGISTERS[6][22] ), .ZN(n37335) );
  AOI22_X1 U505 ( .A1(n37706), .A2(\REGISTERS[14][22] ), .B1(n37707), .B2(
        \REGISTERS[24][22] ), .ZN(n37336) );
  AOI22_X1 U506 ( .A1(n37704), .A2(\REGISTERS[10][22] ), .B1(n37705), .B2(
        \REGISTERS[12][22] ), .ZN(n37337) );
  NAND4_X1 U507 ( .A1(n37334), .A2(n37335), .A3(n37336), .A4(n37337), .ZN(
        n37338) );
  AOI22_X1 U508 ( .A1(n37723), .A2(\REGISTERS[27][22] ), .B1(n37703), .B2(
        \REGISTERS[1][22] ), .ZN(n37339) );
  AOI22_X1 U509 ( .A1(n37695), .A2(\REGISTERS[21][22] ), .B1(n37699), .B2(
        \REGISTERS[20][22] ), .ZN(n37340) );
  AOI22_X1 U510 ( .A1(n37698), .A2(\REGISTERS[7][22] ), .B1(n37700), .B2(
        \REGISTERS[18][22] ), .ZN(n37341) );
  AOI22_X1 U511 ( .A1(n37716), .A2(\REGISTERS[5][22] ), .B1(n37718), .B2(
        \REGISTERS[28][22] ), .ZN(n37342) );
  NAND4_X1 U512 ( .A1(n37339), .A2(n37340), .A3(n37341), .A4(n37342), .ZN(
        n37343) );
  AOI22_X1 U513 ( .A1(n37709), .A2(\REGISTERS[25][22] ), .B1(n37720), .B2(
        \REGISTERS[11][22] ), .ZN(n37344) );
  AOI22_X1 U514 ( .A1(n37725), .A2(\REGISTERS[31][22] ), .B1(n37721), .B2(
        \REGISTERS[2][22] ), .ZN(n37345) );
  AOI222_X1 U515 ( .A1(n37696), .A2(\REGISTERS[29][22] ), .B1(n37697), .B2(
        \REGISTERS[13][22] ), .C1(n37722), .C2(\REGISTERS[19][22] ), .ZN(
        n37346) );
  NAND3_X1 U516 ( .A1(n37344), .A2(n37345), .A3(n37346), .ZN(n37347) );
  AOI22_X1 U517 ( .A1(n37712), .A2(\REGISTERS[26][22] ), .B1(n37715), .B2(
        \REGISTERS[8][22] ), .ZN(n37348) );
  AOI22_X1 U518 ( .A1(n37714), .A2(\REGISTERS[30][22] ), .B1(n37711), .B2(
        \REGISTERS[3][22] ), .ZN(n37349) );
  AOI22_X1 U519 ( .A1(n37719), .A2(\REGISTERS[17][22] ), .B1(n37717), .B2(
        \REGISTERS[4][22] ), .ZN(n37350) );
  AOI22_X1 U520 ( .A1(n37713), .A2(\REGISTERS[22][22] ), .B1(n37724), .B2(
        \REGISTERS[15][22] ), .ZN(n37351) );
  NAND4_X1 U521 ( .A1(n37348), .A2(n37349), .A3(n37350), .A4(n37351), .ZN(
        n37352) );
  OR4_X1 U522 ( .A1(n37338), .A2(n37343), .A3(n37347), .A4(n37352), .ZN(
        OUTB[22]) );
  AOI22_X1 U523 ( .A1(n37702), .A2(\REGISTERS[9][21] ), .B1(n37701), .B2(
        \REGISTERS[16][21] ), .ZN(n37353) );
  AOI22_X1 U524 ( .A1(n37708), .A2(\REGISTERS[23][21] ), .B1(n37710), .B2(
        \REGISTERS[6][21] ), .ZN(n37354) );
  AOI22_X1 U525 ( .A1(n37706), .A2(\REGISTERS[14][21] ), .B1(n37707), .B2(
        \REGISTERS[24][21] ), .ZN(n37355) );
  AOI22_X1 U526 ( .A1(n37704), .A2(\REGISTERS[10][21] ), .B1(n37705), .B2(
        \REGISTERS[12][21] ), .ZN(n37356) );
  NAND4_X1 U527 ( .A1(n37353), .A2(n37354), .A3(n37355), .A4(n37356), .ZN(
        n37357) );
  AOI22_X1 U528 ( .A1(n37723), .A2(\REGISTERS[27][21] ), .B1(n37703), .B2(
        \REGISTERS[1][21] ), .ZN(n37358) );
  AOI22_X1 U529 ( .A1(n37695), .A2(\REGISTERS[21][21] ), .B1(n37699), .B2(
        \REGISTERS[20][21] ), .ZN(n37359) );
  AOI22_X1 U530 ( .A1(n37698), .A2(\REGISTERS[7][21] ), .B1(n37700), .B2(
        \REGISTERS[18][21] ), .ZN(n37360) );
  AOI22_X1 U531 ( .A1(n37716), .A2(\REGISTERS[5][21] ), .B1(n37718), .B2(
        \REGISTERS[28][21] ), .ZN(n37361) );
  NAND4_X1 U532 ( .A1(n37358), .A2(n37359), .A3(n37360), .A4(n37361), .ZN(
        n37362) );
  AOI22_X1 U533 ( .A1(n37709), .A2(\REGISTERS[25][21] ), .B1(n37720), .B2(
        \REGISTERS[11][21] ), .ZN(n37363) );
  AOI22_X1 U534 ( .A1(n37725), .A2(\REGISTERS[31][21] ), .B1(n37721), .B2(
        \REGISTERS[2][21] ), .ZN(n37364) );
  AOI222_X1 U535 ( .A1(n37696), .A2(\REGISTERS[29][21] ), .B1(n37697), .B2(
        \REGISTERS[13][21] ), .C1(n37722), .C2(\REGISTERS[19][21] ), .ZN(
        n37365) );
  NAND3_X1 U536 ( .A1(n37363), .A2(n37364), .A3(n37365), .ZN(n37366) );
  AOI22_X1 U537 ( .A1(n37712), .A2(\REGISTERS[26][21] ), .B1(n37715), .B2(
        \REGISTERS[8][21] ), .ZN(n37367) );
  AOI22_X1 U538 ( .A1(n37714), .A2(\REGISTERS[30][21] ), .B1(n37711), .B2(
        \REGISTERS[3][21] ), .ZN(n37368) );
  AOI22_X1 U539 ( .A1(n37719), .A2(\REGISTERS[17][21] ), .B1(n37717), .B2(
        \REGISTERS[4][21] ), .ZN(n37369) );
  AOI22_X1 U540 ( .A1(n37713), .A2(\REGISTERS[22][21] ), .B1(n37724), .B2(
        \REGISTERS[15][21] ), .ZN(n37370) );
  NAND4_X1 U541 ( .A1(n37367), .A2(n37368), .A3(n37369), .A4(n37370), .ZN(
        n37371) );
  OR4_X1 U542 ( .A1(n37357), .A2(n37362), .A3(n37366), .A4(n37371), .ZN(
        OUTB[21]) );
  AOI22_X1 U543 ( .A1(n37702), .A2(\REGISTERS[9][20] ), .B1(n37701), .B2(
        \REGISTERS[16][20] ), .ZN(n37372) );
  AOI22_X1 U544 ( .A1(n37708), .A2(\REGISTERS[23][20] ), .B1(n37710), .B2(
        \REGISTERS[6][20] ), .ZN(n37373) );
  AOI22_X1 U545 ( .A1(n37706), .A2(\REGISTERS[14][20] ), .B1(n37707), .B2(
        \REGISTERS[24][20] ), .ZN(n37374) );
  AOI22_X1 U546 ( .A1(n37704), .A2(\REGISTERS[10][20] ), .B1(n37705), .B2(
        \REGISTERS[12][20] ), .ZN(n37375) );
  NAND4_X1 U547 ( .A1(n37372), .A2(n37373), .A3(n37374), .A4(n37375), .ZN(
        n37376) );
  AOI22_X1 U548 ( .A1(n37723), .A2(\REGISTERS[27][20] ), .B1(n37703), .B2(
        \REGISTERS[1][20] ), .ZN(n37377) );
  AOI22_X1 U549 ( .A1(n37695), .A2(\REGISTERS[21][20] ), .B1(n37699), .B2(
        \REGISTERS[20][20] ), .ZN(n37378) );
  AOI22_X1 U550 ( .A1(n37698), .A2(\REGISTERS[7][20] ), .B1(n37700), .B2(
        \REGISTERS[18][20] ), .ZN(n37379) );
  AOI22_X1 U551 ( .A1(n37716), .A2(\REGISTERS[5][20] ), .B1(n37718), .B2(
        \REGISTERS[28][20] ), .ZN(n37380) );
  NAND4_X1 U552 ( .A1(n37377), .A2(n37378), .A3(n37379), .A4(n37380), .ZN(
        n37381) );
  AOI22_X1 U553 ( .A1(n37709), .A2(\REGISTERS[25][20] ), .B1(n37720), .B2(
        \REGISTERS[11][20] ), .ZN(n37382) );
  AOI22_X1 U554 ( .A1(n37725), .A2(\REGISTERS[31][20] ), .B1(n37721), .B2(
        \REGISTERS[2][20] ), .ZN(n37383) );
  AOI222_X1 U555 ( .A1(n37696), .A2(\REGISTERS[29][20] ), .B1(n37697), .B2(
        \REGISTERS[13][20] ), .C1(n37722), .C2(\REGISTERS[19][20] ), .ZN(
        n37384) );
  NAND3_X1 U556 ( .A1(n37382), .A2(n37383), .A3(n37384), .ZN(n37385) );
  AOI22_X1 U557 ( .A1(n37712), .A2(\REGISTERS[26][20] ), .B1(n37715), .B2(
        \REGISTERS[8][20] ), .ZN(n37386) );
  AOI22_X1 U558 ( .A1(n37714), .A2(\REGISTERS[30][20] ), .B1(n37711), .B2(
        \REGISTERS[3][20] ), .ZN(n37387) );
  AOI22_X1 U559 ( .A1(n37719), .A2(\REGISTERS[17][20] ), .B1(n37717), .B2(
        \REGISTERS[4][20] ), .ZN(n37388) );
  AOI22_X1 U560 ( .A1(n37713), .A2(\REGISTERS[22][20] ), .B1(n37724), .B2(
        \REGISTERS[15][20] ), .ZN(n37389) );
  NAND4_X1 U561 ( .A1(n37386), .A2(n37387), .A3(n37388), .A4(n37389), .ZN(
        n37390) );
  OR4_X1 U562 ( .A1(n37376), .A2(n37381), .A3(n37385), .A4(n37390), .ZN(
        OUTB[20]) );
  AOI22_X1 U563 ( .A1(n37702), .A2(\REGISTERS[9][19] ), .B1(n37701), .B2(
        \REGISTERS[16][19] ), .ZN(n37391) );
  AOI22_X1 U564 ( .A1(n37708), .A2(\REGISTERS[23][19] ), .B1(n37710), .B2(
        \REGISTERS[6][19] ), .ZN(n37392) );
  AOI22_X1 U565 ( .A1(n37706), .A2(\REGISTERS[14][19] ), .B1(n37707), .B2(
        \REGISTERS[24][19] ), .ZN(n37393) );
  AOI22_X1 U566 ( .A1(n37704), .A2(\REGISTERS[10][19] ), .B1(n37705), .B2(
        \REGISTERS[12][19] ), .ZN(n37394) );
  NAND4_X1 U567 ( .A1(n37391), .A2(n37392), .A3(n37393), .A4(n37394), .ZN(
        n37395) );
  AOI22_X1 U568 ( .A1(n37723), .A2(\REGISTERS[27][19] ), .B1(n37703), .B2(
        \REGISTERS[1][19] ), .ZN(n37396) );
  AOI22_X1 U569 ( .A1(n37695), .A2(\REGISTERS[21][19] ), .B1(n37699), .B2(
        \REGISTERS[20][19] ), .ZN(n37397) );
  AOI22_X1 U570 ( .A1(n37698), .A2(\REGISTERS[7][19] ), .B1(n37700), .B2(
        \REGISTERS[18][19] ), .ZN(n37398) );
  AOI22_X1 U571 ( .A1(n37716), .A2(\REGISTERS[5][19] ), .B1(n37718), .B2(
        \REGISTERS[28][19] ), .ZN(n37399) );
  NAND4_X1 U572 ( .A1(n37396), .A2(n37397), .A3(n37398), .A4(n37399), .ZN(
        n37400) );
  AOI22_X1 U573 ( .A1(n37709), .A2(\REGISTERS[25][19] ), .B1(n37720), .B2(
        \REGISTERS[11][19] ), .ZN(n37401) );
  AOI22_X1 U574 ( .A1(n37725), .A2(\REGISTERS[31][19] ), .B1(n37721), .B2(
        \REGISTERS[2][19] ), .ZN(n37402) );
  AOI222_X1 U575 ( .A1(n37696), .A2(\REGISTERS[29][19] ), .B1(n37697), .B2(
        \REGISTERS[13][19] ), .C1(n37722), .C2(\REGISTERS[19][19] ), .ZN(
        n37403) );
  NAND3_X1 U576 ( .A1(n37401), .A2(n37402), .A3(n37403), .ZN(n37404) );
  AOI22_X1 U577 ( .A1(n37712), .A2(\REGISTERS[26][19] ), .B1(n37715), .B2(
        \REGISTERS[8][19] ), .ZN(n37405) );
  AOI22_X1 U578 ( .A1(n37714), .A2(\REGISTERS[30][19] ), .B1(n37711), .B2(
        \REGISTERS[3][19] ), .ZN(n37406) );
  AOI22_X1 U579 ( .A1(n37719), .A2(\REGISTERS[17][19] ), .B1(n37717), .B2(
        \REGISTERS[4][19] ), .ZN(n37407) );
  AOI22_X1 U580 ( .A1(n37713), .A2(\REGISTERS[22][19] ), .B1(n37724), .B2(
        \REGISTERS[15][19] ), .ZN(n37408) );
  NAND4_X1 U581 ( .A1(n37405), .A2(n37406), .A3(n37407), .A4(n37408), .ZN(
        n37409) );
  OR4_X1 U582 ( .A1(n37395), .A2(n37400), .A3(n37404), .A4(n37409), .ZN(
        OUTB[19]) );
  AOI22_X1 U583 ( .A1(n37702), .A2(\REGISTERS[9][18] ), .B1(n37701), .B2(
        \REGISTERS[16][18] ), .ZN(n37410) );
  AOI22_X1 U584 ( .A1(n37708), .A2(\REGISTERS[23][18] ), .B1(n37710), .B2(
        \REGISTERS[6][18] ), .ZN(n37411) );
  AOI22_X1 U585 ( .A1(n37706), .A2(\REGISTERS[14][18] ), .B1(n37707), .B2(
        \REGISTERS[24][18] ), .ZN(n37412) );
  AOI22_X1 U586 ( .A1(n37704), .A2(\REGISTERS[10][18] ), .B1(n37705), .B2(
        \REGISTERS[12][18] ), .ZN(n37413) );
  NAND4_X1 U587 ( .A1(n37410), .A2(n37411), .A3(n37412), .A4(n37413), .ZN(
        n37414) );
  AOI22_X1 U588 ( .A1(n37723), .A2(\REGISTERS[27][18] ), .B1(n37703), .B2(
        \REGISTERS[1][18] ), .ZN(n37415) );
  AOI22_X1 U589 ( .A1(n37695), .A2(\REGISTERS[21][18] ), .B1(n37699), .B2(
        \REGISTERS[20][18] ), .ZN(n37416) );
  AOI22_X1 U590 ( .A1(n37698), .A2(\REGISTERS[7][18] ), .B1(n37700), .B2(
        \REGISTERS[18][18] ), .ZN(n37417) );
  AOI22_X1 U591 ( .A1(n37716), .A2(\REGISTERS[5][18] ), .B1(n37718), .B2(
        \REGISTERS[28][18] ), .ZN(n37418) );
  NAND4_X1 U592 ( .A1(n37415), .A2(n37416), .A3(n37417), .A4(n37418), .ZN(
        n37419) );
  AOI22_X1 U593 ( .A1(n37709), .A2(\REGISTERS[25][18] ), .B1(n37720), .B2(
        \REGISTERS[11][18] ), .ZN(n37420) );
  AOI22_X1 U594 ( .A1(n37725), .A2(\REGISTERS[31][18] ), .B1(n37721), .B2(
        \REGISTERS[2][18] ), .ZN(n37421) );
  AOI222_X1 U595 ( .A1(n37696), .A2(\REGISTERS[29][18] ), .B1(n37697), .B2(
        \REGISTERS[13][18] ), .C1(n37722), .C2(\REGISTERS[19][18] ), .ZN(
        n37422) );
  NAND3_X1 U596 ( .A1(n37420), .A2(n37421), .A3(n37422), .ZN(n37423) );
  AOI22_X1 U597 ( .A1(n37712), .A2(\REGISTERS[26][18] ), .B1(n37715), .B2(
        \REGISTERS[8][18] ), .ZN(n37424) );
  AOI22_X1 U598 ( .A1(n37714), .A2(\REGISTERS[30][18] ), .B1(n37711), .B2(
        \REGISTERS[3][18] ), .ZN(n37425) );
  AOI22_X1 U599 ( .A1(n37719), .A2(\REGISTERS[17][18] ), .B1(n37717), .B2(
        \REGISTERS[4][18] ), .ZN(n37426) );
  AOI22_X1 U600 ( .A1(n37713), .A2(\REGISTERS[22][18] ), .B1(n37724), .B2(
        \REGISTERS[15][18] ), .ZN(n37427) );
  NAND4_X1 U601 ( .A1(n37424), .A2(n37425), .A3(n37426), .A4(n37427), .ZN(
        n37428) );
  OR4_X1 U602 ( .A1(n37414), .A2(n37419), .A3(n37423), .A4(n37428), .ZN(
        OUTB[18]) );
  AOI22_X1 U603 ( .A1(n37702), .A2(\REGISTERS[9][17] ), .B1(n37701), .B2(
        \REGISTERS[16][17] ), .ZN(n37429) );
  AOI22_X1 U604 ( .A1(n37708), .A2(\REGISTERS[23][17] ), .B1(n37710), .B2(
        \REGISTERS[6][17] ), .ZN(n37430) );
  AOI22_X1 U605 ( .A1(n37706), .A2(\REGISTERS[14][17] ), .B1(n37707), .B2(
        \REGISTERS[24][17] ), .ZN(n37431) );
  AOI22_X1 U606 ( .A1(n37704), .A2(\REGISTERS[10][17] ), .B1(n37705), .B2(
        \REGISTERS[12][17] ), .ZN(n37432) );
  NAND4_X1 U607 ( .A1(n37429), .A2(n37430), .A3(n37431), .A4(n37432), .ZN(
        n37433) );
  AOI22_X1 U608 ( .A1(n37723), .A2(\REGISTERS[27][17] ), .B1(n37703), .B2(
        \REGISTERS[1][17] ), .ZN(n37434) );
  AOI22_X1 U609 ( .A1(n37695), .A2(\REGISTERS[21][17] ), .B1(n37699), .B2(
        \REGISTERS[20][17] ), .ZN(n37435) );
  AOI22_X1 U610 ( .A1(n37698), .A2(\REGISTERS[7][17] ), .B1(n37700), .B2(
        \REGISTERS[18][17] ), .ZN(n37436) );
  AOI22_X1 U611 ( .A1(n37716), .A2(\REGISTERS[5][17] ), .B1(n37718), .B2(
        \REGISTERS[28][17] ), .ZN(n37437) );
  NAND4_X1 U612 ( .A1(n37434), .A2(n37435), .A3(n37436), .A4(n37437), .ZN(
        n37438) );
  AOI22_X1 U613 ( .A1(n37709), .A2(\REGISTERS[25][17] ), .B1(n37720), .B2(
        \REGISTERS[11][17] ), .ZN(n37439) );
  AOI22_X1 U614 ( .A1(n37725), .A2(\REGISTERS[31][17] ), .B1(n37721), .B2(
        \REGISTERS[2][17] ), .ZN(n37440) );
  AOI222_X1 U615 ( .A1(n37696), .A2(\REGISTERS[29][17] ), .B1(n37697), .B2(
        \REGISTERS[13][17] ), .C1(n37722), .C2(\REGISTERS[19][17] ), .ZN(
        n37441) );
  NAND3_X1 U616 ( .A1(n37439), .A2(n37440), .A3(n37441), .ZN(n37442) );
  AOI22_X1 U617 ( .A1(n37712), .A2(\REGISTERS[26][17] ), .B1(n37715), .B2(
        \REGISTERS[8][17] ), .ZN(n37443) );
  AOI22_X1 U618 ( .A1(n37714), .A2(\REGISTERS[30][17] ), .B1(n37711), .B2(
        \REGISTERS[3][17] ), .ZN(n37444) );
  AOI22_X1 U619 ( .A1(n37719), .A2(\REGISTERS[17][17] ), .B1(n37717), .B2(
        \REGISTERS[4][17] ), .ZN(n37445) );
  AOI22_X1 U620 ( .A1(n37713), .A2(\REGISTERS[22][17] ), .B1(n37724), .B2(
        \REGISTERS[15][17] ), .ZN(n37446) );
  NAND4_X1 U621 ( .A1(n37443), .A2(n37444), .A3(n37445), .A4(n37446), .ZN(
        n37447) );
  OR4_X1 U622 ( .A1(n37433), .A2(n37438), .A3(n37442), .A4(n37447), .ZN(
        OUTB[17]) );
  AOI22_X1 U623 ( .A1(n37702), .A2(\REGISTERS[9][16] ), .B1(n37701), .B2(
        \REGISTERS[16][16] ), .ZN(n37448) );
  AOI22_X1 U624 ( .A1(n37708), .A2(\REGISTERS[23][16] ), .B1(n37710), .B2(
        \REGISTERS[6][16] ), .ZN(n37449) );
  AOI22_X1 U625 ( .A1(n37706), .A2(\REGISTERS[14][16] ), .B1(n37707), .B2(
        \REGISTERS[24][16] ), .ZN(n37450) );
  AOI22_X1 U626 ( .A1(n37704), .A2(\REGISTERS[10][16] ), .B1(n37705), .B2(
        \REGISTERS[12][16] ), .ZN(n37451) );
  NAND4_X1 U627 ( .A1(n37448), .A2(n37449), .A3(n37450), .A4(n37451), .ZN(
        n37452) );
  AOI22_X1 U628 ( .A1(n37723), .A2(\REGISTERS[27][16] ), .B1(n37703), .B2(
        \REGISTERS[1][16] ), .ZN(n37453) );
  AOI22_X1 U629 ( .A1(n37695), .A2(\REGISTERS[21][16] ), .B1(n37699), .B2(
        \REGISTERS[20][16] ), .ZN(n37454) );
  AOI22_X1 U630 ( .A1(n37698), .A2(\REGISTERS[7][16] ), .B1(n37700), .B2(
        \REGISTERS[18][16] ), .ZN(n37455) );
  AOI22_X1 U631 ( .A1(n37716), .A2(\REGISTERS[5][16] ), .B1(n37718), .B2(
        \REGISTERS[28][16] ), .ZN(n37456) );
  NAND4_X1 U632 ( .A1(n37453), .A2(n37454), .A3(n37455), .A4(n37456), .ZN(
        n37457) );
  AOI22_X1 U633 ( .A1(n37709), .A2(\REGISTERS[25][16] ), .B1(n37720), .B2(
        \REGISTERS[11][16] ), .ZN(n37458) );
  AOI22_X1 U634 ( .A1(n37725), .A2(\REGISTERS[31][16] ), .B1(n37721), .B2(
        \REGISTERS[2][16] ), .ZN(n37459) );
  AOI222_X1 U635 ( .A1(n37696), .A2(\REGISTERS[29][16] ), .B1(n37697), .B2(
        \REGISTERS[13][16] ), .C1(n37722), .C2(\REGISTERS[19][16] ), .ZN(
        n37460) );
  NAND3_X1 U636 ( .A1(n37458), .A2(n37459), .A3(n37460), .ZN(n37461) );
  AOI22_X1 U637 ( .A1(n37712), .A2(\REGISTERS[26][16] ), .B1(n37715), .B2(
        \REGISTERS[8][16] ), .ZN(n37462) );
  AOI22_X1 U638 ( .A1(n37714), .A2(\REGISTERS[30][16] ), .B1(n37711), .B2(
        \REGISTERS[3][16] ), .ZN(n37463) );
  AOI22_X1 U639 ( .A1(n37719), .A2(\REGISTERS[17][16] ), .B1(n37717), .B2(
        \REGISTERS[4][16] ), .ZN(n37464) );
  AOI22_X1 U640 ( .A1(n37713), .A2(\REGISTERS[22][16] ), .B1(n37724), .B2(
        \REGISTERS[15][16] ), .ZN(n37465) );
  NAND4_X1 U641 ( .A1(n37462), .A2(n37463), .A3(n37464), .A4(n37465), .ZN(
        n37466) );
  OR4_X1 U642 ( .A1(n37452), .A2(n37457), .A3(n37461), .A4(n37466), .ZN(
        OUTB[16]) );
  AOI22_X1 U643 ( .A1(n37702), .A2(\REGISTERS[9][15] ), .B1(n37701), .B2(
        \REGISTERS[16][15] ), .ZN(n37467) );
  AOI22_X1 U644 ( .A1(n37708), .A2(\REGISTERS[23][15] ), .B1(n37710), .B2(
        \REGISTERS[6][15] ), .ZN(n37468) );
  AOI22_X1 U645 ( .A1(n37706), .A2(\REGISTERS[14][15] ), .B1(n37707), .B2(
        \REGISTERS[24][15] ), .ZN(n37469) );
  AOI22_X1 U646 ( .A1(n37704), .A2(\REGISTERS[10][15] ), .B1(n37705), .B2(
        \REGISTERS[12][15] ), .ZN(n37470) );
  NAND4_X1 U647 ( .A1(n37467), .A2(n37468), .A3(n37469), .A4(n37470), .ZN(
        n37471) );
  AOI22_X1 U648 ( .A1(n37723), .A2(\REGISTERS[27][15] ), .B1(n37703), .B2(
        \REGISTERS[1][15] ), .ZN(n37472) );
  AOI22_X1 U649 ( .A1(n37695), .A2(\REGISTERS[21][15] ), .B1(n37699), .B2(
        \REGISTERS[20][15] ), .ZN(n37473) );
  AOI22_X1 U650 ( .A1(n37698), .A2(\REGISTERS[7][15] ), .B1(n37700), .B2(
        \REGISTERS[18][15] ), .ZN(n37474) );
  AOI22_X1 U651 ( .A1(n37716), .A2(\REGISTERS[5][15] ), .B1(n37718), .B2(
        \REGISTERS[28][15] ), .ZN(n37475) );
  NAND4_X1 U652 ( .A1(n37472), .A2(n37473), .A3(n37474), .A4(n37475), .ZN(
        n37476) );
  AOI22_X1 U653 ( .A1(n37709), .A2(\REGISTERS[25][15] ), .B1(n37720), .B2(
        \REGISTERS[11][15] ), .ZN(n37477) );
  AOI22_X1 U654 ( .A1(n37725), .A2(\REGISTERS[31][15] ), .B1(n37721), .B2(
        \REGISTERS[2][15] ), .ZN(n37478) );
  AOI222_X1 U655 ( .A1(n37696), .A2(\REGISTERS[29][15] ), .B1(n37697), .B2(
        \REGISTERS[13][15] ), .C1(n37722), .C2(\REGISTERS[19][15] ), .ZN(
        n37479) );
  NAND3_X1 U656 ( .A1(n37477), .A2(n37478), .A3(n37479), .ZN(n37480) );
  AOI22_X1 U657 ( .A1(n37712), .A2(\REGISTERS[26][15] ), .B1(n37715), .B2(
        \REGISTERS[8][15] ), .ZN(n37481) );
  AOI22_X1 U658 ( .A1(n37714), .A2(\REGISTERS[30][15] ), .B1(n37711), .B2(
        \REGISTERS[3][15] ), .ZN(n37482) );
  AOI22_X1 U659 ( .A1(n37719), .A2(\REGISTERS[17][15] ), .B1(n37717), .B2(
        \REGISTERS[4][15] ), .ZN(n37483) );
  AOI22_X1 U660 ( .A1(n37713), .A2(\REGISTERS[22][15] ), .B1(n37724), .B2(
        \REGISTERS[15][15] ), .ZN(n37484) );
  NAND4_X1 U661 ( .A1(n37481), .A2(n37482), .A3(n37483), .A4(n37484), .ZN(
        n37485) );
  OR4_X1 U662 ( .A1(n37471), .A2(n37476), .A3(n37480), .A4(n37485), .ZN(
        OUTB[15]) );
  AOI22_X1 U663 ( .A1(n37702), .A2(\REGISTERS[9][14] ), .B1(n37701), .B2(
        \REGISTERS[16][14] ), .ZN(n37486) );
  AOI22_X1 U664 ( .A1(n37708), .A2(\REGISTERS[23][14] ), .B1(n37710), .B2(
        \REGISTERS[6][14] ), .ZN(n37487) );
  AOI22_X1 U665 ( .A1(n37706), .A2(\REGISTERS[14][14] ), .B1(n37707), .B2(
        \REGISTERS[24][14] ), .ZN(n37488) );
  AOI22_X1 U666 ( .A1(n37704), .A2(\REGISTERS[10][14] ), .B1(n37705), .B2(
        \REGISTERS[12][14] ), .ZN(n37489) );
  NAND4_X1 U667 ( .A1(n37486), .A2(n37487), .A3(n37488), .A4(n37489), .ZN(
        n37490) );
  AOI22_X1 U668 ( .A1(n37723), .A2(\REGISTERS[27][14] ), .B1(n37703), .B2(
        \REGISTERS[1][14] ), .ZN(n37491) );
  AOI22_X1 U669 ( .A1(n37695), .A2(\REGISTERS[21][14] ), .B1(n37699), .B2(
        \REGISTERS[20][14] ), .ZN(n37492) );
  AOI22_X1 U670 ( .A1(n37698), .A2(\REGISTERS[7][14] ), .B1(n37700), .B2(
        \REGISTERS[18][14] ), .ZN(n37493) );
  AOI22_X1 U671 ( .A1(n37716), .A2(\REGISTERS[5][14] ), .B1(n37718), .B2(
        \REGISTERS[28][14] ), .ZN(n37494) );
  NAND4_X1 U672 ( .A1(n37491), .A2(n37492), .A3(n37493), .A4(n37494), .ZN(
        n37495) );
  AOI22_X1 U673 ( .A1(n37709), .A2(\REGISTERS[25][14] ), .B1(n37720), .B2(
        \REGISTERS[11][14] ), .ZN(n37496) );
  AOI22_X1 U674 ( .A1(n37725), .A2(\REGISTERS[31][14] ), .B1(n37721), .B2(
        \REGISTERS[2][14] ), .ZN(n37497) );
  AOI222_X1 U675 ( .A1(n37696), .A2(\REGISTERS[29][14] ), .B1(n37697), .B2(
        \REGISTERS[13][14] ), .C1(n37722), .C2(\REGISTERS[19][14] ), .ZN(
        n37498) );
  NAND3_X1 U676 ( .A1(n37496), .A2(n37497), .A3(n37498), .ZN(n37499) );
  AOI22_X1 U677 ( .A1(n37712), .A2(\REGISTERS[26][14] ), .B1(n37715), .B2(
        \REGISTERS[8][14] ), .ZN(n37500) );
  AOI22_X1 U678 ( .A1(n37714), .A2(\REGISTERS[30][14] ), .B1(n37711), .B2(
        \REGISTERS[3][14] ), .ZN(n37501) );
  AOI22_X1 U679 ( .A1(n37719), .A2(\REGISTERS[17][14] ), .B1(n37717), .B2(
        \REGISTERS[4][14] ), .ZN(n37502) );
  AOI22_X1 U680 ( .A1(n37713), .A2(\REGISTERS[22][14] ), .B1(n37724), .B2(
        \REGISTERS[15][14] ), .ZN(n37503) );
  NAND4_X1 U681 ( .A1(n37500), .A2(n37501), .A3(n37502), .A4(n37503), .ZN(
        n37504) );
  OR4_X1 U682 ( .A1(n37490), .A2(n37495), .A3(n37499), .A4(n37504), .ZN(
        OUTB[14]) );
  AOI22_X1 U683 ( .A1(n37702), .A2(\REGISTERS[9][13] ), .B1(n37701), .B2(
        \REGISTERS[16][13] ), .ZN(n37505) );
  AOI22_X1 U684 ( .A1(n37708), .A2(\REGISTERS[23][13] ), .B1(n37710), .B2(
        \REGISTERS[6][13] ), .ZN(n37506) );
  AOI22_X1 U685 ( .A1(n37706), .A2(\REGISTERS[14][13] ), .B1(n37707), .B2(
        \REGISTERS[24][13] ), .ZN(n37507) );
  AOI22_X1 U686 ( .A1(n37704), .A2(\REGISTERS[10][13] ), .B1(n37705), .B2(
        \REGISTERS[12][13] ), .ZN(n37508) );
  NAND4_X1 U687 ( .A1(n37505), .A2(n37506), .A3(n37507), .A4(n37508), .ZN(
        n37509) );
  AOI22_X1 U688 ( .A1(n37723), .A2(\REGISTERS[27][13] ), .B1(n37703), .B2(
        \REGISTERS[1][13] ), .ZN(n37510) );
  AOI22_X1 U689 ( .A1(n37695), .A2(\REGISTERS[21][13] ), .B1(n37699), .B2(
        \REGISTERS[20][13] ), .ZN(n37511) );
  AOI22_X1 U690 ( .A1(n37698), .A2(\REGISTERS[7][13] ), .B1(n37700), .B2(
        \REGISTERS[18][13] ), .ZN(n37512) );
  AOI22_X1 U691 ( .A1(n37716), .A2(\REGISTERS[5][13] ), .B1(n37718), .B2(
        \REGISTERS[28][13] ), .ZN(n37513) );
  NAND4_X1 U692 ( .A1(n37510), .A2(n37511), .A3(n37512), .A4(n37513), .ZN(
        n37514) );
  AOI22_X1 U693 ( .A1(n37709), .A2(\REGISTERS[25][13] ), .B1(n37720), .B2(
        \REGISTERS[11][13] ), .ZN(n37515) );
  AOI22_X1 U694 ( .A1(n37725), .A2(\REGISTERS[31][13] ), .B1(n37721), .B2(
        \REGISTERS[2][13] ), .ZN(n37516) );
  AOI222_X1 U695 ( .A1(n37696), .A2(\REGISTERS[29][13] ), .B1(n37697), .B2(
        \REGISTERS[13][13] ), .C1(n37722), .C2(\REGISTERS[19][13] ), .ZN(
        n37517) );
  NAND3_X1 U696 ( .A1(n37515), .A2(n37516), .A3(n37517), .ZN(n37518) );
  AOI22_X1 U697 ( .A1(n37712), .A2(\REGISTERS[26][13] ), .B1(n37715), .B2(
        \REGISTERS[8][13] ), .ZN(n37519) );
  AOI22_X1 U698 ( .A1(n37714), .A2(\REGISTERS[30][13] ), .B1(n37711), .B2(
        \REGISTERS[3][13] ), .ZN(n37520) );
  AOI22_X1 U699 ( .A1(n37719), .A2(\REGISTERS[17][13] ), .B1(n37717), .B2(
        \REGISTERS[4][13] ), .ZN(n37521) );
  AOI22_X1 U700 ( .A1(n37713), .A2(\REGISTERS[22][13] ), .B1(n37724), .B2(
        \REGISTERS[15][13] ), .ZN(n37522) );
  NAND4_X1 U701 ( .A1(n37519), .A2(n37520), .A3(n37521), .A4(n37522), .ZN(
        n37523) );
  OR4_X1 U702 ( .A1(n37509), .A2(n37514), .A3(n37518), .A4(n37523), .ZN(
        OUTB[13]) );
  AOI22_X1 U703 ( .A1(n37702), .A2(\REGISTERS[9][12] ), .B1(n37701), .B2(
        \REGISTERS[16][12] ), .ZN(n37524) );
  AOI22_X1 U704 ( .A1(n37708), .A2(\REGISTERS[23][12] ), .B1(n37710), .B2(
        \REGISTERS[6][12] ), .ZN(n37525) );
  AOI22_X1 U705 ( .A1(n37706), .A2(\REGISTERS[14][12] ), .B1(n37707), .B2(
        \REGISTERS[24][12] ), .ZN(n37526) );
  AOI22_X1 U706 ( .A1(n37704), .A2(\REGISTERS[10][12] ), .B1(n37705), .B2(
        \REGISTERS[12][12] ), .ZN(n37527) );
  NAND4_X1 U707 ( .A1(n37524), .A2(n37525), .A3(n37526), .A4(n37527), .ZN(
        n37528) );
  AOI22_X1 U708 ( .A1(n37723), .A2(\REGISTERS[27][12] ), .B1(n37703), .B2(
        \REGISTERS[1][12] ), .ZN(n37529) );
  AOI22_X1 U709 ( .A1(n37695), .A2(\REGISTERS[21][12] ), .B1(n37699), .B2(
        \REGISTERS[20][12] ), .ZN(n37530) );
  AOI22_X1 U710 ( .A1(n37698), .A2(\REGISTERS[7][12] ), .B1(n37700), .B2(
        \REGISTERS[18][12] ), .ZN(n37531) );
  AOI22_X1 U711 ( .A1(n37716), .A2(\REGISTERS[5][12] ), .B1(n37718), .B2(
        \REGISTERS[28][12] ), .ZN(n37532) );
  NAND4_X1 U712 ( .A1(n37529), .A2(n37530), .A3(n37531), .A4(n37532), .ZN(
        n37533) );
  AOI22_X1 U713 ( .A1(n37709), .A2(\REGISTERS[25][12] ), .B1(n37720), .B2(
        \REGISTERS[11][12] ), .ZN(n37534) );
  AOI22_X1 U714 ( .A1(n37725), .A2(\REGISTERS[31][12] ), .B1(n37721), .B2(
        \REGISTERS[2][12] ), .ZN(n37535) );
  AOI222_X1 U715 ( .A1(n37696), .A2(\REGISTERS[29][12] ), .B1(n37697), .B2(
        \REGISTERS[13][12] ), .C1(n37722), .C2(\REGISTERS[19][12] ), .ZN(
        n37536) );
  NAND3_X1 U716 ( .A1(n37534), .A2(n37535), .A3(n37536), .ZN(n37537) );
  AOI22_X1 U717 ( .A1(n37712), .A2(\REGISTERS[26][12] ), .B1(n37715), .B2(
        \REGISTERS[8][12] ), .ZN(n37538) );
  AOI22_X1 U718 ( .A1(n37714), .A2(\REGISTERS[30][12] ), .B1(n37711), .B2(
        \REGISTERS[3][12] ), .ZN(n37539) );
  AOI22_X1 U719 ( .A1(n37719), .A2(\REGISTERS[17][12] ), .B1(n37717), .B2(
        \REGISTERS[4][12] ), .ZN(n37540) );
  AOI22_X1 U720 ( .A1(n37713), .A2(\REGISTERS[22][12] ), .B1(n37724), .B2(
        \REGISTERS[15][12] ), .ZN(n37541) );
  NAND4_X1 U721 ( .A1(n37538), .A2(n37539), .A3(n37540), .A4(n37541), .ZN(
        n37542) );
  OR4_X1 U722 ( .A1(n37528), .A2(n37533), .A3(n37537), .A4(n37542), .ZN(
        OUTB[12]) );
  AOI22_X1 U723 ( .A1(n37702), .A2(\REGISTERS[9][11] ), .B1(n37701), .B2(
        \REGISTERS[16][11] ), .ZN(n37543) );
  AOI22_X1 U724 ( .A1(n37708), .A2(\REGISTERS[23][11] ), .B1(n37710), .B2(
        \REGISTERS[6][11] ), .ZN(n37544) );
  AOI22_X1 U725 ( .A1(n37706), .A2(\REGISTERS[14][11] ), .B1(n37707), .B2(
        \REGISTERS[24][11] ), .ZN(n37545) );
  AOI22_X1 U726 ( .A1(n37704), .A2(\REGISTERS[10][11] ), .B1(n37705), .B2(
        \REGISTERS[12][11] ), .ZN(n37546) );
  NAND4_X1 U727 ( .A1(n37543), .A2(n37544), .A3(n37545), .A4(n37546), .ZN(
        n37547) );
  AOI22_X1 U728 ( .A1(n37723), .A2(\REGISTERS[27][11] ), .B1(n37703), .B2(
        \REGISTERS[1][11] ), .ZN(n37548) );
  AOI22_X1 U729 ( .A1(n37695), .A2(\REGISTERS[21][11] ), .B1(n37699), .B2(
        \REGISTERS[20][11] ), .ZN(n37549) );
  AOI22_X1 U730 ( .A1(n37698), .A2(\REGISTERS[7][11] ), .B1(n37700), .B2(
        \REGISTERS[18][11] ), .ZN(n37550) );
  AOI22_X1 U731 ( .A1(n37716), .A2(\REGISTERS[5][11] ), .B1(n37718), .B2(
        \REGISTERS[28][11] ), .ZN(n37551) );
  NAND4_X1 U732 ( .A1(n37548), .A2(n37549), .A3(n37550), .A4(n37551), .ZN(
        n37552) );
  AOI22_X1 U733 ( .A1(n37709), .A2(\REGISTERS[25][11] ), .B1(n37720), .B2(
        \REGISTERS[11][11] ), .ZN(n37553) );
  AOI22_X1 U734 ( .A1(n37725), .A2(\REGISTERS[31][11] ), .B1(n37721), .B2(
        \REGISTERS[2][11] ), .ZN(n37554) );
  AOI222_X1 U735 ( .A1(n37696), .A2(\REGISTERS[29][11] ), .B1(n37697), .B2(
        \REGISTERS[13][11] ), .C1(n37722), .C2(\REGISTERS[19][11] ), .ZN(
        n37555) );
  NAND3_X1 U736 ( .A1(n37553), .A2(n37554), .A3(n37555), .ZN(n37556) );
  AOI22_X1 U737 ( .A1(n37712), .A2(\REGISTERS[26][11] ), .B1(n37715), .B2(
        \REGISTERS[8][11] ), .ZN(n37557) );
  AOI22_X1 U738 ( .A1(n37714), .A2(\REGISTERS[30][11] ), .B1(n37711), .B2(
        \REGISTERS[3][11] ), .ZN(n37558) );
  AOI22_X1 U739 ( .A1(n37719), .A2(\REGISTERS[17][11] ), .B1(n37717), .B2(
        \REGISTERS[4][11] ), .ZN(n37559) );
  AOI22_X1 U740 ( .A1(n37713), .A2(\REGISTERS[22][11] ), .B1(n37724), .B2(
        \REGISTERS[15][11] ), .ZN(n37560) );
  NAND4_X1 U741 ( .A1(n37557), .A2(n37558), .A3(n37559), .A4(n37560), .ZN(
        n37561) );
  OR4_X1 U742 ( .A1(n37547), .A2(n37552), .A3(n37556), .A4(n37561), .ZN(
        OUTB[11]) );
  AOI22_X1 U743 ( .A1(n37702), .A2(\REGISTERS[9][10] ), .B1(n37701), .B2(
        \REGISTERS[16][10] ), .ZN(n37562) );
  AOI22_X1 U744 ( .A1(n37708), .A2(\REGISTERS[23][10] ), .B1(n37710), .B2(
        \REGISTERS[6][10] ), .ZN(n37563) );
  AOI22_X1 U745 ( .A1(n37706), .A2(\REGISTERS[14][10] ), .B1(n37707), .B2(
        \REGISTERS[24][10] ), .ZN(n37564) );
  AOI22_X1 U746 ( .A1(n37704), .A2(\REGISTERS[10][10] ), .B1(n37705), .B2(
        \REGISTERS[12][10] ), .ZN(n37565) );
  NAND4_X1 U747 ( .A1(n37562), .A2(n37563), .A3(n37564), .A4(n37565), .ZN(
        n37566) );
  AOI22_X1 U748 ( .A1(n37723), .A2(\REGISTERS[27][10] ), .B1(n37703), .B2(
        \REGISTERS[1][10] ), .ZN(n37567) );
  AOI22_X1 U749 ( .A1(n37695), .A2(\REGISTERS[21][10] ), .B1(n37699), .B2(
        \REGISTERS[20][10] ), .ZN(n37568) );
  AOI22_X1 U750 ( .A1(n37698), .A2(\REGISTERS[7][10] ), .B1(n37700), .B2(
        \REGISTERS[18][10] ), .ZN(n37569) );
  AOI22_X1 U751 ( .A1(n37716), .A2(\REGISTERS[5][10] ), .B1(n37718), .B2(
        \REGISTERS[28][10] ), .ZN(n37570) );
  NAND4_X1 U752 ( .A1(n37567), .A2(n37568), .A3(n37569), .A4(n37570), .ZN(
        n37571) );
  AOI22_X1 U753 ( .A1(n37709), .A2(\REGISTERS[25][10] ), .B1(n37720), .B2(
        \REGISTERS[11][10] ), .ZN(n37572) );
  AOI22_X1 U754 ( .A1(n37725), .A2(\REGISTERS[31][10] ), .B1(n37721), .B2(
        \REGISTERS[2][10] ), .ZN(n37573) );
  AOI222_X1 U755 ( .A1(n37696), .A2(\REGISTERS[29][10] ), .B1(n37697), .B2(
        \REGISTERS[13][10] ), .C1(n37722), .C2(\REGISTERS[19][10] ), .ZN(
        n37574) );
  NAND3_X1 U756 ( .A1(n37572), .A2(n37573), .A3(n37574), .ZN(n37575) );
  AOI22_X1 U757 ( .A1(n37712), .A2(\REGISTERS[26][10] ), .B1(n37715), .B2(
        \REGISTERS[8][10] ), .ZN(n37576) );
  AOI22_X1 U758 ( .A1(n37714), .A2(\REGISTERS[30][10] ), .B1(n37711), .B2(
        \REGISTERS[3][10] ), .ZN(n37577) );
  AOI22_X1 U759 ( .A1(n37719), .A2(\REGISTERS[17][10] ), .B1(n37717), .B2(
        \REGISTERS[4][10] ), .ZN(n37578) );
  AOI22_X1 U760 ( .A1(n37713), .A2(\REGISTERS[22][10] ), .B1(n37724), .B2(
        \REGISTERS[15][10] ), .ZN(n37579) );
  NAND4_X1 U761 ( .A1(n37576), .A2(n37577), .A3(n37578), .A4(n37579), .ZN(
        n37580) );
  OR4_X1 U762 ( .A1(n37566), .A2(n37571), .A3(n37575), .A4(n37580), .ZN(
        OUTB[10]) );
  AOI22_X1 U763 ( .A1(n37702), .A2(\REGISTERS[9][9] ), .B1(n37701), .B2(
        \REGISTERS[16][9] ), .ZN(n37581) );
  AOI22_X1 U764 ( .A1(n37708), .A2(\REGISTERS[23][9] ), .B1(n37710), .B2(
        \REGISTERS[6][9] ), .ZN(n37582) );
  AOI22_X1 U765 ( .A1(n37706), .A2(\REGISTERS[14][9] ), .B1(n37707), .B2(
        \REGISTERS[24][9] ), .ZN(n37583) );
  AOI22_X1 U766 ( .A1(n37704), .A2(\REGISTERS[10][9] ), .B1(n37705), .B2(
        \REGISTERS[12][9] ), .ZN(n37584) );
  NAND4_X1 U767 ( .A1(n37581), .A2(n37582), .A3(n37583), .A4(n37584), .ZN(
        n37585) );
  AOI22_X1 U768 ( .A1(n37723), .A2(\REGISTERS[27][9] ), .B1(n37703), .B2(
        \REGISTERS[1][9] ), .ZN(n37586) );
  AOI22_X1 U769 ( .A1(n37695), .A2(\REGISTERS[21][9] ), .B1(n37699), .B2(
        \REGISTERS[20][9] ), .ZN(n37587) );
  AOI22_X1 U770 ( .A1(n37698), .A2(\REGISTERS[7][9] ), .B1(n37700), .B2(
        \REGISTERS[18][9] ), .ZN(n37588) );
  AOI22_X1 U771 ( .A1(n37716), .A2(\REGISTERS[5][9] ), .B1(n37718), .B2(
        \REGISTERS[28][9] ), .ZN(n37589) );
  NAND4_X1 U772 ( .A1(n37586), .A2(n37587), .A3(n37588), .A4(n37589), .ZN(
        n37590) );
  AOI22_X1 U773 ( .A1(n37709), .A2(\REGISTERS[25][9] ), .B1(n37720), .B2(
        \REGISTERS[11][9] ), .ZN(n37591) );
  AOI22_X1 U774 ( .A1(n37725), .A2(\REGISTERS[31][9] ), .B1(n37721), .B2(
        \REGISTERS[2][9] ), .ZN(n37592) );
  AOI222_X1 U775 ( .A1(n37696), .A2(\REGISTERS[29][9] ), .B1(n37697), .B2(
        \REGISTERS[13][9] ), .C1(n37722), .C2(\REGISTERS[19][9] ), .ZN(n37593)
         );
  NAND3_X1 U776 ( .A1(n37591), .A2(n37592), .A3(n37593), .ZN(n37594) );
  AOI22_X1 U777 ( .A1(n37712), .A2(\REGISTERS[26][9] ), .B1(n37715), .B2(
        \REGISTERS[8][9] ), .ZN(n37595) );
  AOI22_X1 U778 ( .A1(n37714), .A2(\REGISTERS[30][9] ), .B1(n37711), .B2(
        \REGISTERS[3][9] ), .ZN(n37596) );
  AOI22_X1 U779 ( .A1(n37719), .A2(\REGISTERS[17][9] ), .B1(n37717), .B2(
        \REGISTERS[4][9] ), .ZN(n37597) );
  AOI22_X1 U780 ( .A1(n37713), .A2(\REGISTERS[22][9] ), .B1(n37724), .B2(
        \REGISTERS[15][9] ), .ZN(n37598) );
  NAND4_X1 U781 ( .A1(n37595), .A2(n37596), .A3(n37597), .A4(n37598), .ZN(
        n37599) );
  OR4_X1 U782 ( .A1(n37585), .A2(n37590), .A3(n37594), .A4(n37599), .ZN(
        OUTB[9]) );
  AOI22_X1 U783 ( .A1(n37702), .A2(\REGISTERS[9][8] ), .B1(n37701), .B2(
        \REGISTERS[16][8] ), .ZN(n37600) );
  AOI22_X1 U784 ( .A1(n37708), .A2(\REGISTERS[23][8] ), .B1(n37710), .B2(
        \REGISTERS[6][8] ), .ZN(n37601) );
  AOI22_X1 U785 ( .A1(n37706), .A2(\REGISTERS[14][8] ), .B1(n37707), .B2(
        \REGISTERS[24][8] ), .ZN(n37602) );
  AOI22_X1 U786 ( .A1(n37704), .A2(\REGISTERS[10][8] ), .B1(n37705), .B2(
        \REGISTERS[12][8] ), .ZN(n37603) );
  NAND4_X1 U787 ( .A1(n37600), .A2(n37601), .A3(n37602), .A4(n37603), .ZN(
        n37604) );
  AOI22_X1 U788 ( .A1(n37723), .A2(\REGISTERS[27][8] ), .B1(n37703), .B2(
        \REGISTERS[1][8] ), .ZN(n37605) );
  AOI22_X1 U789 ( .A1(n37695), .A2(\REGISTERS[21][8] ), .B1(n37699), .B2(
        \REGISTERS[20][8] ), .ZN(n37606) );
  AOI22_X1 U790 ( .A1(n37698), .A2(\REGISTERS[7][8] ), .B1(n37700), .B2(
        \REGISTERS[18][8] ), .ZN(n37607) );
  AOI22_X1 U791 ( .A1(n37716), .A2(\REGISTERS[5][8] ), .B1(n37718), .B2(
        \REGISTERS[28][8] ), .ZN(n37608) );
  NAND4_X1 U792 ( .A1(n37605), .A2(n37606), .A3(n37607), .A4(n37608), .ZN(
        n37609) );
  AOI22_X1 U793 ( .A1(n37709), .A2(\REGISTERS[25][8] ), .B1(n37720), .B2(
        \REGISTERS[11][8] ), .ZN(n37610) );
  AOI22_X1 U794 ( .A1(n37725), .A2(\REGISTERS[31][8] ), .B1(n37721), .B2(
        \REGISTERS[2][8] ), .ZN(n37611) );
  AOI222_X1 U795 ( .A1(n37696), .A2(\REGISTERS[29][8] ), .B1(n37697), .B2(
        \REGISTERS[13][8] ), .C1(n37722), .C2(\REGISTERS[19][8] ), .ZN(n37612)
         );
  NAND3_X1 U796 ( .A1(n37610), .A2(n37611), .A3(n37612), .ZN(n37613) );
  AOI22_X1 U797 ( .A1(n37712), .A2(\REGISTERS[26][8] ), .B1(n37715), .B2(
        \REGISTERS[8][8] ), .ZN(n37614) );
  AOI22_X1 U798 ( .A1(n37714), .A2(\REGISTERS[30][8] ), .B1(n37711), .B2(
        \REGISTERS[3][8] ), .ZN(n37615) );
  AOI22_X1 U799 ( .A1(n37719), .A2(\REGISTERS[17][8] ), .B1(n37717), .B2(
        \REGISTERS[4][8] ), .ZN(n37616) );
  AOI22_X1 U800 ( .A1(n37713), .A2(\REGISTERS[22][8] ), .B1(n37724), .B2(
        \REGISTERS[15][8] ), .ZN(n37617) );
  NAND4_X1 U801 ( .A1(n37614), .A2(n37615), .A3(n37616), .A4(n37617), .ZN(
        n37618) );
  OR4_X1 U802 ( .A1(n37604), .A2(n37609), .A3(n37613), .A4(n37618), .ZN(
        OUTB[8]) );
  AOI22_X1 U803 ( .A1(n37702), .A2(\REGISTERS[9][3] ), .B1(n37701), .B2(
        \REGISTERS[16][3] ), .ZN(n37619) );
  AOI22_X1 U804 ( .A1(n37708), .A2(\REGISTERS[23][3] ), .B1(n37710), .B2(
        \REGISTERS[6][3] ), .ZN(n37620) );
  AOI22_X1 U805 ( .A1(n37706), .A2(\REGISTERS[14][3] ), .B1(n37707), .B2(
        \REGISTERS[24][3] ), .ZN(n37621) );
  AOI22_X1 U806 ( .A1(n37704), .A2(\REGISTERS[10][3] ), .B1(n37705), .B2(
        \REGISTERS[12][3] ), .ZN(n37622) );
  NAND4_X1 U807 ( .A1(n37619), .A2(n37620), .A3(n37621), .A4(n37622), .ZN(
        n37623) );
  AOI22_X1 U808 ( .A1(n37723), .A2(\REGISTERS[27][3] ), .B1(n37703), .B2(
        \REGISTERS[1][3] ), .ZN(n37624) );
  AOI22_X1 U809 ( .A1(n37695), .A2(\REGISTERS[21][3] ), .B1(n37699), .B2(
        \REGISTERS[20][3] ), .ZN(n37625) );
  AOI22_X1 U810 ( .A1(n37698), .A2(\REGISTERS[7][3] ), .B1(n37700), .B2(
        \REGISTERS[18][3] ), .ZN(n37626) );
  AOI22_X1 U811 ( .A1(n37716), .A2(\REGISTERS[5][3] ), .B1(n37718), .B2(
        \REGISTERS[28][3] ), .ZN(n37627) );
  NAND4_X1 U812 ( .A1(n37624), .A2(n37625), .A3(n37626), .A4(n37627), .ZN(
        n37628) );
  AOI22_X1 U813 ( .A1(n37709), .A2(\REGISTERS[25][3] ), .B1(n37720), .B2(
        \REGISTERS[11][3] ), .ZN(n37629) );
  AOI22_X1 U814 ( .A1(n38277), .A2(\REGISTERS[31][3] ), .B1(n38278), .B2(
        \REGISTERS[2][3] ), .ZN(n37630) );
  AOI222_X1 U815 ( .A1(n37696), .A2(\REGISTERS[29][3] ), .B1(n37697), .B2(
        \REGISTERS[13][3] ), .C1(n37722), .C2(\REGISTERS[19][3] ), .ZN(n37631)
         );
  NAND3_X1 U816 ( .A1(n37629), .A2(n37630), .A3(n37631), .ZN(n37632) );
  AOI22_X1 U817 ( .A1(n37712), .A2(\REGISTERS[26][3] ), .B1(n37715), .B2(
        \REGISTERS[8][3] ), .ZN(n37633) );
  AOI22_X1 U818 ( .A1(n37714), .A2(\REGISTERS[30][3] ), .B1(n37711), .B2(
        \REGISTERS[3][3] ), .ZN(n37634) );
  AOI22_X1 U819 ( .A1(n37719), .A2(\REGISTERS[17][3] ), .B1(n37717), .B2(
        \REGISTERS[4][3] ), .ZN(n37635) );
  AOI22_X1 U820 ( .A1(n37713), .A2(\REGISTERS[22][3] ), .B1(n38289), .B2(
        \REGISTERS[15][3] ), .ZN(n37636) );
  NAND4_X1 U821 ( .A1(n37633), .A2(n37634), .A3(n37635), .A4(n37636), .ZN(
        n37637) );
  OR4_X1 U822 ( .A1(n37623), .A2(n37628), .A3(n37632), .A4(n37637), .ZN(
        OUTB[3]) );
  AOI22_X1 U823 ( .A1(n37702), .A2(\REGISTERS[9][2] ), .B1(n37701), .B2(
        \REGISTERS[16][2] ), .ZN(n37638) );
  AOI22_X1 U824 ( .A1(n37708), .A2(\REGISTERS[23][2] ), .B1(n37710), .B2(
        \REGISTERS[6][2] ), .ZN(n37639) );
  AOI22_X1 U825 ( .A1(n37706), .A2(\REGISTERS[14][2] ), .B1(n37707), .B2(
        \REGISTERS[24][2] ), .ZN(n37640) );
  AOI22_X1 U826 ( .A1(n37704), .A2(\REGISTERS[10][2] ), .B1(n37705), .B2(
        \REGISTERS[12][2] ), .ZN(n37641) );
  NAND4_X1 U827 ( .A1(n37638), .A2(n37639), .A3(n37640), .A4(n37641), .ZN(
        n37642) );
  AOI22_X1 U828 ( .A1(n37723), .A2(\REGISTERS[27][2] ), .B1(n37703), .B2(
        \REGISTERS[1][2] ), .ZN(n37643) );
  AOI22_X1 U829 ( .A1(n37695), .A2(\REGISTERS[21][2] ), .B1(n37699), .B2(
        \REGISTERS[20][2] ), .ZN(n37644) );
  AOI22_X1 U830 ( .A1(n37698), .A2(\REGISTERS[7][2] ), .B1(n37700), .B2(
        \REGISTERS[18][2] ), .ZN(n37645) );
  AOI22_X1 U831 ( .A1(n37716), .A2(\REGISTERS[5][2] ), .B1(n37718), .B2(
        \REGISTERS[28][2] ), .ZN(n37646) );
  NAND4_X1 U832 ( .A1(n37643), .A2(n37644), .A3(n37645), .A4(n37646), .ZN(
        n37647) );
  AOI22_X1 U833 ( .A1(n37709), .A2(\REGISTERS[25][2] ), .B1(n37720), .B2(
        \REGISTERS[11][2] ), .ZN(n37648) );
  AOI22_X1 U834 ( .A1(n37725), .A2(\REGISTERS[31][2] ), .B1(n37721), .B2(
        \REGISTERS[2][2] ), .ZN(n37649) );
  AOI222_X1 U835 ( .A1(n37696), .A2(\REGISTERS[29][2] ), .B1(n37697), .B2(
        \REGISTERS[13][2] ), .C1(n37722), .C2(\REGISTERS[19][2] ), .ZN(n37650)
         );
  NAND3_X1 U836 ( .A1(n37648), .A2(n37649), .A3(n37650), .ZN(n37651) );
  AOI22_X1 U837 ( .A1(n37712), .A2(\REGISTERS[26][2] ), .B1(n37715), .B2(
        \REGISTERS[8][2] ), .ZN(n37652) );
  AOI22_X1 U838 ( .A1(n37714), .A2(\REGISTERS[30][2] ), .B1(n37711), .B2(
        \REGISTERS[3][2] ), .ZN(n37653) );
  AOI22_X1 U839 ( .A1(n37719), .A2(\REGISTERS[17][2] ), .B1(n37717), .B2(
        \REGISTERS[4][2] ), .ZN(n37654) );
  AOI22_X1 U840 ( .A1(n37713), .A2(\REGISTERS[22][2] ), .B1(n37724), .B2(
        \REGISTERS[15][2] ), .ZN(n37655) );
  NAND4_X1 U841 ( .A1(n37652), .A2(n37653), .A3(n37654), .A4(n37655), .ZN(
        n37656) );
  OR4_X1 U842 ( .A1(n37642), .A2(n37647), .A3(n37651), .A4(n37656), .ZN(
        OUTB[2]) );
  AOI22_X1 U843 ( .A1(n37702), .A2(\REGISTERS[9][1] ), .B1(n37701), .B2(
        \REGISTERS[16][1] ), .ZN(n37657) );
  AOI22_X1 U844 ( .A1(n37708), .A2(\REGISTERS[23][1] ), .B1(n37710), .B2(
        \REGISTERS[6][1] ), .ZN(n37658) );
  AOI22_X1 U845 ( .A1(n37706), .A2(\REGISTERS[14][1] ), .B1(n37707), .B2(
        \REGISTERS[24][1] ), .ZN(n37659) );
  AOI22_X1 U846 ( .A1(n37704), .A2(\REGISTERS[10][1] ), .B1(n37705), .B2(
        \REGISTERS[12][1] ), .ZN(n37660) );
  NAND4_X1 U847 ( .A1(n37657), .A2(n37658), .A3(n37659), .A4(n37660), .ZN(
        n37661) );
  AOI22_X1 U848 ( .A1(n37723), .A2(\REGISTERS[27][1] ), .B1(n37703), .B2(
        \REGISTERS[1][1] ), .ZN(n37662) );
  AOI22_X1 U849 ( .A1(n37695), .A2(\REGISTERS[21][1] ), .B1(n37699), .B2(
        \REGISTERS[20][1] ), .ZN(n37663) );
  AOI22_X1 U850 ( .A1(n37698), .A2(\REGISTERS[7][1] ), .B1(n37700), .B2(
        \REGISTERS[18][1] ), .ZN(n37664) );
  AOI22_X1 U851 ( .A1(n37716), .A2(\REGISTERS[5][1] ), .B1(n37718), .B2(
        \REGISTERS[28][1] ), .ZN(n37665) );
  NAND4_X1 U852 ( .A1(n37662), .A2(n37663), .A3(n37664), .A4(n37665), .ZN(
        n37666) );
  AOI22_X1 U853 ( .A1(n37709), .A2(\REGISTERS[25][1] ), .B1(n37720), .B2(
        \REGISTERS[11][1] ), .ZN(n37667) );
  AOI22_X1 U854 ( .A1(n37725), .A2(\REGISTERS[31][1] ), .B1(n37721), .B2(
        \REGISTERS[2][1] ), .ZN(n37668) );
  AOI222_X1 U855 ( .A1(n37696), .A2(\REGISTERS[29][1] ), .B1(n37697), .B2(
        \REGISTERS[13][1] ), .C1(n37722), .C2(\REGISTERS[19][1] ), .ZN(n37669)
         );
  NAND3_X1 U856 ( .A1(n37667), .A2(n37668), .A3(n37669), .ZN(n37670) );
  AOI22_X1 U857 ( .A1(n37712), .A2(\REGISTERS[26][1] ), .B1(n37715), .B2(
        \REGISTERS[8][1] ), .ZN(n37671) );
  AOI22_X1 U858 ( .A1(n37714), .A2(\REGISTERS[30][1] ), .B1(n37711), .B2(
        \REGISTERS[3][1] ), .ZN(n37672) );
  AOI22_X1 U859 ( .A1(n37719), .A2(\REGISTERS[17][1] ), .B1(n37717), .B2(
        \REGISTERS[4][1] ), .ZN(n37673) );
  AOI22_X1 U860 ( .A1(n37713), .A2(\REGISTERS[22][1] ), .B1(n37724), .B2(
        \REGISTERS[15][1] ), .ZN(n37674) );
  NAND4_X1 U861 ( .A1(n37671), .A2(n37672), .A3(n37673), .A4(n37674), .ZN(
        n37675) );
  OR4_X1 U862 ( .A1(n37661), .A2(n37666), .A3(n37670), .A4(n37675), .ZN(
        OUTB[1]) );
  AOI22_X1 U863 ( .A1(n37702), .A2(\REGISTERS[9][0] ), .B1(n37701), .B2(
        \REGISTERS[16][0] ), .ZN(n37676) );
  AOI22_X1 U864 ( .A1(n37708), .A2(\REGISTERS[23][0] ), .B1(n37710), .B2(
        \REGISTERS[6][0] ), .ZN(n37677) );
  AOI22_X1 U865 ( .A1(n37706), .A2(\REGISTERS[14][0] ), .B1(n37707), .B2(
        \REGISTERS[24][0] ), .ZN(n37678) );
  AOI22_X1 U866 ( .A1(n37704), .A2(\REGISTERS[10][0] ), .B1(n37705), .B2(
        \REGISTERS[12][0] ), .ZN(n37679) );
  NAND4_X1 U867 ( .A1(n37676), .A2(n37677), .A3(n37678), .A4(n37679), .ZN(
        n37680) );
  AOI22_X1 U868 ( .A1(n37723), .A2(\REGISTERS[27][0] ), .B1(n37703), .B2(
        \REGISTERS[1][0] ), .ZN(n37681) );
  AOI22_X1 U869 ( .A1(n37695), .A2(\REGISTERS[21][0] ), .B1(n37699), .B2(
        \REGISTERS[20][0] ), .ZN(n37682) );
  AOI22_X1 U870 ( .A1(n37698), .A2(\REGISTERS[7][0] ), .B1(n37700), .B2(
        \REGISTERS[18][0] ), .ZN(n37683) );
  AOI22_X1 U871 ( .A1(n37716), .A2(\REGISTERS[5][0] ), .B1(n37718), .B2(
        \REGISTERS[28][0] ), .ZN(n37684) );
  NAND4_X1 U872 ( .A1(n37681), .A2(n37682), .A3(n37683), .A4(n37684), .ZN(
        n37685) );
  AOI22_X1 U873 ( .A1(n37709), .A2(\REGISTERS[25][0] ), .B1(n37720), .B2(
        \REGISTERS[11][0] ), .ZN(n37686) );
  AOI22_X1 U874 ( .A1(n37725), .A2(\REGISTERS[31][0] ), .B1(n37721), .B2(
        \REGISTERS[2][0] ), .ZN(n37687) );
  AOI222_X1 U875 ( .A1(n37696), .A2(\REGISTERS[29][0] ), .B1(n37697), .B2(
        \REGISTERS[13][0] ), .C1(n37722), .C2(\REGISTERS[19][0] ), .ZN(n37688)
         );
  NAND3_X1 U876 ( .A1(n37686), .A2(n37687), .A3(n37688), .ZN(n37689) );
  AOI22_X1 U877 ( .A1(n37712), .A2(\REGISTERS[26][0] ), .B1(n37715), .B2(
        \REGISTERS[8][0] ), .ZN(n37690) );
  AOI22_X1 U878 ( .A1(n37714), .A2(\REGISTERS[30][0] ), .B1(n37711), .B2(
        \REGISTERS[3][0] ), .ZN(n37691) );
  AOI22_X1 U879 ( .A1(n37719), .A2(\REGISTERS[17][0] ), .B1(n37717), .B2(
        \REGISTERS[4][0] ), .ZN(n37692) );
  AOI22_X1 U880 ( .A1(n37713), .A2(\REGISTERS[22][0] ), .B1(n37724), .B2(
        \REGISTERS[15][0] ), .ZN(n37693) );
  NAND4_X1 U881 ( .A1(n37690), .A2(n37691), .A3(n37692), .A4(n37693), .ZN(
        n37694) );
  OR4_X1 U882 ( .A1(n37680), .A2(n37685), .A3(n37689), .A4(n37694), .ZN(
        OUTB[0]) );
  BUF_X2 U883 ( .A(n38300), .Z(n37695) );
  BUF_X2 U884 ( .A(n38279), .Z(n37696) );
  BUF_X2 U885 ( .A(n38280), .Z(n37697) );
  BUF_X2 U886 ( .A(n38302), .Z(n37698) );
  BUF_X2 U887 ( .A(n38301), .Z(n37699) );
  BUF_X2 U888 ( .A(n38303), .Z(n37700) );
  BUF_X2 U889 ( .A(n38291), .Z(n37701) );
  BUF_X2 U890 ( .A(n38290), .Z(n37702) );
  BUF_X2 U891 ( .A(n38299), .Z(n37703) );
  BUF_X2 U892 ( .A(n38296), .Z(n37704) );
  BUF_X2 U893 ( .A(n38297), .Z(n37705) );
  BUF_X2 U894 ( .A(n38294), .Z(n37706) );
  BUF_X2 U895 ( .A(n38295), .Z(n37707) );
  BUF_X2 U896 ( .A(n38292), .Z(n37708) );
  BUF_X2 U897 ( .A(n38275), .Z(n37709) );
  BUF_X2 U898 ( .A(n38293), .Z(n37710) );
  BUF_X2 U899 ( .A(n38285), .Z(n37711) );
  BUF_X2 U900 ( .A(n38282), .Z(n37712) );
  BUF_X2 U901 ( .A(n38288), .Z(n37713) );
  BUF_X2 U902 ( .A(n38284), .Z(n37714) );
  BUF_X2 U903 ( .A(n38283), .Z(n37715) );
  BUF_X2 U904 ( .A(n38304), .Z(n37716) );
  BUF_X2 U905 ( .A(n38287), .Z(n37717) );
  BUF_X2 U906 ( .A(n38305), .Z(n37718) );
  BUF_X2 U907 ( .A(n38286), .Z(n37719) );
  BUF_X2 U908 ( .A(n38276), .Z(n37720) );
  BUF_X2 U909 ( .A(n38278), .Z(n37721) );
  BUF_X2 U910 ( .A(n38281), .Z(n37722) );
  BUF_X2 U911 ( .A(n38298), .Z(n37723) );
  BUF_X2 U912 ( .A(n38289), .Z(n37724) );
  BUF_X2 U913 ( .A(n38277), .Z(n37725) );
  NOR3_X2 U914 ( .A1(ADD_RDA[2]), .A2(n37811), .A3(n37813), .ZN(n38221) );
  BUF_X1 U915 ( .A(n38230), .Z(n37743) );
  BUF_X1 U916 ( .A(n38221), .Z(n37738) );
  BUF_X1 U917 ( .A(n38231), .Z(n37744) );
  BUF_X1 U918 ( .A(n38218), .Z(n37735) );
  BUF_X1 U919 ( .A(n38246), .Z(n37755) );
  BUF_X1 U920 ( .A(n38243), .Z(n37752) );
  BUF_X1 U921 ( .A(n38241), .Z(n37750) );
  BUF_X1 U922 ( .A(n38210), .Z(n37731) );
  BUF_X1 U923 ( .A(n38208), .Z(n37729) );
  BUF_X1 U924 ( .A(n38206), .Z(n37727) );
  BUF_X1 U925 ( .A(n38240), .Z(n37749) );
  BUF_X1 U926 ( .A(n38232), .Z(n37745) );
  BUF_X1 U927 ( .A(n38228), .Z(n37741) );
  BUF_X1 U928 ( .A(n38211), .Z(n37732) );
  BUF_X1 U929 ( .A(n38247), .Z(n37756) );
  BUF_X1 U930 ( .A(n38245), .Z(n37754) );
  BUF_X1 U931 ( .A(n38235), .Z(n37748) );
  BUF_X1 U932 ( .A(n38233), .Z(n37746) );
  BUF_X1 U933 ( .A(n38229), .Z(n37742) );
  BUF_X1 U934 ( .A(n38223), .Z(n37740) );
  BUF_X1 U935 ( .A(n38219), .Z(n37736) );
  BUF_X1 U936 ( .A(n38217), .Z(n37734) );
  BUF_X1 U937 ( .A(n38209), .Z(n37730) );
  BUF_X1 U938 ( .A(n38234), .Z(n37747) );
  BUF_X1 U939 ( .A(n38222), .Z(n37739) );
  BUF_X1 U940 ( .A(n38244), .Z(n37753) );
  BUF_X1 U941 ( .A(n38242), .Z(n37751) );
  BUF_X1 U942 ( .A(n38220), .Z(n37737) );
  BUF_X1 U943 ( .A(n38216), .Z(n37733) );
  BUF_X1 U944 ( .A(n38207), .Z(n37728) );
  BUF_X1 U945 ( .A(n38205), .Z(n37726) );
  INV_X1 U946 ( .A(ADD_RDA[1]), .ZN(n37811) );
  INV_X1 U947 ( .A(ADD_RDA[3]), .ZN(n37817) );
  INV_X1 U948 ( .A(ADD_RDA[2]), .ZN(n37812) );
  OR4_X1 U949 ( .A1(n38184), .A2(n38183), .A3(n38182), .A4(n38181), .ZN(
        OUTA[6]) );
  OR4_X1 U950 ( .A1(n38144), .A2(n38143), .A3(n38142), .A4(n38141), .ZN(
        OUTA[3]) );
  OR4_X1 U951 ( .A1(n38164), .A2(n38163), .A3(n38162), .A4(n38161), .ZN(
        OUTA[5]) );
  OR4_X1 U952 ( .A1(n38124), .A2(n38123), .A3(n38122), .A4(n38121), .ZN(
        OUTA[31]) );
  OR4_X1 U953 ( .A1(n38104), .A2(n38103), .A3(n38102), .A4(n38101), .ZN(
        OUTA[30]) );
  OR4_X1 U954 ( .A1(n37924), .A2(n37923), .A3(n37922), .A4(n37921), .ZN(
        OUTA[22]) );
  OR4_X1 U955 ( .A1(n37984), .A2(n37983), .A3(n37982), .A4(n37981), .ZN(
        OUTA[25]) );
  OR4_X1 U956 ( .A1(n37964), .A2(n37963), .A3(n37962), .A4(n37961), .ZN(
        OUTA[24]) );
  OR4_X1 U957 ( .A1(n37864), .A2(n37863), .A3(n37862), .A4(n37861), .ZN(
        OUTA[19]) );
  OR4_X1 U958 ( .A1(n37884), .A2(n37883), .A3(n37882), .A4(n37881), .ZN(
        OUTA[20]) );
  OR4_X1 U959 ( .A1(n37844), .A2(n37843), .A3(n37842), .A4(n37841), .ZN(
        OUTA[18]) );
  OR4_X1 U960 ( .A1(n37944), .A2(n37943), .A3(n37942), .A4(n37941), .ZN(
        OUTA[23]) );
  OR4_X1 U961 ( .A1(n37904), .A2(n37903), .A3(n37902), .A4(n37901), .ZN(
        OUTA[21]) );
  OR4_X1 U962 ( .A1(n38024), .A2(n38023), .A3(n38022), .A4(n38021), .ZN(
        OUTA[27]) );
  OR4_X1 U963 ( .A1(n38204), .A2(n38203), .A3(n38202), .A4(n38201), .ZN(
        OUTA[8]) );
  OR4_X1 U964 ( .A1(n38084), .A2(n38083), .A3(n38082), .A4(n38081), .ZN(
        OUTA[2]) );
  OR4_X1 U965 ( .A1(n38064), .A2(n38063), .A3(n38062), .A4(n38061), .ZN(
        OUTA[29]) );
  OR4_X1 U966 ( .A1(n38004), .A2(n38003), .A3(n38002), .A4(n38001), .ZN(
        OUTA[26]) );
  OR4_X1 U967 ( .A1(n38255), .A2(n38254), .A3(n38253), .A4(n38252), .ZN(
        OUTA[9]) );
  OR4_X1 U968 ( .A1(n38044), .A2(n38043), .A3(n38042), .A4(n38041), .ZN(
        OUTA[28]) );
  NOR2_X1 U969 ( .A1(n37809), .A2(n37818), .ZN(n38211) );
  BUF_X1 U970 ( .A(N291), .Z(n37771) );
  BUF_X1 U971 ( .A(N290), .Z(n37772) );
  BUF_X1 U972 ( .A(N292), .Z(n37770) );
  BUF_X1 U973 ( .A(N293), .Z(n37769) );
  BUF_X1 U974 ( .A(N294), .Z(n37768) );
  BUF_X1 U975 ( .A(N285), .Z(n37777) );
  BUF_X1 U976 ( .A(N284), .Z(n37778) );
  BUF_X1 U977 ( .A(N286), .Z(n37776) );
  BUF_X1 U978 ( .A(N287), .Z(n37775) );
  BUF_X1 U979 ( .A(N288), .Z(n37774) );
  BUF_X1 U980 ( .A(N289), .Z(n37773) );
  BUF_X1 U981 ( .A(N302), .Z(n37760) );
  BUF_X1 U982 ( .A(N303), .Z(n37759) );
  BUF_X1 U983 ( .A(N304), .Z(n37758) );
  BUF_X1 U984 ( .A(N305), .Z(n37757) );
  BUF_X1 U985 ( .A(N295), .Z(n37767) );
  BUF_X1 U986 ( .A(N296), .Z(n37766) );
  BUF_X1 U987 ( .A(N297), .Z(n37765) );
  BUF_X1 U988 ( .A(N298), .Z(n37764) );
  BUF_X1 U989 ( .A(N299), .Z(n37763) );
  BUF_X1 U990 ( .A(N300), .Z(n37762) );
  BUF_X1 U991 ( .A(N301), .Z(n37761) );
  BUF_X1 U992 ( .A(N281), .Z(n37781) );
  BUF_X1 U993 ( .A(N279), .Z(n37783) );
  BUF_X1 U994 ( .A(N243), .Z(n37787) );
  BUF_X1 U995 ( .A(N280), .Z(n37782) );
  BUF_X1 U996 ( .A(N278), .Z(n37784) );
  BUF_X1 U997 ( .A(N283), .Z(n37779) );
  BUF_X1 U998 ( .A(N276), .Z(n37786) );
  BUF_X1 U999 ( .A(N282), .Z(n37780) );
  INV_X1 U1000 ( .A(ADD_WR[0]), .ZN(n37790) );
  BUF_X1 U1001 ( .A(N277), .Z(n37785) );
  AND2_X1 U1002 ( .A1(RESET), .A2(DATAIN[0]), .ZN(N244) );
  AND2_X1 U1003 ( .A1(RESET), .A2(DATAIN[31]), .ZN(N275) );
  AND2_X1 U1004 ( .A1(RESET), .A2(DATAIN[1]), .ZN(N245) );
  AND2_X1 U1005 ( .A1(RESET), .A2(DATAIN[30]), .ZN(N274) );
  AND2_X1 U1006 ( .A1(RESET), .A2(DATAIN[29]), .ZN(N273) );
  AND2_X1 U1007 ( .A1(RESET), .A2(DATAIN[2]), .ZN(N246) );
  AND2_X1 U1008 ( .A1(RESET), .A2(DATAIN[28]), .ZN(N272) );
  AND2_X1 U1009 ( .A1(RESET), .A2(DATAIN[27]), .ZN(N271) );
  AND2_X1 U1010 ( .A1(RESET), .A2(DATAIN[3]), .ZN(N247) );
  AND2_X1 U1011 ( .A1(RESET), .A2(DATAIN[26]), .ZN(N270) );
  AND2_X1 U1012 ( .A1(RESET), .A2(DATAIN[25]), .ZN(N269) );
  AND2_X1 U1013 ( .A1(RESET), .A2(DATAIN[4]), .ZN(N248) );
  AND2_X1 U1014 ( .A1(RESET), .A2(DATAIN[24]), .ZN(N268) );
  AND2_X1 U1015 ( .A1(RESET), .A2(DATAIN[23]), .ZN(N267) );
  AND2_X1 U1016 ( .A1(RESET), .A2(DATAIN[5]), .ZN(N249) );
  AND2_X1 U1017 ( .A1(RESET), .A2(DATAIN[22]), .ZN(N266) );
  AND2_X1 U1018 ( .A1(RESET), .A2(DATAIN[21]), .ZN(N265) );
  AND2_X1 U1019 ( .A1(RESET), .A2(DATAIN[6]), .ZN(N250) );
  AND2_X1 U1020 ( .A1(RESET), .A2(DATAIN[20]), .ZN(N264) );
  AND2_X1 U1021 ( .A1(RESET), .A2(DATAIN[19]), .ZN(N263) );
  AND2_X1 U1022 ( .A1(RESET), .A2(DATAIN[7]), .ZN(N251) );
  AND2_X1 U1023 ( .A1(RESET), .A2(DATAIN[18]), .ZN(N262) );
  AND2_X1 U1024 ( .A1(RESET), .A2(DATAIN[17]), .ZN(N261) );
  AND2_X1 U1025 ( .A1(RESET), .A2(DATAIN[8]), .ZN(N252) );
  AND2_X1 U1026 ( .A1(RESET), .A2(DATAIN[15]), .ZN(N259) );
  AND2_X1 U1027 ( .A1(RESET), .A2(DATAIN[9]), .ZN(N253) );
  AND2_X1 U1028 ( .A1(RESET), .A2(DATAIN[16]), .ZN(N260) );
  AND2_X1 U1029 ( .A1(RESET), .A2(DATAIN[14]), .ZN(N258) );
  AND2_X1 U1030 ( .A1(RESET), .A2(DATAIN[10]), .ZN(N254) );
  AND2_X1 U1031 ( .A1(RESET), .A2(DATAIN[13]), .ZN(N257) );
  AND2_X1 U1032 ( .A1(RESET), .A2(DATAIN[11]), .ZN(N255) );
  AND2_X1 U1033 ( .A1(RESET), .A2(DATAIN[12]), .ZN(N256) );
  NOR2_X1 U1034 ( .A1(n38262), .A2(n38271), .ZN(n38289) );
  NOR2_X1 U1035 ( .A1(n38267), .A2(n38271), .ZN(n38277) );
  NAND3_X1 U1036 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(ADD_WR[2]), .ZN(n37798)
         );
  NAND3_X1 U1037 ( .A1(WE), .A2(ADD_WR[3]), .A3(ADD_WR[4]), .ZN(n37792) );
  OAI21_X1 U1038 ( .B1(n37798), .B2(n37792), .A(RESET), .ZN(N243) );
  NAND3_X1 U1039 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n37790), .ZN(n37799) );
  OAI21_X1 U1040 ( .B1(n37792), .B2(n37799), .A(RESET), .ZN(N276) );
  INV_X1 U1041 ( .A(ADD_WR[1]), .ZN(n37788) );
  NAND3_X1 U1042 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n37788), .ZN(n37800) );
  OAI21_X1 U1043 ( .B1(n37792), .B2(n37800), .A(RESET), .ZN(N277) );
  NAND3_X1 U1044 ( .A1(ADD_WR[2]), .A2(n37790), .A3(n37788), .ZN(n37801) );
  OAI21_X1 U1045 ( .B1(n37792), .B2(n37801), .A(RESET), .ZN(N278) );
  NOR2_X1 U1046 ( .A1(ADD_WR[2]), .A2(n37788), .ZN(n37789) );
  NAND2_X1 U1047 ( .A1(ADD_WR[0]), .A2(n37789), .ZN(n37802) );
  OAI21_X1 U1048 ( .B1(n37792), .B2(n37802), .A(RESET), .ZN(N279) );
  NAND2_X1 U1049 ( .A1(n37789), .A2(n37790), .ZN(n37803) );
  OAI21_X1 U1050 ( .B1(n37792), .B2(n37803), .A(RESET), .ZN(N280) );
  NOR2_X1 U1051 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .ZN(n37791) );
  NAND2_X1 U1052 ( .A1(ADD_WR[0]), .A2(n37791), .ZN(n37805) );
  OAI21_X1 U1053 ( .B1(n37792), .B2(n37805), .A(RESET), .ZN(N281) );
  NAND2_X1 U1054 ( .A1(n37791), .A2(n37790), .ZN(n37795) );
  OAI21_X1 U1055 ( .B1(n37792), .B2(n37795), .A(RESET), .ZN(N282) );
  INV_X1 U1056 ( .A(ADD_WR[3]), .ZN(n37797) );
  NAND3_X1 U1057 ( .A1(WE), .A2(ADD_WR[4]), .A3(n37797), .ZN(n37793) );
  OAI21_X1 U1058 ( .B1(n37798), .B2(n37793), .A(RESET), .ZN(N283) );
  OAI21_X1 U1059 ( .B1(n37799), .B2(n37793), .A(RESET), .ZN(N284) );
  OAI21_X1 U1060 ( .B1(n37800), .B2(n37793), .A(RESET), .ZN(N285) );
  OAI21_X1 U1061 ( .B1(n37801), .B2(n37793), .A(RESET), .ZN(N286) );
  OAI21_X1 U1062 ( .B1(n37802), .B2(n37793), .A(RESET), .ZN(N287) );
  OAI21_X1 U1063 ( .B1(n37803), .B2(n37793), .A(RESET), .ZN(N288) );
  OAI21_X1 U1064 ( .B1(n37805), .B2(n37793), .A(RESET), .ZN(N289) );
  OAI21_X1 U1065 ( .B1(n37795), .B2(n37793), .A(RESET), .ZN(N290) );
  INV_X1 U1066 ( .A(ADD_WR[4]), .ZN(n37796) );
  NAND3_X1 U1067 ( .A1(ADD_WR[3]), .A2(WE), .A3(n37796), .ZN(n37794) );
  OAI21_X1 U1068 ( .B1(n37798), .B2(n37794), .A(RESET), .ZN(N291) );
  OAI21_X1 U1069 ( .B1(n37799), .B2(n37794), .A(RESET), .ZN(N292) );
  OAI21_X1 U1070 ( .B1(n37800), .B2(n37794), .A(RESET), .ZN(N293) );
  OAI21_X1 U1071 ( .B1(n37801), .B2(n37794), .A(RESET), .ZN(N294) );
  OAI21_X1 U1072 ( .B1(n37802), .B2(n37794), .A(RESET), .ZN(N295) );
  OAI21_X1 U1073 ( .B1(n37803), .B2(n37794), .A(RESET), .ZN(N296) );
  OAI21_X1 U1074 ( .B1(n37805), .B2(n37794), .A(RESET), .ZN(N297) );
  OAI21_X1 U1075 ( .B1(n37795), .B2(n37794), .A(RESET), .ZN(N298) );
  NAND3_X1 U1076 ( .A1(WE), .A2(n37797), .A3(n37796), .ZN(n37804) );
  OAI21_X1 U1077 ( .B1(n37798), .B2(n37804), .A(RESET), .ZN(N299) );
  OAI21_X1 U1078 ( .B1(n37799), .B2(n37804), .A(RESET), .ZN(N300) );
  OAI21_X1 U1079 ( .B1(n37800), .B2(n37804), .A(RESET), .ZN(N301) );
  OAI21_X1 U1080 ( .B1(n37801), .B2(n37804), .A(RESET), .ZN(N302) );
  OAI21_X1 U1081 ( .B1(n37802), .B2(n37804), .A(RESET), .ZN(N303) );
  OAI21_X1 U1082 ( .B1(n37803), .B2(n37804), .A(RESET), .ZN(N304) );
  OAI21_X1 U1083 ( .B1(n37805), .B2(n37804), .A(RESET), .ZN(N305) );
  INV_X1 U1084 ( .A(ADD_RDA[4]), .ZN(n37806) );
  NAND3_X1 U1085 ( .A1(ADD_RDA[3]), .A2(ADD_RDA[0]), .A3(n37806), .ZN(n37809)
         );
  NAND3_X1 U1086 ( .A1(RESET), .A2(ADD_RDA[1]), .A3(n37812), .ZN(n37824) );
  NOR2_X1 U1087 ( .A1(n37809), .A2(n37824), .ZN(n38206) );
  INV_X1 U1088 ( .A(ADD_RDA[0]), .ZN(n37807) );
  NAND3_X1 U1089 ( .A1(ADD_RDA[4]), .A2(n37817), .A3(n37807), .ZN(n37808) );
  NAND3_X1 U1090 ( .A1(RESET), .A2(n37812), .A3(n37811), .ZN(n37820) );
  NOR2_X1 U1091 ( .A1(n37808), .A2(n37820), .ZN(n38205) );
  NAND3_X1 U1092 ( .A1(ADD_RDA[0]), .A2(n37817), .A3(n37806), .ZN(n37816) );
  NOR2_X1 U1093 ( .A1(n37820), .A2(n37816), .ZN(n38208) );
  NAND3_X1 U1094 ( .A1(ADD_RDA[4]), .A2(ADD_RDA[3]), .A3(n37807), .ZN(n37815)
         );
  NOR2_X1 U1095 ( .A1(n37820), .A2(n37815), .ZN(n38207) );
  NAND3_X1 U1096 ( .A1(ADD_RDA[2]), .A2(RESET), .A3(n37811), .ZN(n37818) );
  NOR2_X1 U1097 ( .A1(ADD_RDA[4]), .A2(ADD_RDA[0]), .ZN(n37810) );
  NAND2_X1 U1098 ( .A1(ADD_RDA[3]), .A2(n37810), .ZN(n37822) );
  NOR2_X1 U1099 ( .A1(n37818), .A2(n37822), .ZN(n38210) );
  NAND3_X1 U1100 ( .A1(RESET), .A2(ADD_RDA[2]), .A3(ADD_RDA[1]), .ZN(n37821)
         );
  NOR2_X1 U1101 ( .A1(n37809), .A2(n37821), .ZN(n38209) );
  NOR2_X1 U1102 ( .A1(n37818), .A2(n37808), .ZN(n38217) );
  NOR2_X1 U1103 ( .A1(n37808), .A2(n37821), .ZN(n38216) );
  NOR2_X1 U1104 ( .A1(n37824), .A2(n37808), .ZN(n38219) );
  NOR2_X1 U1105 ( .A1(n37809), .A2(n37820), .ZN(n38218) );
  NAND3_X1 U1106 ( .A1(RESET), .A2(n37810), .A3(n37817), .ZN(n37813) );
  NAND3_X1 U1107 ( .A1(ADD_RDA[3]), .A2(ADD_RDA[4]), .A3(ADD_RDA[0]), .ZN(
        n37819) );
  NOR2_X1 U1108 ( .A1(n37821), .A2(n37819), .ZN(n38220) );
  NOR2_X1 U1109 ( .A1(n37824), .A2(n37816), .ZN(n38223) );
  NOR2_X1 U1110 ( .A1(n37820), .A2(n37822), .ZN(n38222) );
  NOR2_X1 U1111 ( .A1(n37815), .A2(n37821), .ZN(n38229) );
  NOR2_X1 U1112 ( .A1(n37818), .A2(n37819), .ZN(n38228) );
  NOR2_X1 U1113 ( .A1(n37824), .A2(n37819), .ZN(n38231) );
  NOR3_X1 U1114 ( .A1(ADD_RDA[1]), .A2(n37812), .A3(n37813), .ZN(n38230) );
  NOR2_X1 U1115 ( .A1(n37824), .A2(n37822), .ZN(n38233) );
  NOR2_X1 U1116 ( .A1(n37818), .A2(n37815), .ZN(n38232) );
  NAND2_X1 U1117 ( .A1(ADD_RDA[2]), .A2(ADD_RDA[1]), .ZN(n37814) );
  NOR2_X1 U1118 ( .A1(n37814), .A2(n37813), .ZN(n38235) );
  NOR2_X1 U1119 ( .A1(n37816), .A2(n37821), .ZN(n38234) );
  NOR2_X1 U1120 ( .A1(n37824), .A2(n37815), .ZN(n38241) );
  NOR2_X1 U1121 ( .A1(n37818), .A2(n37816), .ZN(n38240) );
  NAND3_X1 U1122 ( .A1(ADD_RDA[4]), .A2(ADD_RDA[0]), .A3(n37817), .ZN(n37823)
         );
  NOR2_X1 U1123 ( .A1(n37818), .A2(n37823), .ZN(n38243) );
  NOR2_X1 U1124 ( .A1(n37820), .A2(n37819), .ZN(n38242) );
  NOR2_X1 U1125 ( .A1(n37821), .A2(n37823), .ZN(n38245) );
  NOR2_X1 U1126 ( .A1(n37820), .A2(n37823), .ZN(n38244) );
  NOR2_X1 U1127 ( .A1(n37822), .A2(n37821), .ZN(n38247) );
  NOR2_X1 U1128 ( .A1(n37824), .A2(n37823), .ZN(n38246) );
  AOI22_X1 U1129 ( .A1(n37727), .A2(\REGISTERS[11][18] ), .B1(n37726), .B2(
        \REGISTERS[16][18] ), .ZN(n37828) );
  AOI22_X1 U1130 ( .A1(n37729), .A2(\REGISTERS[1][18] ), .B1(n37728), .B2(
        \REGISTERS[24][18] ), .ZN(n37827) );
  AOI22_X1 U1131 ( .A1(n37731), .A2(\REGISTERS[12][18] ), .B1(n37730), .B2(
        \REGISTERS[15][18] ), .ZN(n37826) );
  NAND2_X1 U1132 ( .A1(n37732), .A2(\REGISTERS[13][18] ), .ZN(n37825) );
  NAND4_X1 U1133 ( .A1(n37828), .A2(n37827), .A3(n37826), .A4(n37825), .ZN(
        n37844) );
  AOI22_X1 U1134 ( .A1(n37734), .A2(\REGISTERS[20][18] ), .B1(n37733), .B2(
        \REGISTERS[22][18] ), .ZN(n37832) );
  AOI22_X1 U1135 ( .A1(n37736), .A2(\REGISTERS[18][18] ), .B1(n37735), .B2(
        \REGISTERS[9][18] ), .ZN(n37831) );
  AOI22_X1 U1136 ( .A1(n37738), .A2(\REGISTERS[2][18] ), .B1(n37737), .B2(
        \REGISTERS[31][18] ), .ZN(n37830) );
  AOI22_X1 U1137 ( .A1(n37740), .A2(\REGISTERS[3][18] ), .B1(n37739), .B2(
        \REGISTERS[8][18] ), .ZN(n37829) );
  NAND4_X1 U1138 ( .A1(n37832), .A2(n37831), .A3(n37830), .A4(n37829), .ZN(
        n37843) );
  AOI22_X1 U1139 ( .A1(n37742), .A2(\REGISTERS[30][18] ), .B1(n37741), .B2(
        \REGISTERS[29][18] ), .ZN(n37836) );
  AOI22_X1 U1140 ( .A1(n37744), .A2(\REGISTERS[27][18] ), .B1(n37743), .B2(
        \REGISTERS[4][18] ), .ZN(n37835) );
  AOI22_X1 U1141 ( .A1(n37746), .A2(\REGISTERS[10][18] ), .B1(n37745), .B2(
        \REGISTERS[28][18] ), .ZN(n37834) );
  AOI22_X1 U1142 ( .A1(n37748), .A2(\REGISTERS[6][18] ), .B1(n37747), .B2(
        \REGISTERS[7][18] ), .ZN(n37833) );
  NAND4_X1 U1143 ( .A1(n37836), .A2(n37835), .A3(n37834), .A4(n37833), .ZN(
        n37842) );
  AOI22_X1 U1144 ( .A1(n37750), .A2(\REGISTERS[26][18] ), .B1(n37749), .B2(
        \REGISTERS[5][18] ), .ZN(n37840) );
  AOI22_X1 U1145 ( .A1(n37752), .A2(\REGISTERS[21][18] ), .B1(n37751), .B2(
        \REGISTERS[25][18] ), .ZN(n37839) );
  AOI22_X1 U1146 ( .A1(n37754), .A2(\REGISTERS[23][18] ), .B1(n37753), .B2(
        \REGISTERS[17][18] ), .ZN(n37838) );
  AOI22_X1 U1147 ( .A1(n37756), .A2(\REGISTERS[14][18] ), .B1(n37755), .B2(
        \REGISTERS[19][18] ), .ZN(n37837) );
  NAND4_X1 U1148 ( .A1(n37840), .A2(n37839), .A3(n37838), .A4(n37837), .ZN(
        n37841) );
  AOI22_X1 U1149 ( .A1(n37727), .A2(\REGISTERS[11][19] ), .B1(n37726), .B2(
        \REGISTERS[16][19] ), .ZN(n37848) );
  AOI22_X1 U1150 ( .A1(n37729), .A2(\REGISTERS[1][19] ), .B1(n37728), .B2(
        \REGISTERS[24][19] ), .ZN(n37847) );
  AOI22_X1 U1151 ( .A1(n37731), .A2(\REGISTERS[12][19] ), .B1(n37730), .B2(
        \REGISTERS[15][19] ), .ZN(n37846) );
  NAND2_X1 U1152 ( .A1(n37732), .A2(\REGISTERS[13][19] ), .ZN(n37845) );
  NAND4_X1 U1153 ( .A1(n37848), .A2(n37847), .A3(n37846), .A4(n37845), .ZN(
        n37864) );
  AOI22_X1 U1154 ( .A1(n37734), .A2(\REGISTERS[20][19] ), .B1(n37733), .B2(
        \REGISTERS[22][19] ), .ZN(n37852) );
  AOI22_X1 U1155 ( .A1(n37736), .A2(\REGISTERS[18][19] ), .B1(n37735), .B2(
        \REGISTERS[9][19] ), .ZN(n37851) );
  AOI22_X1 U1156 ( .A1(n37738), .A2(\REGISTERS[2][19] ), .B1(n37737), .B2(
        \REGISTERS[31][19] ), .ZN(n37850) );
  AOI22_X1 U1157 ( .A1(n37740), .A2(\REGISTERS[3][19] ), .B1(n37739), .B2(
        \REGISTERS[8][19] ), .ZN(n37849) );
  NAND4_X1 U1158 ( .A1(n37852), .A2(n37851), .A3(n37850), .A4(n37849), .ZN(
        n37863) );
  AOI22_X1 U1159 ( .A1(n37742), .A2(\REGISTERS[30][19] ), .B1(n37741), .B2(
        \REGISTERS[29][19] ), .ZN(n37856) );
  AOI22_X1 U1160 ( .A1(n37744), .A2(\REGISTERS[27][19] ), .B1(n37743), .B2(
        \REGISTERS[4][19] ), .ZN(n37855) );
  AOI22_X1 U1161 ( .A1(n37746), .A2(\REGISTERS[10][19] ), .B1(n37745), .B2(
        \REGISTERS[28][19] ), .ZN(n37854) );
  AOI22_X1 U1162 ( .A1(n37748), .A2(\REGISTERS[6][19] ), .B1(n37747), .B2(
        \REGISTERS[7][19] ), .ZN(n37853) );
  NAND4_X1 U1163 ( .A1(n37856), .A2(n37855), .A3(n37854), .A4(n37853), .ZN(
        n37862) );
  AOI22_X1 U1164 ( .A1(n37750), .A2(\REGISTERS[26][19] ), .B1(n37749), .B2(
        \REGISTERS[5][19] ), .ZN(n37860) );
  AOI22_X1 U1165 ( .A1(n37752), .A2(\REGISTERS[21][19] ), .B1(n37751), .B2(
        \REGISTERS[25][19] ), .ZN(n37859) );
  AOI22_X1 U1166 ( .A1(n37754), .A2(\REGISTERS[23][19] ), .B1(n37753), .B2(
        \REGISTERS[17][19] ), .ZN(n37858) );
  AOI22_X1 U1167 ( .A1(n37756), .A2(\REGISTERS[14][19] ), .B1(n37755), .B2(
        \REGISTERS[19][19] ), .ZN(n37857) );
  NAND4_X1 U1168 ( .A1(n37860), .A2(n37859), .A3(n37858), .A4(n37857), .ZN(
        n37861) );
  AOI22_X1 U1169 ( .A1(n37727), .A2(\REGISTERS[11][20] ), .B1(n37726), .B2(
        \REGISTERS[16][20] ), .ZN(n37868) );
  AOI22_X1 U1170 ( .A1(n37729), .A2(\REGISTERS[1][20] ), .B1(n37728), .B2(
        \REGISTERS[24][20] ), .ZN(n37867) );
  AOI22_X1 U1171 ( .A1(n37731), .A2(\REGISTERS[12][20] ), .B1(n37730), .B2(
        \REGISTERS[15][20] ), .ZN(n37866) );
  NAND2_X1 U1172 ( .A1(n37732), .A2(\REGISTERS[13][20] ), .ZN(n37865) );
  NAND4_X1 U1173 ( .A1(n37868), .A2(n37867), .A3(n37866), .A4(n37865), .ZN(
        n37884) );
  AOI22_X1 U1174 ( .A1(n37734), .A2(\REGISTERS[20][20] ), .B1(n37733), .B2(
        \REGISTERS[22][20] ), .ZN(n37872) );
  AOI22_X1 U1175 ( .A1(n37736), .A2(\REGISTERS[18][20] ), .B1(n37735), .B2(
        \REGISTERS[9][20] ), .ZN(n37871) );
  AOI22_X1 U1176 ( .A1(n38221), .A2(\REGISTERS[2][20] ), .B1(n37737), .B2(
        \REGISTERS[31][20] ), .ZN(n37870) );
  AOI22_X1 U1177 ( .A1(n37740), .A2(\REGISTERS[3][20] ), .B1(n37739), .B2(
        \REGISTERS[8][20] ), .ZN(n37869) );
  NAND4_X1 U1178 ( .A1(n37872), .A2(n37871), .A3(n37870), .A4(n37869), .ZN(
        n37883) );
  AOI22_X1 U1179 ( .A1(n37742), .A2(\REGISTERS[30][20] ), .B1(n37741), .B2(
        \REGISTERS[29][20] ), .ZN(n37876) );
  AOI22_X1 U1180 ( .A1(n37744), .A2(\REGISTERS[27][20] ), .B1(n37743), .B2(
        \REGISTERS[4][20] ), .ZN(n37875) );
  AOI22_X1 U1181 ( .A1(n37746), .A2(\REGISTERS[10][20] ), .B1(n37745), .B2(
        \REGISTERS[28][20] ), .ZN(n37874) );
  AOI22_X1 U1182 ( .A1(n37748), .A2(\REGISTERS[6][20] ), .B1(n37747), .B2(
        \REGISTERS[7][20] ), .ZN(n37873) );
  NAND4_X1 U1183 ( .A1(n37876), .A2(n37875), .A3(n37874), .A4(n37873), .ZN(
        n37882) );
  AOI22_X1 U1184 ( .A1(n37750), .A2(\REGISTERS[26][20] ), .B1(n37749), .B2(
        \REGISTERS[5][20] ), .ZN(n37880) );
  AOI22_X1 U1185 ( .A1(n37752), .A2(\REGISTERS[21][20] ), .B1(n37751), .B2(
        \REGISTERS[25][20] ), .ZN(n37879) );
  AOI22_X1 U1186 ( .A1(n37754), .A2(\REGISTERS[23][20] ), .B1(n37753), .B2(
        \REGISTERS[17][20] ), .ZN(n37878) );
  AOI22_X1 U1187 ( .A1(n37756), .A2(\REGISTERS[14][20] ), .B1(n37755), .B2(
        \REGISTERS[19][20] ), .ZN(n37877) );
  NAND4_X1 U1188 ( .A1(n37880), .A2(n37879), .A3(n37878), .A4(n37877), .ZN(
        n37881) );
  AOI22_X1 U1189 ( .A1(n37727), .A2(\REGISTERS[11][21] ), .B1(n37726), .B2(
        \REGISTERS[16][21] ), .ZN(n37888) );
  AOI22_X1 U1190 ( .A1(n37729), .A2(\REGISTERS[1][21] ), .B1(n37728), .B2(
        \REGISTERS[24][21] ), .ZN(n37887) );
  AOI22_X1 U1191 ( .A1(n37731), .A2(\REGISTERS[12][21] ), .B1(n37730), .B2(
        \REGISTERS[15][21] ), .ZN(n37886) );
  NAND2_X1 U1192 ( .A1(n37732), .A2(\REGISTERS[13][21] ), .ZN(n37885) );
  NAND4_X1 U1193 ( .A1(n37888), .A2(n37887), .A3(n37886), .A4(n37885), .ZN(
        n37904) );
  AOI22_X1 U1194 ( .A1(n37734), .A2(\REGISTERS[20][21] ), .B1(n37733), .B2(
        \REGISTERS[22][21] ), .ZN(n37892) );
  AOI22_X1 U1195 ( .A1(n37736), .A2(\REGISTERS[18][21] ), .B1(n37735), .B2(
        \REGISTERS[9][21] ), .ZN(n37891) );
  AOI22_X1 U1196 ( .A1(n37738), .A2(\REGISTERS[2][21] ), .B1(n37737), .B2(
        \REGISTERS[31][21] ), .ZN(n37890) );
  AOI22_X1 U1197 ( .A1(n37740), .A2(\REGISTERS[3][21] ), .B1(n37739), .B2(
        \REGISTERS[8][21] ), .ZN(n37889) );
  NAND4_X1 U1198 ( .A1(n37892), .A2(n37891), .A3(n37890), .A4(n37889), .ZN(
        n37903) );
  AOI22_X1 U1199 ( .A1(n37742), .A2(\REGISTERS[30][21] ), .B1(n37741), .B2(
        \REGISTERS[29][21] ), .ZN(n37896) );
  AOI22_X1 U1200 ( .A1(n37744), .A2(\REGISTERS[27][21] ), .B1(n37743), .B2(
        \REGISTERS[4][21] ), .ZN(n37895) );
  AOI22_X1 U1201 ( .A1(n37746), .A2(\REGISTERS[10][21] ), .B1(n37745), .B2(
        \REGISTERS[28][21] ), .ZN(n37894) );
  AOI22_X1 U1202 ( .A1(n37748), .A2(\REGISTERS[6][21] ), .B1(n37747), .B2(
        \REGISTERS[7][21] ), .ZN(n37893) );
  NAND4_X1 U1203 ( .A1(n37896), .A2(n37895), .A3(n37894), .A4(n37893), .ZN(
        n37902) );
  AOI22_X1 U1204 ( .A1(n37750), .A2(\REGISTERS[26][21] ), .B1(n37749), .B2(
        \REGISTERS[5][21] ), .ZN(n37900) );
  AOI22_X1 U1205 ( .A1(n37752), .A2(\REGISTERS[21][21] ), .B1(n37751), .B2(
        \REGISTERS[25][21] ), .ZN(n37899) );
  AOI22_X1 U1206 ( .A1(n37754), .A2(\REGISTERS[23][21] ), .B1(n37753), .B2(
        \REGISTERS[17][21] ), .ZN(n37898) );
  AOI22_X1 U1207 ( .A1(n37756), .A2(\REGISTERS[14][21] ), .B1(n37755), .B2(
        \REGISTERS[19][21] ), .ZN(n37897) );
  NAND4_X1 U1208 ( .A1(n37900), .A2(n37899), .A3(n37898), .A4(n37897), .ZN(
        n37901) );
  AOI22_X1 U1209 ( .A1(n37727), .A2(\REGISTERS[11][22] ), .B1(n37726), .B2(
        \REGISTERS[16][22] ), .ZN(n37908) );
  AOI22_X1 U1210 ( .A1(n37729), .A2(\REGISTERS[1][22] ), .B1(n37728), .B2(
        \REGISTERS[24][22] ), .ZN(n37907) );
  AOI22_X1 U1211 ( .A1(n37731), .A2(\REGISTERS[12][22] ), .B1(n37730), .B2(
        \REGISTERS[15][22] ), .ZN(n37906) );
  NAND2_X1 U1212 ( .A1(n37732), .A2(\REGISTERS[13][22] ), .ZN(n37905) );
  NAND4_X1 U1213 ( .A1(n37908), .A2(n37907), .A3(n37906), .A4(n37905), .ZN(
        n37924) );
  AOI22_X1 U1214 ( .A1(n37734), .A2(\REGISTERS[20][22] ), .B1(n37733), .B2(
        \REGISTERS[22][22] ), .ZN(n37912) );
  AOI22_X1 U1215 ( .A1(n37736), .A2(\REGISTERS[18][22] ), .B1(n37735), .B2(
        \REGISTERS[9][22] ), .ZN(n37911) );
  AOI22_X1 U1216 ( .A1(n37738), .A2(\REGISTERS[2][22] ), .B1(n37737), .B2(
        \REGISTERS[31][22] ), .ZN(n37910) );
  AOI22_X1 U1217 ( .A1(n37740), .A2(\REGISTERS[3][22] ), .B1(n37739), .B2(
        \REGISTERS[8][22] ), .ZN(n37909) );
  NAND4_X1 U1218 ( .A1(n37912), .A2(n37911), .A3(n37910), .A4(n37909), .ZN(
        n37923) );
  AOI22_X1 U1219 ( .A1(n37742), .A2(\REGISTERS[30][22] ), .B1(n37741), .B2(
        \REGISTERS[29][22] ), .ZN(n37916) );
  AOI22_X1 U1220 ( .A1(n37744), .A2(\REGISTERS[27][22] ), .B1(n37743), .B2(
        \REGISTERS[4][22] ), .ZN(n37915) );
  AOI22_X1 U1221 ( .A1(n37746), .A2(\REGISTERS[10][22] ), .B1(n37745), .B2(
        \REGISTERS[28][22] ), .ZN(n37914) );
  AOI22_X1 U1222 ( .A1(n37748), .A2(\REGISTERS[6][22] ), .B1(n37747), .B2(
        \REGISTERS[7][22] ), .ZN(n37913) );
  NAND4_X1 U1223 ( .A1(n37916), .A2(n37915), .A3(n37914), .A4(n37913), .ZN(
        n37922) );
  AOI22_X1 U1224 ( .A1(n37750), .A2(\REGISTERS[26][22] ), .B1(n37749), .B2(
        \REGISTERS[5][22] ), .ZN(n37920) );
  AOI22_X1 U1225 ( .A1(n37752), .A2(\REGISTERS[21][22] ), .B1(n37751), .B2(
        \REGISTERS[25][22] ), .ZN(n37919) );
  AOI22_X1 U1226 ( .A1(n37754), .A2(\REGISTERS[23][22] ), .B1(n37753), .B2(
        \REGISTERS[17][22] ), .ZN(n37918) );
  AOI22_X1 U1227 ( .A1(n37756), .A2(\REGISTERS[14][22] ), .B1(n37755), .B2(
        \REGISTERS[19][22] ), .ZN(n37917) );
  NAND4_X1 U1228 ( .A1(n37920), .A2(n37919), .A3(n37918), .A4(n37917), .ZN(
        n37921) );
  AOI22_X1 U1229 ( .A1(n37727), .A2(\REGISTERS[11][23] ), .B1(n37726), .B2(
        \REGISTERS[16][23] ), .ZN(n37928) );
  AOI22_X1 U1230 ( .A1(n37729), .A2(\REGISTERS[1][23] ), .B1(n37728), .B2(
        \REGISTERS[24][23] ), .ZN(n37927) );
  AOI22_X1 U1231 ( .A1(n37731), .A2(\REGISTERS[12][23] ), .B1(n37730), .B2(
        \REGISTERS[15][23] ), .ZN(n37926) );
  NAND2_X1 U1232 ( .A1(n37732), .A2(\REGISTERS[13][23] ), .ZN(n37925) );
  NAND4_X1 U1233 ( .A1(n37928), .A2(n37927), .A3(n37926), .A4(n37925), .ZN(
        n37944) );
  AOI22_X1 U1234 ( .A1(n37734), .A2(\REGISTERS[20][23] ), .B1(n37733), .B2(
        \REGISTERS[22][23] ), .ZN(n37932) );
  AOI22_X1 U1235 ( .A1(n37736), .A2(\REGISTERS[18][23] ), .B1(n37735), .B2(
        \REGISTERS[9][23] ), .ZN(n37931) );
  AOI22_X1 U1236 ( .A1(n37738), .A2(\REGISTERS[2][23] ), .B1(n37737), .B2(
        \REGISTERS[31][23] ), .ZN(n37930) );
  AOI22_X1 U1237 ( .A1(n37740), .A2(\REGISTERS[3][23] ), .B1(n37739), .B2(
        \REGISTERS[8][23] ), .ZN(n37929) );
  NAND4_X1 U1238 ( .A1(n37932), .A2(n37931), .A3(n37930), .A4(n37929), .ZN(
        n37943) );
  AOI22_X1 U1239 ( .A1(n37742), .A2(\REGISTERS[30][23] ), .B1(n37741), .B2(
        \REGISTERS[29][23] ), .ZN(n37936) );
  AOI22_X1 U1240 ( .A1(n37744), .A2(\REGISTERS[27][23] ), .B1(n37743), .B2(
        \REGISTERS[4][23] ), .ZN(n37935) );
  AOI22_X1 U1241 ( .A1(n37746), .A2(\REGISTERS[10][23] ), .B1(n37745), .B2(
        \REGISTERS[28][23] ), .ZN(n37934) );
  AOI22_X1 U1242 ( .A1(n37748), .A2(\REGISTERS[6][23] ), .B1(n37747), .B2(
        \REGISTERS[7][23] ), .ZN(n37933) );
  NAND4_X1 U1243 ( .A1(n37936), .A2(n37935), .A3(n37934), .A4(n37933), .ZN(
        n37942) );
  AOI22_X1 U1244 ( .A1(n37750), .A2(\REGISTERS[26][23] ), .B1(n37749), .B2(
        \REGISTERS[5][23] ), .ZN(n37940) );
  AOI22_X1 U1245 ( .A1(n37752), .A2(\REGISTERS[21][23] ), .B1(n37751), .B2(
        \REGISTERS[25][23] ), .ZN(n37939) );
  AOI22_X1 U1246 ( .A1(n37754), .A2(\REGISTERS[23][23] ), .B1(n37753), .B2(
        \REGISTERS[17][23] ), .ZN(n37938) );
  AOI22_X1 U1247 ( .A1(n37756), .A2(\REGISTERS[14][23] ), .B1(n37755), .B2(
        \REGISTERS[19][23] ), .ZN(n37937) );
  NAND4_X1 U1248 ( .A1(n37940), .A2(n37939), .A3(n37938), .A4(n37937), .ZN(
        n37941) );
  AOI22_X1 U1249 ( .A1(n37727), .A2(\REGISTERS[11][24] ), .B1(n37726), .B2(
        \REGISTERS[16][24] ), .ZN(n37948) );
  AOI22_X1 U1250 ( .A1(n37729), .A2(\REGISTERS[1][24] ), .B1(n37728), .B2(
        \REGISTERS[24][24] ), .ZN(n37947) );
  AOI22_X1 U1251 ( .A1(n37731), .A2(\REGISTERS[12][24] ), .B1(n37730), .B2(
        \REGISTERS[15][24] ), .ZN(n37946) );
  NAND2_X1 U1252 ( .A1(n37732), .A2(\REGISTERS[13][24] ), .ZN(n37945) );
  NAND4_X1 U1253 ( .A1(n37948), .A2(n37947), .A3(n37946), .A4(n37945), .ZN(
        n37964) );
  AOI22_X1 U1254 ( .A1(n37734), .A2(\REGISTERS[20][24] ), .B1(n37733), .B2(
        \REGISTERS[22][24] ), .ZN(n37952) );
  AOI22_X1 U1255 ( .A1(n37736), .A2(\REGISTERS[18][24] ), .B1(n37735), .B2(
        \REGISTERS[9][24] ), .ZN(n37951) );
  AOI22_X1 U1256 ( .A1(n37738), .A2(\REGISTERS[2][24] ), .B1(n37737), .B2(
        \REGISTERS[31][24] ), .ZN(n37950) );
  AOI22_X1 U1257 ( .A1(n37740), .A2(\REGISTERS[3][24] ), .B1(n37739), .B2(
        \REGISTERS[8][24] ), .ZN(n37949) );
  NAND4_X1 U1258 ( .A1(n37952), .A2(n37951), .A3(n37950), .A4(n37949), .ZN(
        n37963) );
  AOI22_X1 U1259 ( .A1(n37742), .A2(\REGISTERS[30][24] ), .B1(n37741), .B2(
        \REGISTERS[29][24] ), .ZN(n37956) );
  AOI22_X1 U1260 ( .A1(n37744), .A2(\REGISTERS[27][24] ), .B1(n37743), .B2(
        \REGISTERS[4][24] ), .ZN(n37955) );
  AOI22_X1 U1261 ( .A1(n37746), .A2(\REGISTERS[10][24] ), .B1(n37745), .B2(
        \REGISTERS[28][24] ), .ZN(n37954) );
  AOI22_X1 U1262 ( .A1(n37748), .A2(\REGISTERS[6][24] ), .B1(n37747), .B2(
        \REGISTERS[7][24] ), .ZN(n37953) );
  NAND4_X1 U1263 ( .A1(n37956), .A2(n37955), .A3(n37954), .A4(n37953), .ZN(
        n37962) );
  AOI22_X1 U1264 ( .A1(n37750), .A2(\REGISTERS[26][24] ), .B1(n37749), .B2(
        \REGISTERS[5][24] ), .ZN(n37960) );
  AOI22_X1 U1265 ( .A1(n37752), .A2(\REGISTERS[21][24] ), .B1(n37751), .B2(
        \REGISTERS[25][24] ), .ZN(n37959) );
  AOI22_X1 U1266 ( .A1(n37754), .A2(\REGISTERS[23][24] ), .B1(n37753), .B2(
        \REGISTERS[17][24] ), .ZN(n37958) );
  AOI22_X1 U1267 ( .A1(n37756), .A2(\REGISTERS[14][24] ), .B1(n37755), .B2(
        \REGISTERS[19][24] ), .ZN(n37957) );
  NAND4_X1 U1268 ( .A1(n37960), .A2(n37959), .A3(n37958), .A4(n37957), .ZN(
        n37961) );
  AOI22_X1 U1269 ( .A1(n37727), .A2(\REGISTERS[11][25] ), .B1(n37726), .B2(
        \REGISTERS[16][25] ), .ZN(n37968) );
  AOI22_X1 U1270 ( .A1(n37729), .A2(\REGISTERS[1][25] ), .B1(n37728), .B2(
        \REGISTERS[24][25] ), .ZN(n37967) );
  AOI22_X1 U1271 ( .A1(n37731), .A2(\REGISTERS[12][25] ), .B1(n37730), .B2(
        \REGISTERS[15][25] ), .ZN(n37966) );
  NAND2_X1 U1272 ( .A1(n37732), .A2(\REGISTERS[13][25] ), .ZN(n37965) );
  NAND4_X1 U1273 ( .A1(n37968), .A2(n37967), .A3(n37966), .A4(n37965), .ZN(
        n37984) );
  AOI22_X1 U1274 ( .A1(n37734), .A2(\REGISTERS[20][25] ), .B1(n37733), .B2(
        \REGISTERS[22][25] ), .ZN(n37972) );
  AOI22_X1 U1275 ( .A1(n37736), .A2(\REGISTERS[18][25] ), .B1(n37735), .B2(
        \REGISTERS[9][25] ), .ZN(n37971) );
  AOI22_X1 U1276 ( .A1(n37738), .A2(\REGISTERS[2][25] ), .B1(n37737), .B2(
        \REGISTERS[31][25] ), .ZN(n37970) );
  AOI22_X1 U1277 ( .A1(n37740), .A2(\REGISTERS[3][25] ), .B1(n37739), .B2(
        \REGISTERS[8][25] ), .ZN(n37969) );
  NAND4_X1 U1278 ( .A1(n37972), .A2(n37971), .A3(n37970), .A4(n37969), .ZN(
        n37983) );
  AOI22_X1 U1279 ( .A1(n37742), .A2(\REGISTERS[30][25] ), .B1(n37741), .B2(
        \REGISTERS[29][25] ), .ZN(n37976) );
  AOI22_X1 U1280 ( .A1(n37744), .A2(\REGISTERS[27][25] ), .B1(n37743), .B2(
        \REGISTERS[4][25] ), .ZN(n37975) );
  AOI22_X1 U1281 ( .A1(n37746), .A2(\REGISTERS[10][25] ), .B1(n37745), .B2(
        \REGISTERS[28][25] ), .ZN(n37974) );
  AOI22_X1 U1282 ( .A1(n37748), .A2(\REGISTERS[6][25] ), .B1(n37747), .B2(
        \REGISTERS[7][25] ), .ZN(n37973) );
  NAND4_X1 U1283 ( .A1(n37976), .A2(n37975), .A3(n37974), .A4(n37973), .ZN(
        n37982) );
  AOI22_X1 U1284 ( .A1(n37750), .A2(\REGISTERS[26][25] ), .B1(n37749), .B2(
        \REGISTERS[5][25] ), .ZN(n37980) );
  AOI22_X1 U1285 ( .A1(n37752), .A2(\REGISTERS[21][25] ), .B1(n37751), .B2(
        \REGISTERS[25][25] ), .ZN(n37979) );
  AOI22_X1 U1286 ( .A1(n37754), .A2(\REGISTERS[23][25] ), .B1(n37753), .B2(
        \REGISTERS[17][25] ), .ZN(n37978) );
  AOI22_X1 U1287 ( .A1(n37756), .A2(\REGISTERS[14][25] ), .B1(n37755), .B2(
        \REGISTERS[19][25] ), .ZN(n37977) );
  NAND4_X1 U1288 ( .A1(n37980), .A2(n37979), .A3(n37978), .A4(n37977), .ZN(
        n37981) );
  AOI22_X1 U1289 ( .A1(n37727), .A2(\REGISTERS[11][26] ), .B1(n38205), .B2(
        \REGISTERS[16][26] ), .ZN(n37988) );
  AOI22_X1 U1290 ( .A1(n37729), .A2(\REGISTERS[1][26] ), .B1(n38207), .B2(
        \REGISTERS[24][26] ), .ZN(n37987) );
  AOI22_X1 U1291 ( .A1(n37731), .A2(\REGISTERS[12][26] ), .B1(n38209), .B2(
        \REGISTERS[15][26] ), .ZN(n37986) );
  NAND2_X1 U1292 ( .A1(n37732), .A2(\REGISTERS[13][26] ), .ZN(n37985) );
  NAND4_X1 U1293 ( .A1(n37988), .A2(n37987), .A3(n37986), .A4(n37985), .ZN(
        n38004) );
  AOI22_X1 U1294 ( .A1(n37734), .A2(\REGISTERS[20][26] ), .B1(n38216), .B2(
        \REGISTERS[22][26] ), .ZN(n37992) );
  AOI22_X1 U1295 ( .A1(n37736), .A2(\REGISTERS[18][26] ), .B1(n38218), .B2(
        \REGISTERS[9][26] ), .ZN(n37991) );
  AOI22_X1 U1296 ( .A1(n37738), .A2(\REGISTERS[2][26] ), .B1(n38220), .B2(
        \REGISTERS[31][26] ), .ZN(n37990) );
  AOI22_X1 U1297 ( .A1(n37740), .A2(\REGISTERS[3][26] ), .B1(n38222), .B2(
        \REGISTERS[8][26] ), .ZN(n37989) );
  NAND4_X1 U1298 ( .A1(n37992), .A2(n37991), .A3(n37990), .A4(n37989), .ZN(
        n38003) );
  AOI22_X1 U1299 ( .A1(n37742), .A2(\REGISTERS[30][26] ), .B1(n38228), .B2(
        \REGISTERS[29][26] ), .ZN(n37996) );
  AOI22_X1 U1300 ( .A1(n38231), .A2(\REGISTERS[27][26] ), .B1(n37743), .B2(
        \REGISTERS[4][26] ), .ZN(n37995) );
  AOI22_X1 U1301 ( .A1(n37746), .A2(\REGISTERS[10][26] ), .B1(n38232), .B2(
        \REGISTERS[28][26] ), .ZN(n37994) );
  AOI22_X1 U1302 ( .A1(n37748), .A2(\REGISTERS[6][26] ), .B1(n38234), .B2(
        \REGISTERS[7][26] ), .ZN(n37993) );
  NAND4_X1 U1303 ( .A1(n37996), .A2(n37995), .A3(n37994), .A4(n37993), .ZN(
        n38002) );
  AOI22_X1 U1304 ( .A1(n37750), .A2(\REGISTERS[26][26] ), .B1(n38240), .B2(
        \REGISTERS[5][26] ), .ZN(n38000) );
  AOI22_X1 U1305 ( .A1(n37752), .A2(\REGISTERS[21][26] ), .B1(n37751), .B2(
        \REGISTERS[25][26] ), .ZN(n37999) );
  AOI22_X1 U1306 ( .A1(n37754), .A2(\REGISTERS[23][26] ), .B1(n37753), .B2(
        \REGISTERS[17][26] ), .ZN(n37998) );
  AOI22_X1 U1307 ( .A1(n37756), .A2(\REGISTERS[14][26] ), .B1(n37755), .B2(
        \REGISTERS[19][26] ), .ZN(n37997) );
  NAND4_X1 U1308 ( .A1(n38000), .A2(n37999), .A3(n37998), .A4(n37997), .ZN(
        n38001) );
  AOI22_X1 U1309 ( .A1(n38206), .A2(\REGISTERS[11][27] ), .B1(n38205), .B2(
        \REGISTERS[16][27] ), .ZN(n38008) );
  AOI22_X1 U1310 ( .A1(n38208), .A2(\REGISTERS[1][27] ), .B1(n38207), .B2(
        \REGISTERS[24][27] ), .ZN(n38007) );
  AOI22_X1 U1311 ( .A1(n38210), .A2(\REGISTERS[12][27] ), .B1(n38209), .B2(
        \REGISTERS[15][27] ), .ZN(n38006) );
  NAND2_X1 U1312 ( .A1(n38211), .A2(\REGISTERS[13][27] ), .ZN(n38005) );
  NAND4_X1 U1313 ( .A1(n38008), .A2(n38007), .A3(n38006), .A4(n38005), .ZN(
        n38024) );
  AOI22_X1 U1314 ( .A1(n38217), .A2(\REGISTERS[20][27] ), .B1(n38216), .B2(
        \REGISTERS[22][27] ), .ZN(n38012) );
  AOI22_X1 U1315 ( .A1(n38219), .A2(\REGISTERS[18][27] ), .B1(n37735), .B2(
        \REGISTERS[9][27] ), .ZN(n38011) );
  AOI22_X1 U1316 ( .A1(n37738), .A2(\REGISTERS[2][27] ), .B1(n38220), .B2(
        \REGISTERS[31][27] ), .ZN(n38010) );
  AOI22_X1 U1317 ( .A1(n38223), .A2(\REGISTERS[3][27] ), .B1(n37739), .B2(
        \REGISTERS[8][27] ), .ZN(n38009) );
  NAND4_X1 U1318 ( .A1(n38012), .A2(n38011), .A3(n38010), .A4(n38009), .ZN(
        n38023) );
  AOI22_X1 U1319 ( .A1(n38229), .A2(\REGISTERS[30][27] ), .B1(n38228), .B2(
        \REGISTERS[29][27] ), .ZN(n38016) );
  AOI22_X1 U1320 ( .A1(n37744), .A2(\REGISTERS[27][27] ), .B1(n37743), .B2(
        \REGISTERS[4][27] ), .ZN(n38015) );
  AOI22_X1 U1321 ( .A1(n38233), .A2(\REGISTERS[10][27] ), .B1(n38232), .B2(
        \REGISTERS[28][27] ), .ZN(n38014) );
  AOI22_X1 U1322 ( .A1(n38235), .A2(\REGISTERS[6][27] ), .B1(n37747), .B2(
        \REGISTERS[7][27] ), .ZN(n38013) );
  NAND4_X1 U1323 ( .A1(n38016), .A2(n38015), .A3(n38014), .A4(n38013), .ZN(
        n38022) );
  AOI22_X1 U1324 ( .A1(n37750), .A2(\REGISTERS[26][27] ), .B1(n38240), .B2(
        \REGISTERS[5][27] ), .ZN(n38020) );
  AOI22_X1 U1325 ( .A1(n37752), .A2(\REGISTERS[21][27] ), .B1(n38242), .B2(
        \REGISTERS[25][27] ), .ZN(n38019) );
  AOI22_X1 U1326 ( .A1(n38245), .A2(\REGISTERS[23][27] ), .B1(n38244), .B2(
        \REGISTERS[17][27] ), .ZN(n38018) );
  AOI22_X1 U1327 ( .A1(n38247), .A2(\REGISTERS[14][27] ), .B1(n38246), .B2(
        \REGISTERS[19][27] ), .ZN(n38017) );
  NAND4_X1 U1328 ( .A1(n38020), .A2(n38019), .A3(n38018), .A4(n38017), .ZN(
        n38021) );
  AOI22_X1 U1329 ( .A1(n38206), .A2(\REGISTERS[11][28] ), .B1(n37726), .B2(
        \REGISTERS[16][28] ), .ZN(n38028) );
  AOI22_X1 U1330 ( .A1(n38208), .A2(\REGISTERS[1][28] ), .B1(n37728), .B2(
        \REGISTERS[24][28] ), .ZN(n38027) );
  AOI22_X1 U1331 ( .A1(n38210), .A2(\REGISTERS[12][28] ), .B1(n38209), .B2(
        \REGISTERS[15][28] ), .ZN(n38026) );
  NAND2_X1 U1332 ( .A1(n38211), .A2(\REGISTERS[13][28] ), .ZN(n38025) );
  NAND4_X1 U1333 ( .A1(n38028), .A2(n38027), .A3(n38026), .A4(n38025), .ZN(
        n38044) );
  AOI22_X1 U1334 ( .A1(n37734), .A2(\REGISTERS[20][28] ), .B1(n37733), .B2(
        \REGISTERS[22][28] ), .ZN(n38032) );
  AOI22_X1 U1335 ( .A1(n37736), .A2(\REGISTERS[18][28] ), .B1(n38218), .B2(
        \REGISTERS[9][28] ), .ZN(n38031) );
  AOI22_X1 U1336 ( .A1(n37738), .A2(\REGISTERS[2][28] ), .B1(n38220), .B2(
        \REGISTERS[31][28] ), .ZN(n38030) );
  AOI22_X1 U1337 ( .A1(n37740), .A2(\REGISTERS[3][28] ), .B1(n38222), .B2(
        \REGISTERS[8][28] ), .ZN(n38029) );
  NAND4_X1 U1338 ( .A1(n38032), .A2(n38031), .A3(n38030), .A4(n38029), .ZN(
        n38043) );
  AOI22_X1 U1339 ( .A1(n37742), .A2(\REGISTERS[30][28] ), .B1(n38228), .B2(
        \REGISTERS[29][28] ), .ZN(n38036) );
  AOI22_X1 U1340 ( .A1(n38231), .A2(\REGISTERS[27][28] ), .B1(n37743), .B2(
        \REGISTERS[4][28] ), .ZN(n38035) );
  AOI22_X1 U1341 ( .A1(n37746), .A2(\REGISTERS[10][28] ), .B1(n38232), .B2(
        \REGISTERS[28][28] ), .ZN(n38034) );
  AOI22_X1 U1342 ( .A1(n37748), .A2(\REGISTERS[6][28] ), .B1(n38234), .B2(
        \REGISTERS[7][28] ), .ZN(n38033) );
  NAND4_X1 U1343 ( .A1(n38036), .A2(n38035), .A3(n38034), .A4(n38033), .ZN(
        n38042) );
  AOI22_X1 U1344 ( .A1(n38241), .A2(\REGISTERS[26][28] ), .B1(n38240), .B2(
        \REGISTERS[5][28] ), .ZN(n38040) );
  AOI22_X1 U1345 ( .A1(n38243), .A2(\REGISTERS[21][28] ), .B1(n38242), .B2(
        \REGISTERS[25][28] ), .ZN(n38039) );
  AOI22_X1 U1346 ( .A1(n37754), .A2(\REGISTERS[23][28] ), .B1(n38244), .B2(
        \REGISTERS[17][28] ), .ZN(n38038) );
  AOI22_X1 U1347 ( .A1(n37756), .A2(\REGISTERS[14][28] ), .B1(n38246), .B2(
        \REGISTERS[19][28] ), .ZN(n38037) );
  NAND4_X1 U1348 ( .A1(n38040), .A2(n38039), .A3(n38038), .A4(n38037), .ZN(
        n38041) );
  AOI22_X1 U1349 ( .A1(n38206), .A2(\REGISTERS[11][29] ), .B1(n38205), .B2(
        \REGISTERS[16][29] ), .ZN(n38048) );
  AOI22_X1 U1350 ( .A1(n38208), .A2(\REGISTERS[1][29] ), .B1(n38207), .B2(
        \REGISTERS[24][29] ), .ZN(n38047) );
  AOI22_X1 U1351 ( .A1(n38210), .A2(\REGISTERS[12][29] ), .B1(n38209), .B2(
        \REGISTERS[15][29] ), .ZN(n38046) );
  NAND2_X1 U1352 ( .A1(n38211), .A2(\REGISTERS[13][29] ), .ZN(n38045) );
  NAND4_X1 U1353 ( .A1(n38048), .A2(n38047), .A3(n38046), .A4(n38045), .ZN(
        n38064) );
  AOI22_X1 U1354 ( .A1(n38217), .A2(\REGISTERS[20][29] ), .B1(n38216), .B2(
        \REGISTERS[22][29] ), .ZN(n38052) );
  AOI22_X1 U1355 ( .A1(n38219), .A2(\REGISTERS[18][29] ), .B1(n38218), .B2(
        \REGISTERS[9][29] ), .ZN(n38051) );
  AOI22_X1 U1356 ( .A1(n37738), .A2(\REGISTERS[2][29] ), .B1(n38220), .B2(
        \REGISTERS[31][29] ), .ZN(n38050) );
  AOI22_X1 U1357 ( .A1(n38223), .A2(\REGISTERS[3][29] ), .B1(n38222), .B2(
        \REGISTERS[8][29] ), .ZN(n38049) );
  NAND4_X1 U1358 ( .A1(n38052), .A2(n38051), .A3(n38050), .A4(n38049), .ZN(
        n38063) );
  AOI22_X1 U1359 ( .A1(n38229), .A2(\REGISTERS[30][29] ), .B1(n38228), .B2(
        \REGISTERS[29][29] ), .ZN(n38056) );
  AOI22_X1 U1360 ( .A1(n38231), .A2(\REGISTERS[27][29] ), .B1(n37743), .B2(
        \REGISTERS[4][29] ), .ZN(n38055) );
  AOI22_X1 U1361 ( .A1(n38233), .A2(\REGISTERS[10][29] ), .B1(n38232), .B2(
        \REGISTERS[28][29] ), .ZN(n38054) );
  AOI22_X1 U1362 ( .A1(n38235), .A2(\REGISTERS[6][29] ), .B1(n38234), .B2(
        \REGISTERS[7][29] ), .ZN(n38053) );
  NAND4_X1 U1363 ( .A1(n38056), .A2(n38055), .A3(n38054), .A4(n38053), .ZN(
        n38062) );
  AOI22_X1 U1364 ( .A1(n38241), .A2(\REGISTERS[26][29] ), .B1(n38240), .B2(
        \REGISTERS[5][29] ), .ZN(n38060) );
  AOI22_X1 U1365 ( .A1(n38243), .A2(\REGISTERS[21][29] ), .B1(n38242), .B2(
        \REGISTERS[25][29] ), .ZN(n38059) );
  AOI22_X1 U1366 ( .A1(n38245), .A2(\REGISTERS[23][29] ), .B1(n38244), .B2(
        \REGISTERS[17][29] ), .ZN(n38058) );
  AOI22_X1 U1367 ( .A1(n38247), .A2(\REGISTERS[14][29] ), .B1(n38246), .B2(
        \REGISTERS[19][29] ), .ZN(n38057) );
  NAND4_X1 U1368 ( .A1(n38060), .A2(n38059), .A3(n38058), .A4(n38057), .ZN(
        n38061) );
  AOI22_X1 U1369 ( .A1(n38206), .A2(\REGISTERS[11][2] ), .B1(n38205), .B2(
        \REGISTERS[16][2] ), .ZN(n38068) );
  AOI22_X1 U1370 ( .A1(n38208), .A2(\REGISTERS[1][2] ), .B1(n38207), .B2(
        \REGISTERS[24][2] ), .ZN(n38067) );
  AOI22_X1 U1371 ( .A1(n38210), .A2(\REGISTERS[12][2] ), .B1(n38209), .B2(
        \REGISTERS[15][2] ), .ZN(n38066) );
  NAND2_X1 U1372 ( .A1(n38211), .A2(\REGISTERS[13][2] ), .ZN(n38065) );
  NAND4_X1 U1373 ( .A1(n38068), .A2(n38067), .A3(n38066), .A4(n38065), .ZN(
        n38084) );
  AOI22_X1 U1374 ( .A1(n38217), .A2(\REGISTERS[20][2] ), .B1(n38216), .B2(
        \REGISTERS[22][2] ), .ZN(n38072) );
  AOI22_X1 U1375 ( .A1(n38219), .A2(\REGISTERS[18][2] ), .B1(n38218), .B2(
        \REGISTERS[9][2] ), .ZN(n38071) );
  AOI22_X1 U1376 ( .A1(n38221), .A2(\REGISTERS[2][2] ), .B1(n38220), .B2(
        \REGISTERS[31][2] ), .ZN(n38070) );
  AOI22_X1 U1377 ( .A1(n38223), .A2(\REGISTERS[3][2] ), .B1(n38222), .B2(
        \REGISTERS[8][2] ), .ZN(n38069) );
  NAND4_X1 U1378 ( .A1(n38072), .A2(n38071), .A3(n38070), .A4(n38069), .ZN(
        n38083) );
  AOI22_X1 U1379 ( .A1(n38229), .A2(\REGISTERS[30][2] ), .B1(n38228), .B2(
        \REGISTERS[29][2] ), .ZN(n38076) );
  AOI22_X1 U1380 ( .A1(n38231), .A2(\REGISTERS[27][2] ), .B1(n37743), .B2(
        \REGISTERS[4][2] ), .ZN(n38075) );
  AOI22_X1 U1381 ( .A1(n38233), .A2(\REGISTERS[10][2] ), .B1(n38232), .B2(
        \REGISTERS[28][2] ), .ZN(n38074) );
  AOI22_X1 U1382 ( .A1(n38235), .A2(\REGISTERS[6][2] ), .B1(n38234), .B2(
        \REGISTERS[7][2] ), .ZN(n38073) );
  NAND4_X1 U1383 ( .A1(n38076), .A2(n38075), .A3(n38074), .A4(n38073), .ZN(
        n38082) );
  AOI22_X1 U1384 ( .A1(n38241), .A2(\REGISTERS[26][2] ), .B1(n38240), .B2(
        \REGISTERS[5][2] ), .ZN(n38080) );
  AOI22_X1 U1385 ( .A1(n38243), .A2(\REGISTERS[21][2] ), .B1(n38242), .B2(
        \REGISTERS[25][2] ), .ZN(n38079) );
  AOI22_X1 U1386 ( .A1(n38245), .A2(\REGISTERS[23][2] ), .B1(n38244), .B2(
        \REGISTERS[17][2] ), .ZN(n38078) );
  AOI22_X1 U1387 ( .A1(n38247), .A2(\REGISTERS[14][2] ), .B1(n38246), .B2(
        \REGISTERS[19][2] ), .ZN(n38077) );
  NAND4_X1 U1388 ( .A1(n38080), .A2(n38079), .A3(n38078), .A4(n38077), .ZN(
        n38081) );
  AOI22_X1 U1389 ( .A1(n37727), .A2(\REGISTERS[11][30] ), .B1(n38205), .B2(
        \REGISTERS[16][30] ), .ZN(n38088) );
  AOI22_X1 U1390 ( .A1(n37729), .A2(\REGISTERS[1][30] ), .B1(n38207), .B2(
        \REGISTERS[24][30] ), .ZN(n38087) );
  AOI22_X1 U1391 ( .A1(n37731), .A2(\REGISTERS[12][30] ), .B1(n37730), .B2(
        \REGISTERS[15][30] ), .ZN(n38086) );
  NAND2_X1 U1392 ( .A1(n38211), .A2(\REGISTERS[13][30] ), .ZN(n38085) );
  NAND4_X1 U1393 ( .A1(n38088), .A2(n38087), .A3(n38086), .A4(n38085), .ZN(
        n38104) );
  AOI22_X1 U1394 ( .A1(n38217), .A2(\REGISTERS[20][30] ), .B1(n38216), .B2(
        \REGISTERS[22][30] ), .ZN(n38092) );
  AOI22_X1 U1395 ( .A1(n38219), .A2(\REGISTERS[18][30] ), .B1(n38218), .B2(
        \REGISTERS[9][30] ), .ZN(n38091) );
  AOI22_X1 U1396 ( .A1(n38221), .A2(\REGISTERS[2][30] ), .B1(n38220), .B2(
        \REGISTERS[31][30] ), .ZN(n38090) );
  AOI22_X1 U1397 ( .A1(n38223), .A2(\REGISTERS[3][30] ), .B1(n38222), .B2(
        \REGISTERS[8][30] ), .ZN(n38089) );
  NAND4_X1 U1398 ( .A1(n38092), .A2(n38091), .A3(n38090), .A4(n38089), .ZN(
        n38103) );
  AOI22_X1 U1399 ( .A1(n38229), .A2(\REGISTERS[30][30] ), .B1(n38228), .B2(
        \REGISTERS[29][30] ), .ZN(n38096) );
  AOI22_X1 U1400 ( .A1(n37744), .A2(\REGISTERS[27][30] ), .B1(n38230), .B2(
        \REGISTERS[4][30] ), .ZN(n38095) );
  AOI22_X1 U1401 ( .A1(n38233), .A2(\REGISTERS[10][30] ), .B1(n38232), .B2(
        \REGISTERS[28][30] ), .ZN(n38094) );
  AOI22_X1 U1402 ( .A1(n38235), .A2(\REGISTERS[6][30] ), .B1(n38234), .B2(
        \REGISTERS[7][30] ), .ZN(n38093) );
  NAND4_X1 U1403 ( .A1(n38096), .A2(n38095), .A3(n38094), .A4(n38093), .ZN(
        n38102) );
  AOI22_X1 U1404 ( .A1(n38241), .A2(\REGISTERS[26][30] ), .B1(n38240), .B2(
        \REGISTERS[5][30] ), .ZN(n38100) );
  AOI22_X1 U1405 ( .A1(n38243), .A2(\REGISTERS[21][30] ), .B1(n38242), .B2(
        \REGISTERS[25][30] ), .ZN(n38099) );
  AOI22_X1 U1406 ( .A1(n38245), .A2(\REGISTERS[23][30] ), .B1(n38244), .B2(
        \REGISTERS[17][30] ), .ZN(n38098) );
  AOI22_X1 U1407 ( .A1(n38247), .A2(\REGISTERS[14][30] ), .B1(n38246), .B2(
        \REGISTERS[19][30] ), .ZN(n38097) );
  NAND4_X1 U1408 ( .A1(n38100), .A2(n38099), .A3(n38098), .A4(n38097), .ZN(
        n38101) );
  AOI22_X1 U1409 ( .A1(n38206), .A2(\REGISTERS[11][31] ), .B1(n38205), .B2(
        \REGISTERS[16][31] ), .ZN(n38108) );
  AOI22_X1 U1410 ( .A1(n38208), .A2(\REGISTERS[1][31] ), .B1(n38207), .B2(
        \REGISTERS[24][31] ), .ZN(n38107) );
  AOI22_X1 U1411 ( .A1(n38210), .A2(\REGISTERS[12][31] ), .B1(n38209), .B2(
        \REGISTERS[15][31] ), .ZN(n38106) );
  NAND2_X1 U1412 ( .A1(n38211), .A2(\REGISTERS[13][31] ), .ZN(n38105) );
  NAND4_X1 U1413 ( .A1(n38108), .A2(n38107), .A3(n38106), .A4(n38105), .ZN(
        n38124) );
  AOI22_X1 U1414 ( .A1(n38217), .A2(\REGISTERS[20][31] ), .B1(n38216), .B2(
        \REGISTERS[22][31] ), .ZN(n38112) );
  AOI22_X1 U1415 ( .A1(n38219), .A2(\REGISTERS[18][31] ), .B1(n38218), .B2(
        \REGISTERS[9][31] ), .ZN(n38111) );
  AOI22_X1 U1416 ( .A1(n37738), .A2(\REGISTERS[2][31] ), .B1(n38220), .B2(
        \REGISTERS[31][31] ), .ZN(n38110) );
  AOI22_X1 U1417 ( .A1(n38223), .A2(\REGISTERS[3][31] ), .B1(n38222), .B2(
        \REGISTERS[8][31] ), .ZN(n38109) );
  NAND4_X1 U1418 ( .A1(n38112), .A2(n38111), .A3(n38110), .A4(n38109), .ZN(
        n38123) );
  AOI22_X1 U1419 ( .A1(n38229), .A2(\REGISTERS[30][31] ), .B1(n38228), .B2(
        \REGISTERS[29][31] ), .ZN(n38116) );
  AOI22_X1 U1420 ( .A1(n38231), .A2(\REGISTERS[27][31] ), .B1(n38230), .B2(
        \REGISTERS[4][31] ), .ZN(n38115) );
  AOI22_X1 U1421 ( .A1(n38233), .A2(\REGISTERS[10][31] ), .B1(n38232), .B2(
        \REGISTERS[28][31] ), .ZN(n38114) );
  AOI22_X1 U1422 ( .A1(n38235), .A2(\REGISTERS[6][31] ), .B1(n38234), .B2(
        \REGISTERS[7][31] ), .ZN(n38113) );
  NAND4_X1 U1423 ( .A1(n38116), .A2(n38115), .A3(n38114), .A4(n38113), .ZN(
        n38122) );
  AOI22_X1 U1424 ( .A1(n38241), .A2(\REGISTERS[26][31] ), .B1(n38240), .B2(
        \REGISTERS[5][31] ), .ZN(n38120) );
  AOI22_X1 U1425 ( .A1(n38243), .A2(\REGISTERS[21][31] ), .B1(n38242), .B2(
        \REGISTERS[25][31] ), .ZN(n38119) );
  AOI22_X1 U1426 ( .A1(n38245), .A2(\REGISTERS[23][31] ), .B1(n38244), .B2(
        \REGISTERS[17][31] ), .ZN(n38118) );
  AOI22_X1 U1427 ( .A1(n38247), .A2(\REGISTERS[14][31] ), .B1(n38246), .B2(
        \REGISTERS[19][31] ), .ZN(n38117) );
  NAND4_X1 U1428 ( .A1(n38120), .A2(n38119), .A3(n38118), .A4(n38117), .ZN(
        n38121) );
  AOI22_X1 U1429 ( .A1(n38206), .A2(\REGISTERS[11][3] ), .B1(n38205), .B2(
        \REGISTERS[16][3] ), .ZN(n38128) );
  AOI22_X1 U1430 ( .A1(n38208), .A2(\REGISTERS[1][3] ), .B1(n38207), .B2(
        \REGISTERS[24][3] ), .ZN(n38127) );
  AOI22_X1 U1431 ( .A1(n38210), .A2(\REGISTERS[12][3] ), .B1(n38209), .B2(
        \REGISTERS[15][3] ), .ZN(n38126) );
  NAND2_X1 U1432 ( .A1(n38211), .A2(\REGISTERS[13][3] ), .ZN(n38125) );
  NAND4_X1 U1433 ( .A1(n38128), .A2(n38127), .A3(n38126), .A4(n38125), .ZN(
        n38144) );
  AOI22_X1 U1434 ( .A1(n38217), .A2(\REGISTERS[20][3] ), .B1(n38216), .B2(
        \REGISTERS[22][3] ), .ZN(n38132) );
  AOI22_X1 U1435 ( .A1(n38219), .A2(\REGISTERS[18][3] ), .B1(n38218), .B2(
        \REGISTERS[9][3] ), .ZN(n38131) );
  AOI22_X1 U1436 ( .A1(n38221), .A2(\REGISTERS[2][3] ), .B1(n38220), .B2(
        \REGISTERS[31][3] ), .ZN(n38130) );
  AOI22_X1 U1437 ( .A1(n38223), .A2(\REGISTERS[3][3] ), .B1(n38222), .B2(
        \REGISTERS[8][3] ), .ZN(n38129) );
  NAND4_X1 U1438 ( .A1(n38132), .A2(n38131), .A3(n38130), .A4(n38129), .ZN(
        n38143) );
  AOI22_X1 U1439 ( .A1(n38229), .A2(\REGISTERS[30][3] ), .B1(n38228), .B2(
        \REGISTERS[29][3] ), .ZN(n38136) );
  AOI22_X1 U1440 ( .A1(n38231), .A2(\REGISTERS[27][3] ), .B1(n38230), .B2(
        \REGISTERS[4][3] ), .ZN(n38135) );
  AOI22_X1 U1441 ( .A1(n38233), .A2(\REGISTERS[10][3] ), .B1(n38232), .B2(
        \REGISTERS[28][3] ), .ZN(n38134) );
  AOI22_X1 U1442 ( .A1(n38235), .A2(\REGISTERS[6][3] ), .B1(n38234), .B2(
        \REGISTERS[7][3] ), .ZN(n38133) );
  NAND4_X1 U1443 ( .A1(n38136), .A2(n38135), .A3(n38134), .A4(n38133), .ZN(
        n38142) );
  AOI22_X1 U1444 ( .A1(n38241), .A2(\REGISTERS[26][3] ), .B1(n38240), .B2(
        \REGISTERS[5][3] ), .ZN(n38140) );
  AOI22_X1 U1445 ( .A1(n38243), .A2(\REGISTERS[21][3] ), .B1(n38242), .B2(
        \REGISTERS[25][3] ), .ZN(n38139) );
  AOI22_X1 U1446 ( .A1(n38245), .A2(\REGISTERS[23][3] ), .B1(n38244), .B2(
        \REGISTERS[17][3] ), .ZN(n38138) );
  AOI22_X1 U1447 ( .A1(n38247), .A2(\REGISTERS[14][3] ), .B1(n38246), .B2(
        \REGISTERS[19][3] ), .ZN(n38137) );
  NAND4_X1 U1448 ( .A1(n38140), .A2(n38139), .A3(n38138), .A4(n38137), .ZN(
        n38141) );
  AOI22_X1 U1449 ( .A1(n38206), .A2(\REGISTERS[11][5] ), .B1(n38205), .B2(
        \REGISTERS[16][5] ), .ZN(n38148) );
  AOI22_X1 U1450 ( .A1(n38208), .A2(\REGISTERS[1][5] ), .B1(n38207), .B2(
        \REGISTERS[24][5] ), .ZN(n38147) );
  AOI22_X1 U1451 ( .A1(n38210), .A2(\REGISTERS[12][5] ), .B1(n38209), .B2(
        \REGISTERS[15][5] ), .ZN(n38146) );
  NAND2_X1 U1452 ( .A1(n38211), .A2(\REGISTERS[13][5] ), .ZN(n38145) );
  NAND4_X1 U1453 ( .A1(n38148), .A2(n38147), .A3(n38146), .A4(n38145), .ZN(
        n38164) );
  AOI22_X1 U1454 ( .A1(n38217), .A2(\REGISTERS[20][5] ), .B1(n38216), .B2(
        \REGISTERS[22][5] ), .ZN(n38152) );
  AOI22_X1 U1455 ( .A1(n38219), .A2(\REGISTERS[18][5] ), .B1(n38218), .B2(
        \REGISTERS[9][5] ), .ZN(n38151) );
  AOI22_X1 U1456 ( .A1(n38221), .A2(\REGISTERS[2][5] ), .B1(n38220), .B2(
        \REGISTERS[31][5] ), .ZN(n38150) );
  AOI22_X1 U1457 ( .A1(n38223), .A2(\REGISTERS[3][5] ), .B1(n38222), .B2(
        \REGISTERS[8][5] ), .ZN(n38149) );
  NAND4_X1 U1458 ( .A1(n38152), .A2(n38151), .A3(n38150), .A4(n38149), .ZN(
        n38163) );
  AOI22_X1 U1459 ( .A1(n38229), .A2(\REGISTERS[30][5] ), .B1(n38228), .B2(
        \REGISTERS[29][5] ), .ZN(n38156) );
  AOI22_X1 U1460 ( .A1(n38231), .A2(\REGISTERS[27][5] ), .B1(n38230), .B2(
        \REGISTERS[4][5] ), .ZN(n38155) );
  AOI22_X1 U1461 ( .A1(n38233), .A2(\REGISTERS[10][5] ), .B1(n38232), .B2(
        \REGISTERS[28][5] ), .ZN(n38154) );
  AOI22_X1 U1462 ( .A1(n38235), .A2(\REGISTERS[6][5] ), .B1(n38234), .B2(
        \REGISTERS[7][5] ), .ZN(n38153) );
  NAND4_X1 U1463 ( .A1(n38156), .A2(n38155), .A3(n38154), .A4(n38153), .ZN(
        n38162) );
  AOI22_X1 U1464 ( .A1(n38241), .A2(\REGISTERS[26][5] ), .B1(n38240), .B2(
        \REGISTERS[5][5] ), .ZN(n38160) );
  AOI22_X1 U1465 ( .A1(n38243), .A2(\REGISTERS[21][5] ), .B1(n38242), .B2(
        \REGISTERS[25][5] ), .ZN(n38159) );
  AOI22_X1 U1466 ( .A1(n38245), .A2(\REGISTERS[23][5] ), .B1(n38244), .B2(
        \REGISTERS[17][5] ), .ZN(n38158) );
  AOI22_X1 U1467 ( .A1(n38247), .A2(\REGISTERS[14][5] ), .B1(n38246), .B2(
        \REGISTERS[19][5] ), .ZN(n38157) );
  NAND4_X1 U1468 ( .A1(n38160), .A2(n38159), .A3(n38158), .A4(n38157), .ZN(
        n38161) );
  AOI22_X1 U1469 ( .A1(n38206), .A2(\REGISTERS[11][6] ), .B1(n38205), .B2(
        \REGISTERS[16][6] ), .ZN(n38168) );
  AOI22_X1 U1470 ( .A1(n38208), .A2(\REGISTERS[1][6] ), .B1(n38207), .B2(
        \REGISTERS[24][6] ), .ZN(n38167) );
  AOI22_X1 U1471 ( .A1(n38210), .A2(\REGISTERS[12][6] ), .B1(n38209), .B2(
        \REGISTERS[15][6] ), .ZN(n38166) );
  NAND2_X1 U1472 ( .A1(n38211), .A2(\REGISTERS[13][6] ), .ZN(n38165) );
  NAND4_X1 U1473 ( .A1(n38168), .A2(n38167), .A3(n38166), .A4(n38165), .ZN(
        n38184) );
  AOI22_X1 U1474 ( .A1(n38217), .A2(\REGISTERS[20][6] ), .B1(n38216), .B2(
        \REGISTERS[22][6] ), .ZN(n38172) );
  AOI22_X1 U1475 ( .A1(n38219), .A2(\REGISTERS[18][6] ), .B1(n38218), .B2(
        \REGISTERS[9][6] ), .ZN(n38171) );
  AOI22_X1 U1476 ( .A1(n38221), .A2(\REGISTERS[2][6] ), .B1(n38220), .B2(
        \REGISTERS[31][6] ), .ZN(n38170) );
  AOI22_X1 U1477 ( .A1(n38223), .A2(\REGISTERS[3][6] ), .B1(n38222), .B2(
        \REGISTERS[8][6] ), .ZN(n38169) );
  NAND4_X1 U1478 ( .A1(n38172), .A2(n38171), .A3(n38170), .A4(n38169), .ZN(
        n38183) );
  AOI22_X1 U1479 ( .A1(n38229), .A2(\REGISTERS[30][6] ), .B1(n38228), .B2(
        \REGISTERS[29][6] ), .ZN(n38176) );
  AOI22_X1 U1480 ( .A1(n38231), .A2(\REGISTERS[27][6] ), .B1(n38230), .B2(
        \REGISTERS[4][6] ), .ZN(n38175) );
  AOI22_X1 U1481 ( .A1(n38233), .A2(\REGISTERS[10][6] ), .B1(n38232), .B2(
        \REGISTERS[28][6] ), .ZN(n38174) );
  AOI22_X1 U1482 ( .A1(n38235), .A2(\REGISTERS[6][6] ), .B1(n38234), .B2(
        \REGISTERS[7][6] ), .ZN(n38173) );
  NAND4_X1 U1483 ( .A1(n38176), .A2(n38175), .A3(n38174), .A4(n38173), .ZN(
        n38182) );
  AOI22_X1 U1484 ( .A1(n38241), .A2(\REGISTERS[26][6] ), .B1(n38240), .B2(
        \REGISTERS[5][6] ), .ZN(n38180) );
  AOI22_X1 U1485 ( .A1(n38243), .A2(\REGISTERS[21][6] ), .B1(n38242), .B2(
        \REGISTERS[25][6] ), .ZN(n38179) );
  AOI22_X1 U1486 ( .A1(n38245), .A2(\REGISTERS[23][6] ), .B1(n38244), .B2(
        \REGISTERS[17][6] ), .ZN(n38178) );
  AOI22_X1 U1487 ( .A1(n38247), .A2(\REGISTERS[14][6] ), .B1(n38246), .B2(
        \REGISTERS[19][6] ), .ZN(n38177) );
  NAND4_X1 U1488 ( .A1(n38180), .A2(n38179), .A3(n38178), .A4(n38177), .ZN(
        n38181) );
  AOI22_X1 U1489 ( .A1(n38206), .A2(\REGISTERS[11][8] ), .B1(n38205), .B2(
        \REGISTERS[16][8] ), .ZN(n38188) );
  AOI22_X1 U1490 ( .A1(n38208), .A2(\REGISTERS[1][8] ), .B1(n38207), .B2(
        \REGISTERS[24][8] ), .ZN(n38187) );
  AOI22_X1 U1491 ( .A1(n38210), .A2(\REGISTERS[12][8] ), .B1(n38209), .B2(
        \REGISTERS[15][8] ), .ZN(n38186) );
  NAND2_X1 U1492 ( .A1(n37732), .A2(\REGISTERS[13][8] ), .ZN(n38185) );
  NAND4_X1 U1493 ( .A1(n38188), .A2(n38187), .A3(n38186), .A4(n38185), .ZN(
        n38204) );
  AOI22_X1 U1494 ( .A1(n38217), .A2(\REGISTERS[20][8] ), .B1(n38216), .B2(
        \REGISTERS[22][8] ), .ZN(n38192) );
  AOI22_X1 U1495 ( .A1(n38219), .A2(\REGISTERS[18][8] ), .B1(n38218), .B2(
        \REGISTERS[9][8] ), .ZN(n38191) );
  AOI22_X1 U1496 ( .A1(n37738), .A2(\REGISTERS[2][8] ), .B1(n38220), .B2(
        \REGISTERS[31][8] ), .ZN(n38190) );
  AOI22_X1 U1497 ( .A1(n38223), .A2(\REGISTERS[3][8] ), .B1(n38222), .B2(
        \REGISTERS[8][8] ), .ZN(n38189) );
  NAND4_X1 U1498 ( .A1(n38192), .A2(n38191), .A3(n38190), .A4(n38189), .ZN(
        n38203) );
  AOI22_X1 U1499 ( .A1(n38229), .A2(\REGISTERS[30][8] ), .B1(n38228), .B2(
        \REGISTERS[29][8] ), .ZN(n38196) );
  AOI22_X1 U1500 ( .A1(n38231), .A2(\REGISTERS[27][8] ), .B1(n37743), .B2(
        \REGISTERS[4][8] ), .ZN(n38195) );
  AOI22_X1 U1501 ( .A1(n38233), .A2(\REGISTERS[10][8] ), .B1(n38232), .B2(
        \REGISTERS[28][8] ), .ZN(n38194) );
  AOI22_X1 U1502 ( .A1(n38235), .A2(\REGISTERS[6][8] ), .B1(n38234), .B2(
        \REGISTERS[7][8] ), .ZN(n38193) );
  NAND4_X1 U1503 ( .A1(n38196), .A2(n38195), .A3(n38194), .A4(n38193), .ZN(
        n38202) );
  AOI22_X1 U1504 ( .A1(n38241), .A2(\REGISTERS[26][8] ), .B1(n38240), .B2(
        \REGISTERS[5][8] ), .ZN(n38200) );
  AOI22_X1 U1505 ( .A1(n38243), .A2(\REGISTERS[21][8] ), .B1(n38242), .B2(
        \REGISTERS[25][8] ), .ZN(n38199) );
  AOI22_X1 U1506 ( .A1(n38245), .A2(\REGISTERS[23][8] ), .B1(n38244), .B2(
        \REGISTERS[17][8] ), .ZN(n38198) );
  AOI22_X1 U1507 ( .A1(n38247), .A2(\REGISTERS[14][8] ), .B1(n38246), .B2(
        \REGISTERS[19][8] ), .ZN(n38197) );
  NAND4_X1 U1508 ( .A1(n38200), .A2(n38199), .A3(n38198), .A4(n38197), .ZN(
        n38201) );
  AOI22_X1 U1509 ( .A1(n38206), .A2(\REGISTERS[11][9] ), .B1(n38205), .B2(
        \REGISTERS[16][9] ), .ZN(n38215) );
  AOI22_X1 U1510 ( .A1(n38208), .A2(\REGISTERS[1][9] ), .B1(n38207), .B2(
        \REGISTERS[24][9] ), .ZN(n38214) );
  AOI22_X1 U1511 ( .A1(n38210), .A2(\REGISTERS[12][9] ), .B1(n38209), .B2(
        \REGISTERS[15][9] ), .ZN(n38213) );
  NAND2_X1 U1512 ( .A1(n37732), .A2(\REGISTERS[13][9] ), .ZN(n38212) );
  NAND4_X1 U1513 ( .A1(n38215), .A2(n38214), .A3(n38213), .A4(n38212), .ZN(
        n38255) );
  AOI22_X1 U1514 ( .A1(n38217), .A2(\REGISTERS[20][9] ), .B1(n38216), .B2(
        \REGISTERS[22][9] ), .ZN(n38227) );
  AOI22_X1 U1515 ( .A1(n38219), .A2(\REGISTERS[18][9] ), .B1(n38218), .B2(
        \REGISTERS[9][9] ), .ZN(n38226) );
  AOI22_X1 U1516 ( .A1(n37738), .A2(\REGISTERS[2][9] ), .B1(n37737), .B2(
        \REGISTERS[31][9] ), .ZN(n38225) );
  AOI22_X1 U1517 ( .A1(n38223), .A2(\REGISTERS[3][9] ), .B1(n38222), .B2(
        \REGISTERS[8][9] ), .ZN(n38224) );
  NAND4_X1 U1518 ( .A1(n38227), .A2(n38226), .A3(n38225), .A4(n38224), .ZN(
        n38254) );
  AOI22_X1 U1519 ( .A1(n38229), .A2(\REGISTERS[30][9] ), .B1(n37741), .B2(
        \REGISTERS[29][9] ), .ZN(n38239) );
  AOI22_X1 U1520 ( .A1(n38231), .A2(\REGISTERS[27][9] ), .B1(n37743), .B2(
        \REGISTERS[4][9] ), .ZN(n38238) );
  AOI22_X1 U1521 ( .A1(n38233), .A2(\REGISTERS[10][9] ), .B1(n37745), .B2(
        \REGISTERS[28][9] ), .ZN(n38237) );
  AOI22_X1 U1522 ( .A1(n38235), .A2(\REGISTERS[6][9] ), .B1(n38234), .B2(
        \REGISTERS[7][9] ), .ZN(n38236) );
  NAND4_X1 U1523 ( .A1(n38239), .A2(n38238), .A3(n38237), .A4(n38236), .ZN(
        n38253) );
  AOI22_X1 U1524 ( .A1(n38241), .A2(\REGISTERS[26][9] ), .B1(n37749), .B2(
        \REGISTERS[5][9] ), .ZN(n38251) );
  AOI22_X1 U1525 ( .A1(n38243), .A2(\REGISTERS[21][9] ), .B1(n38242), .B2(
        \REGISTERS[25][9] ), .ZN(n38250) );
  AOI22_X1 U1526 ( .A1(n38245), .A2(\REGISTERS[23][9] ), .B1(n38244), .B2(
        \REGISTERS[17][9] ), .ZN(n38249) );
  AOI22_X1 U1527 ( .A1(n38247), .A2(\REGISTERS[14][9] ), .B1(n38246), .B2(
        \REGISTERS[19][9] ), .ZN(n38248) );
  NAND4_X1 U1528 ( .A1(n38251), .A2(n38250), .A3(n38249), .A4(n38248), .ZN(
        n38252) );
  INV_X1 U1529 ( .A(ADD_RDB[2]), .ZN(n38260) );
  NAND3_X1 U1530 ( .A1(RESET), .A2(ADD_RDB[1]), .A3(n38260), .ZN(n38270) );
  INV_X1 U1531 ( .A(ADD_RDB[4]), .ZN(n38259) );
  NAND3_X1 U1532 ( .A1(ADD_RDB[3]), .A2(ADD_RDB[0]), .A3(n38259), .ZN(n38262)
         );
  NOR2_X1 U1533 ( .A1(n38270), .A2(n38262), .ZN(n38276) );
  NAND3_X1 U1534 ( .A1(ADD_RDB[4]), .A2(ADD_RDB[3]), .A3(ADD_RDB[0]), .ZN(
        n38267) );
  INV_X1 U1535 ( .A(ADD_RDB[1]), .ZN(n38256) );
  NAND3_X1 U1536 ( .A1(RESET), .A2(n38260), .A3(n38256), .ZN(n38266) );
  NOR2_X1 U1537 ( .A1(n38267), .A2(n38266), .ZN(n38275) );
  NOR2_X1 U1538 ( .A1(ADD_RDB[3]), .A2(ADD_RDB[0]), .ZN(n38261) );
  NAND3_X1 U1539 ( .A1(RESET), .A2(n38261), .A3(n38259), .ZN(n38264) );
  NOR3_X1 U1540 ( .A1(ADD_RDB[2]), .A2(n38256), .A3(n38264), .ZN(n38278) );
  NAND3_X1 U1541 ( .A1(RESET), .A2(ADD_RDB[2]), .A3(ADD_RDB[1]), .ZN(n38271)
         );
  NAND3_X1 U1542 ( .A1(ADD_RDB[2]), .A2(RESET), .A3(n38256), .ZN(n38274) );
  NOR2_X1 U1543 ( .A1(n38262), .A2(n38274), .ZN(n38280) );
  NOR2_X1 U1544 ( .A1(n38267), .A2(n38274), .ZN(n38279) );
  INV_X1 U1545 ( .A(ADD_RDB[3]), .ZN(n38258) );
  NAND3_X1 U1546 ( .A1(ADD_RDB[4]), .A2(ADD_RDB[0]), .A3(n38258), .ZN(n38268)
         );
  NOR2_X1 U1547 ( .A1(n38270), .A2(n38268), .ZN(n38281) );
  INV_X1 U1548 ( .A(ADD_RDB[0]), .ZN(n38257) );
  NAND3_X1 U1549 ( .A1(ADD_RDB[3]), .A2(n38259), .A3(n38257), .ZN(n38265) );
  NOR2_X1 U1550 ( .A1(n38266), .A2(n38265), .ZN(n38283) );
  NAND3_X1 U1551 ( .A1(ADD_RDB[3]), .A2(ADD_RDB[4]), .A3(n38257), .ZN(n38272)
         );
  NOR2_X1 U1552 ( .A1(n38270), .A2(n38272), .ZN(n38282) );
  NAND3_X1 U1553 ( .A1(ADD_RDB[0]), .A2(n38259), .A3(n38258), .ZN(n38273) );
  NOR2_X1 U1554 ( .A1(n38270), .A2(n38273), .ZN(n38285) );
  NOR2_X1 U1555 ( .A1(n38271), .A2(n38272), .ZN(n38284) );
  NOR3_X1 U1556 ( .A1(ADD_RDB[1]), .A2(n38260), .A3(n38264), .ZN(n38287) );
  NOR2_X1 U1557 ( .A1(n38268), .A2(n38266), .ZN(n38286) );
  NAND2_X1 U1558 ( .A1(ADD_RDB[4]), .A2(n38261), .ZN(n38269) );
  NOR2_X1 U1559 ( .A1(n38271), .A2(n38269), .ZN(n38288) );
  NOR2_X1 U1560 ( .A1(n38266), .A2(n38269), .ZN(n38291) );
  NOR2_X1 U1561 ( .A1(n38262), .A2(n38266), .ZN(n38290) );
  NAND2_X1 U1562 ( .A1(ADD_RDB[2]), .A2(ADD_RDB[1]), .ZN(n38263) );
  NOR2_X1 U1563 ( .A1(n38264), .A2(n38263), .ZN(n38293) );
  NOR2_X1 U1564 ( .A1(n38268), .A2(n38271), .ZN(n38292) );
  NOR2_X1 U1565 ( .A1(n38266), .A2(n38272), .ZN(n38295) );
  NOR2_X1 U1566 ( .A1(n38271), .A2(n38265), .ZN(n38294) );
  NOR2_X1 U1567 ( .A1(n38274), .A2(n38265), .ZN(n38297) );
  NOR2_X1 U1568 ( .A1(n38270), .A2(n38265), .ZN(n38296) );
  NOR2_X1 U1569 ( .A1(n38266), .A2(n38273), .ZN(n38299) );
  NOR2_X1 U1570 ( .A1(n38270), .A2(n38267), .ZN(n38298) );
  NOR2_X1 U1571 ( .A1(n38274), .A2(n38269), .ZN(n38301) );
  NOR2_X1 U1572 ( .A1(n38268), .A2(n38274), .ZN(n38300) );
  NOR2_X1 U1573 ( .A1(n38270), .A2(n38269), .ZN(n38303) );
  NOR2_X1 U1574 ( .A1(n38271), .A2(n38273), .ZN(n38302) );
  NOR2_X1 U1575 ( .A1(n38274), .A2(n38272), .ZN(n38305) );
  NOR2_X1 U1576 ( .A1(n38274), .A2(n38273), .ZN(n38304) );
endmodule


module branch_predictor ( RST, PC_IN, PC_FAIL, IR_IN, IR_FAIL, WRONG_PRE, 
        RIGHT_PRE, NPC_OUT, LINK_ADD, SEL, TAKEN );
  input [31:0] PC_IN;
  input [31:0] PC_FAIL;
  input [31:0] IR_IN;
  input [15:0] IR_FAIL;
  output [31:0] NPC_OUT;
  output [31:0] LINK_ADD;
  input RST, WRONG_PRE, RIGHT_PRE;
  output SEL, TAKEN;
  wire   \CACHE_mem[0][1] , \CACHE_mem[0][0] , \CACHE_mem[1][1] ,
         \CACHE_mem[1][0] , \CACHE_mem[2][1] , \CACHE_mem[2][0] ,
         \CACHE_mem[3][1] , \CACHE_mem[3][0] , \CACHE_mem[4][1] ,
         \CACHE_mem[4][0] , \CACHE_mem[5][1] , \CACHE_mem[5][0] ,
         \CACHE_mem[6][1] , \CACHE_mem[6][0] , \CACHE_mem[7][1] ,
         \CACHE_mem[7][0] , \CACHE_mem[8][1] , \CACHE_mem[8][0] ,
         \CACHE_mem[9][1] , \CACHE_mem[9][0] , \CACHE_mem[10][1] ,
         \CACHE_mem[10][0] , \CACHE_mem[11][1] , \CACHE_mem[11][0] ,
         \CACHE_mem[12][1] , \CACHE_mem[12][0] , \CACHE_mem[13][1] ,
         \CACHE_mem[13][0] , \CACHE_mem[14][1] , \CACHE_mem[14][0] ,
         \CACHE_mem[15][1] , \CACHE_mem[15][0] , \CACHE_mem[16][1] ,
         \CACHE_mem[16][0] , \CACHE_mem[17][1] , \CACHE_mem[17][0] ,
         \CACHE_mem[18][1] , \CACHE_mem[18][0] , \CACHE_mem[19][1] ,
         \CACHE_mem[19][0] , \CACHE_mem[20][1] , \CACHE_mem[20][0] ,
         \CACHE_mem[21][1] , \CACHE_mem[21][0] , \CACHE_mem[22][1] ,
         \CACHE_mem[22][0] , \CACHE_mem[23][1] , \CACHE_mem[23][0] ,
         \CACHE_mem[24][1] , \CACHE_mem[24][0] , \CACHE_mem[25][1] ,
         \CACHE_mem[25][0] , \CACHE_mem[26][1] , \CACHE_mem[26][0] ,
         \CACHE_mem[27][1] , \CACHE_mem[27][0] , \CACHE_mem[28][1] ,
         \CACHE_mem[28][0] , \CACHE_mem[29][1] , \CACHE_mem[29][0] ,
         \CACHE_mem[30][1] , \CACHE_mem[30][0] , \CACHE_mem[31][1] ,
         \CACHE_mem[31][0] , N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N323, N356, N357, N358, N362, N387, N388, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n60,
         \add_65/carry[31] , \add_65/carry[30] , \add_65/carry[29] ,
         \add_65/carry[28] , \add_65/carry[27] , \add_65/carry[26] ,
         \add_65/carry[25] , \add_65/carry[24] , \add_65/carry[23] ,
         \add_65/carry[22] , \add_65/carry[21] , \add_65/carry[20] ,
         \add_65/carry[19] , \add_65/carry[18] , \add_65/carry[17] ,
         \add_65/carry[16] , \add_65/carry[15] , \add_65/carry[14] ,
         \add_65/carry[13] , \add_65/carry[12] , \add_65/carry[11] ,
         \add_65/carry[10] , \add_65/carry[9] , \add_65/carry[8] ,
         \add_65/carry[7] , \add_65/carry[6] , \add_65/carry[5] ,
         \add_65/carry[4] , \add_65/carry[3] , \add_65/carry[2] , \add_59/n1 ,
         \add_59/carry[31] , \add_59/carry[30] , \add_59/carry[29] ,
         \add_59/carry[28] , \add_59/carry[27] , \add_59/carry[26] ,
         \add_59/carry[25] , \add_59/carry[24] , \add_59/carry[23] ,
         \add_59/carry[22] , \add_59/carry[21] , \add_59/carry[20] ,
         \add_59/carry[19] , \add_59/carry[18] , \add_59/carry[17] ,
         \add_59/carry[16] , \add_59/carry[15] , \add_59/carry[14] ,
         \add_59/carry[13] , \add_59/carry[12] , \add_59/carry[11] ,
         \add_59/carry[10] , \add_59/carry[9] , \add_59/carry[8] ,
         \add_59/carry[7] , \add_59/carry[6] , \add_59/carry[5] ,
         \add_59/carry[4] , \add_59/carry[3] , \add_59/carry[2] ,
         \add_53_aco/n2 , \add_53_aco/carry[31] , \add_53_aco/carry[30] ,
         \add_53_aco/carry[29] , \add_53_aco/carry[28] ,
         \add_53_aco/carry[27] , \add_53_aco/carry[26] ,
         \add_53_aco/carry[25] , \add_53_aco/carry[24] ,
         \add_53_aco/carry[23] , \add_53_aco/carry[22] ,
         \add_53_aco/carry[21] , \add_53_aco/carry[20] ,
         \add_53_aco/carry[19] , \add_53_aco/carry[18] ,
         \add_53_aco/carry[17] , \add_53_aco/carry[16] ,
         \add_53_aco/carry[15] , \add_53_aco/carry[14] ,
         \add_53_aco/carry[13] , \add_53_aco/carry[12] ,
         \add_53_aco/carry[11] , \add_53_aco/carry[10] , \add_53_aco/carry[9] ,
         \add_53_aco/carry[8] , \add_53_aco/carry[7] , \add_53_aco/carry[6] ,
         \add_53_aco/carry[5] , \add_53_aco/carry[4] , \add_53_aco/carry[3] ,
         \add_53_aco/carry[2] , n62, n286, n291, n59, n1, n2, n3, n4, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n280, n281, n282, n283,
         n284, n285, n287, n288, n289, n290, n292, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549;
  assign N113 = PC_IN[0];
  assign N114 = PC_IN[1];

  DLH_X1 \NPC_OUT_reg[31]  ( .G(N323), .D(n1), .Q(NPC_OUT[31]) );
  DLH_X1 \NPC_OUT_reg[30]  ( .G(N323), .D(n2), .Q(NPC_OUT[30]) );
  DLH_X1 \NPC_OUT_reg[29]  ( .G(N323), .D(n3), .Q(NPC_OUT[29]) );
  DLH_X1 \NPC_OUT_reg[28]  ( .G(N323), .D(n4), .Q(NPC_OUT[28]) );
  DLH_X1 \NPC_OUT_reg[27]  ( .G(N323), .D(n20), .Q(NPC_OUT[27]) );
  DLH_X1 \NPC_OUT_reg[26]  ( .G(N323), .D(n21), .Q(NPC_OUT[26]) );
  DLH_X1 \NPC_OUT_reg[25]  ( .G(N323), .D(n22), .Q(NPC_OUT[25]) );
  DLH_X1 \NPC_OUT_reg[24]  ( .G(N323), .D(n23), .Q(NPC_OUT[24]) );
  DLH_X1 \NPC_OUT_reg[23]  ( .G(N323), .D(n24), .Q(NPC_OUT[23]) );
  DLH_X1 \NPC_OUT_reg[22]  ( .G(N323), .D(n25), .Q(NPC_OUT[22]) );
  DLH_X1 \NPC_OUT_reg[21]  ( .G(N323), .D(n26), .Q(NPC_OUT[21]) );
  DLH_X1 \NPC_OUT_reg[20]  ( .G(N323), .D(n27), .Q(NPC_OUT[20]) );
  DLH_X1 \NPC_OUT_reg[19]  ( .G(N323), .D(n28), .Q(NPC_OUT[19]) );
  DLH_X1 \NPC_OUT_reg[18]  ( .G(N323), .D(n29), .Q(NPC_OUT[18]) );
  DLH_X1 \NPC_OUT_reg[17]  ( .G(N323), .D(n30), .Q(NPC_OUT[17]) );
  DLH_X1 \NPC_OUT_reg[16]  ( .G(N323), .D(n31), .Q(NPC_OUT[16]) );
  DLH_X1 \NPC_OUT_reg[15]  ( .G(N323), .D(n32), .Q(NPC_OUT[15]) );
  DLH_X1 \NPC_OUT_reg[14]  ( .G(N323), .D(n33), .Q(NPC_OUT[14]) );
  DLH_X1 \NPC_OUT_reg[13]  ( .G(N323), .D(n34), .Q(NPC_OUT[13]) );
  DLH_X1 \NPC_OUT_reg[12]  ( .G(N323), .D(n35), .Q(NPC_OUT[12]) );
  DLH_X1 \NPC_OUT_reg[11]  ( .G(N323), .D(n36), .Q(NPC_OUT[11]) );
  DLH_X1 \NPC_OUT_reg[10]  ( .G(N323), .D(n37), .Q(NPC_OUT[10]) );
  DLH_X1 \NPC_OUT_reg[9]  ( .G(N323), .D(n38), .Q(NPC_OUT[9]) );
  DLH_X1 \NPC_OUT_reg[8]  ( .G(N323), .D(n39), .Q(NPC_OUT[8]) );
  DLH_X1 \NPC_OUT_reg[7]  ( .G(N323), .D(n40), .Q(NPC_OUT[7]) );
  DLH_X1 \NPC_OUT_reg[6]  ( .G(N323), .D(n41), .Q(NPC_OUT[6]) );
  DLH_X1 \NPC_OUT_reg[5]  ( .G(N323), .D(n42), .Q(NPC_OUT[5]) );
  DLH_X1 \NPC_OUT_reg[4]  ( .G(N323), .D(n43), .Q(NPC_OUT[4]) );
  DLH_X1 \NPC_OUT_reg[3]  ( .G(N323), .D(n44), .Q(NPC_OUT[3]) );
  DLH_X1 \NPC_OUT_reg[2]  ( .G(N323), .D(n45), .Q(NPC_OUT[2]) );
  DLH_X1 \NPC_OUT_reg[1]  ( .G(N323), .D(n46), .Q(NPC_OUT[1]) );
  DLH_X1 \NPC_OUT_reg[0]  ( .G(N323), .D(n60), .Q(NPC_OUT[0]) );
  DLH_X1 \LINK_ADD_reg[31]  ( .G(N356), .D(N388), .Q(LINK_ADD[31]) );
  DLH_X1 \LINK_ADD_reg[30]  ( .G(N356), .D(N387), .Q(LINK_ADD[30]) );
  DLH_X1 \LINK_ADD_reg[29]  ( .G(n5323), .D(n58), .Q(LINK_ADD[29]) );
  DLH_X1 \LINK_ADD_reg[28]  ( .G(n5323), .D(n282), .Q(LINK_ADD[28]) );
  DLH_X1 \LINK_ADD_reg[27]  ( .G(n5323), .D(n57), .Q(LINK_ADD[27]) );
  DLH_X1 \LINK_ADD_reg[26]  ( .G(n5323), .D(n288), .Q(LINK_ADD[26]) );
  DLH_X1 \LINK_ADD_reg[25]  ( .G(n5323), .D(n56), .Q(LINK_ADD[25]) );
  DLH_X1 \LINK_ADD_reg[24]  ( .G(n5323), .D(n287), .Q(LINK_ADD[24]) );
  DLH_X1 \LINK_ADD_reg[23]  ( .G(n5323), .D(n55), .Q(LINK_ADD[23]) );
  DLH_X1 \LINK_ADD_reg[22]  ( .G(n5323), .D(n292), .Q(LINK_ADD[22]) );
  DLH_X1 \LINK_ADD_reg[21]  ( .G(n5323), .D(n54), .Q(LINK_ADD[21]) );
  DLH_X1 \LINK_ADD_reg[20]  ( .G(n5323), .D(n290), .Q(LINK_ADD[20]) );
  DLH_X1 \LINK_ADD_reg[19]  ( .G(n5323), .D(n53), .Q(LINK_ADD[19]) );
  DLH_X1 \LINK_ADD_reg[18]  ( .G(n5323), .D(n283), .Q(LINK_ADD[18]) );
  DLH_X1 \LINK_ADD_reg[17]  ( .G(n5323), .D(n52), .Q(LINK_ADD[17]) );
  DLH_X1 \LINK_ADD_reg[16]  ( .G(n5323), .D(n289), .Q(LINK_ADD[16]) );
  DLH_X1 \LINK_ADD_reg[15]  ( .G(n5323), .D(n51), .Q(LINK_ADD[15]) );
  DLH_X1 \LINK_ADD_reg[14]  ( .G(n5323), .D(n281), .Q(LINK_ADD[14]) );
  DLH_X1 \LINK_ADD_reg[13]  ( .G(n5323), .D(n50), .Q(LINK_ADD[13]) );
  DLH_X1 \LINK_ADD_reg[12]  ( .G(n5323), .D(n284), .Q(LINK_ADD[12]) );
  DLH_X1 \LINK_ADD_reg[11]  ( .G(n5323), .D(n49), .Q(LINK_ADD[11]) );
  DLH_X1 \LINK_ADD_reg[10]  ( .G(n5323), .D(n285), .Q(LINK_ADD[10]) );
  DLH_X1 \LINK_ADD_reg[9]  ( .G(n5323), .D(n48), .Q(LINK_ADD[9]) );
  DLH_X1 \LINK_ADD_reg[8]  ( .G(n5323), .D(n280), .Q(LINK_ADD[8]) );
  DLH_X1 \LINK_ADD_reg[7]  ( .G(N356), .D(n47), .Q(LINK_ADD[7]) );
  DLH_X1 \LINK_ADD_reg[6]  ( .G(N356), .D(n291), .Q(LINK_ADD[6]) );
  DLH_X1 \LINK_ADD_reg[5]  ( .G(N356), .D(N362), .Q(LINK_ADD[5]) );
  DLH_X1 \LINK_ADD_reg[4]  ( .G(N356), .D(n286), .Q(LINK_ADD[4]) );
  DLH_X1 \LINK_ADD_reg[3]  ( .G(N356), .D(n59), .Q(LINK_ADD[3]) );
  DLH_X1 \LINK_ADD_reg[2]  ( .G(N356), .D(n62), .Q(LINK_ADD[2]) );
  DLH_X1 \LINK_ADD_reg[1]  ( .G(N356), .D(N358), .Q(LINK_ADD[1]) );
  DLH_X1 \LINK_ADD_reg[0]  ( .G(N356), .D(N357), .Q(LINK_ADD[0]) );
  DLH_X1 \CACHE_mem_reg[0][1]  ( .G(N643), .D(N645), .Q(\CACHE_mem[0][1] ) );
  DLH_X1 \CACHE_mem_reg[0][0]  ( .G(N643), .D(N644), .Q(\CACHE_mem[0][0] ) );
  DLH_X1 \CACHE_mem_reg[1][1]  ( .G(N642), .D(N645), .Q(\CACHE_mem[1][1] ) );
  DLH_X1 \CACHE_mem_reg[1][0]  ( .G(N642), .D(N644), .Q(\CACHE_mem[1][0] ) );
  DLH_X1 \CACHE_mem_reg[2][1]  ( .G(N641), .D(N645), .Q(\CACHE_mem[2][1] ) );
  DLH_X1 \CACHE_mem_reg[2][0]  ( .G(N641), .D(N644), .Q(\CACHE_mem[2][0] ) );
  DLH_X1 \CACHE_mem_reg[3][1]  ( .G(N640), .D(N645), .Q(\CACHE_mem[3][1] ) );
  DLH_X1 \CACHE_mem_reg[3][0]  ( .G(N640), .D(N644), .Q(\CACHE_mem[3][0] ) );
  DLH_X1 \CACHE_mem_reg[4][1]  ( .G(N639), .D(N645), .Q(\CACHE_mem[4][1] ) );
  DLH_X1 \CACHE_mem_reg[4][0]  ( .G(N639), .D(N644), .Q(\CACHE_mem[4][0] ) );
  DLH_X1 \CACHE_mem_reg[5][1]  ( .G(N638), .D(N645), .Q(\CACHE_mem[5][1] ) );
  DLH_X1 \CACHE_mem_reg[5][0]  ( .G(N638), .D(N644), .Q(\CACHE_mem[5][0] ) );
  DLH_X1 \CACHE_mem_reg[6][1]  ( .G(N637), .D(N645), .Q(\CACHE_mem[6][1] ) );
  DLH_X1 \CACHE_mem_reg[6][0]  ( .G(N637), .D(N644), .Q(\CACHE_mem[6][0] ) );
  DLH_X1 \CACHE_mem_reg[7][1]  ( .G(N636), .D(N645), .Q(\CACHE_mem[7][1] ) );
  DLH_X1 \CACHE_mem_reg[7][0]  ( .G(N636), .D(N644), .Q(\CACHE_mem[7][0] ) );
  DLH_X1 \CACHE_mem_reg[8][1]  ( .G(N635), .D(N645), .Q(\CACHE_mem[8][1] ) );
  DLH_X1 \CACHE_mem_reg[8][0]  ( .G(N635), .D(N644), .Q(\CACHE_mem[8][0] ) );
  DLH_X1 \CACHE_mem_reg[9][1]  ( .G(N634), .D(N645), .Q(\CACHE_mem[9][1] ) );
  DLH_X1 \CACHE_mem_reg[9][0]  ( .G(N634), .D(N644), .Q(\CACHE_mem[9][0] ) );
  DLH_X1 \CACHE_mem_reg[10][1]  ( .G(N633), .D(N645), .Q(\CACHE_mem[10][1] )
         );
  DLH_X1 \CACHE_mem_reg[10][0]  ( .G(N633), .D(N644), .Q(\CACHE_mem[10][0] )
         );
  DLH_X1 \CACHE_mem_reg[11][1]  ( .G(N632), .D(N645), .Q(\CACHE_mem[11][1] )
         );
  DLH_X1 \CACHE_mem_reg[11][0]  ( .G(N632), .D(N644), .Q(\CACHE_mem[11][0] )
         );
  DLH_X1 \CACHE_mem_reg[12][1]  ( .G(N631), .D(N645), .Q(\CACHE_mem[12][1] )
         );
  DLH_X1 \CACHE_mem_reg[12][0]  ( .G(N631), .D(N644), .Q(\CACHE_mem[12][0] )
         );
  DLH_X1 \CACHE_mem_reg[13][1]  ( .G(N630), .D(N645), .Q(\CACHE_mem[13][1] )
         );
  DLH_X1 \CACHE_mem_reg[13][0]  ( .G(N630), .D(N644), .Q(\CACHE_mem[13][0] )
         );
  DLH_X1 \CACHE_mem_reg[14][1]  ( .G(N629), .D(N645), .Q(\CACHE_mem[14][1] )
         );
  DLH_X1 \CACHE_mem_reg[14][0]  ( .G(N629), .D(N644), .Q(\CACHE_mem[14][0] )
         );
  DLH_X1 \CACHE_mem_reg[15][1]  ( .G(N628), .D(N645), .Q(\CACHE_mem[15][1] )
         );
  DLH_X1 \CACHE_mem_reg[15][0]  ( .G(N628), .D(N644), .Q(\CACHE_mem[15][0] )
         );
  DLH_X1 \CACHE_mem_reg[16][1]  ( .G(N627), .D(N645), .Q(\CACHE_mem[16][1] )
         );
  DLH_X1 \CACHE_mem_reg[16][0]  ( .G(N627), .D(N644), .Q(\CACHE_mem[16][0] )
         );
  DLH_X1 \CACHE_mem_reg[17][1]  ( .G(N626), .D(N645), .Q(\CACHE_mem[17][1] )
         );
  DLH_X1 \CACHE_mem_reg[17][0]  ( .G(N626), .D(N644), .Q(\CACHE_mem[17][0] )
         );
  DLH_X1 \CACHE_mem_reg[18][1]  ( .G(N625), .D(N645), .Q(\CACHE_mem[18][1] )
         );
  DLH_X1 \CACHE_mem_reg[18][0]  ( .G(N625), .D(N644), .Q(\CACHE_mem[18][0] )
         );
  DLH_X1 \CACHE_mem_reg[19][1]  ( .G(N624), .D(N645), .Q(\CACHE_mem[19][1] )
         );
  DLH_X1 \CACHE_mem_reg[19][0]  ( .G(N624), .D(N644), .Q(\CACHE_mem[19][0] )
         );
  DLH_X1 \CACHE_mem_reg[20][1]  ( .G(N623), .D(N645), .Q(\CACHE_mem[20][1] )
         );
  DLH_X1 \CACHE_mem_reg[20][0]  ( .G(N623), .D(N644), .Q(\CACHE_mem[20][0] )
         );
  DLH_X1 \CACHE_mem_reg[21][1]  ( .G(N622), .D(N645), .Q(\CACHE_mem[21][1] )
         );
  DLH_X1 \CACHE_mem_reg[21][0]  ( .G(N622), .D(N644), .Q(\CACHE_mem[21][0] )
         );
  DLH_X1 \CACHE_mem_reg[22][1]  ( .G(N621), .D(N645), .Q(\CACHE_mem[22][1] )
         );
  DLH_X1 \CACHE_mem_reg[22][0]  ( .G(N621), .D(N644), .Q(\CACHE_mem[22][0] )
         );
  DLH_X1 \CACHE_mem_reg[23][1]  ( .G(N620), .D(N645), .Q(\CACHE_mem[23][1] )
         );
  DLH_X1 \CACHE_mem_reg[23][0]  ( .G(N620), .D(N644), .Q(\CACHE_mem[23][0] )
         );
  DLH_X1 \CACHE_mem_reg[24][1]  ( .G(N619), .D(N645), .Q(\CACHE_mem[24][1] )
         );
  DLH_X1 \CACHE_mem_reg[24][0]  ( .G(N619), .D(N644), .Q(\CACHE_mem[24][0] )
         );
  DLH_X1 \CACHE_mem_reg[25][1]  ( .G(N618), .D(N645), .Q(\CACHE_mem[25][1] )
         );
  DLH_X1 \CACHE_mem_reg[25][0]  ( .G(N618), .D(N644), .Q(\CACHE_mem[25][0] )
         );
  DLH_X1 \CACHE_mem_reg[26][1]  ( .G(N617), .D(N645), .Q(\CACHE_mem[26][1] )
         );
  DLH_X1 \CACHE_mem_reg[26][0]  ( .G(N617), .D(N644), .Q(\CACHE_mem[26][0] )
         );
  DLH_X1 \CACHE_mem_reg[27][1]  ( .G(N616), .D(N645), .Q(\CACHE_mem[27][1] )
         );
  DLH_X1 \CACHE_mem_reg[27][0]  ( .G(N616), .D(N644), .Q(\CACHE_mem[27][0] )
         );
  DLH_X1 \CACHE_mem_reg[28][1]  ( .G(N615), .D(N645), .Q(\CACHE_mem[28][1] )
         );
  DLH_X1 \CACHE_mem_reg[28][0]  ( .G(N615), .D(N644), .Q(\CACHE_mem[28][0] )
         );
  DLH_X1 \CACHE_mem_reg[29][1]  ( .G(N614), .D(N645), .Q(\CACHE_mem[29][1] )
         );
  DLH_X1 \CACHE_mem_reg[29][0]  ( .G(N614), .D(N644), .Q(\CACHE_mem[29][0] )
         );
  DLH_X1 \CACHE_mem_reg[30][1]  ( .G(N613), .D(N645), .Q(\CACHE_mem[30][1] )
         );
  DLH_X1 \CACHE_mem_reg[30][0]  ( .G(N613), .D(N644), .Q(\CACHE_mem[30][0] )
         );
  DLH_X1 \CACHE_mem_reg[31][1]  ( .G(N612), .D(N645), .Q(\CACHE_mem[31][1] )
         );
  DLH_X1 \CACHE_mem_reg[31][0]  ( .G(N612), .D(N644), .Q(\CACHE_mem[31][0] )
         );
  FA_X1 \add_65/U1_1  ( .A(N114), .B(IR_IN[1]), .CI(\add_59/n1 ), .CO(
        \add_65/carry[2] ), .S(N220) );
  FA_X1 \add_65/U1_2  ( .A(PC_IN[2]), .B(IR_IN[2]), .CI(\add_65/carry[2] ), 
        .CO(\add_65/carry[3] ), .S(N221) );
  FA_X1 \add_65/U1_3  ( .A(PC_IN[3]), .B(IR_IN[3]), .CI(\add_65/carry[3] ), 
        .CO(\add_65/carry[4] ), .S(N222) );
  FA_X1 \add_65/U1_4  ( .A(PC_IN[4]), .B(IR_IN[4]), .CI(\add_65/carry[4] ), 
        .CO(\add_65/carry[5] ), .S(N223) );
  FA_X1 \add_65/U1_5  ( .A(PC_IN[5]), .B(IR_IN[5]), .CI(\add_65/carry[5] ), 
        .CO(\add_65/carry[6] ), .S(N224) );
  FA_X1 \add_65/U1_6  ( .A(PC_IN[6]), .B(IR_IN[6]), .CI(\add_65/carry[6] ), 
        .CO(\add_65/carry[7] ), .S(N225) );
  FA_X1 \add_65/U1_7  ( .A(PC_IN[7]), .B(IR_IN[7]), .CI(\add_65/carry[7] ), 
        .CO(\add_65/carry[8] ), .S(N226) );
  FA_X1 \add_65/U1_8  ( .A(PC_IN[8]), .B(IR_IN[8]), .CI(\add_65/carry[8] ), 
        .CO(\add_65/carry[9] ), .S(N227) );
  FA_X1 \add_65/U1_9  ( .A(PC_IN[9]), .B(IR_IN[9]), .CI(\add_65/carry[9] ), 
        .CO(\add_65/carry[10] ), .S(N228) );
  FA_X1 \add_65/U1_10  ( .A(PC_IN[10]), .B(IR_IN[10]), .CI(\add_65/carry[10] ), 
        .CO(\add_65/carry[11] ), .S(N229) );
  FA_X1 \add_65/U1_11  ( .A(PC_IN[11]), .B(IR_IN[11]), .CI(\add_65/carry[11] ), 
        .CO(\add_65/carry[12] ), .S(N230) );
  FA_X1 \add_65/U1_12  ( .A(PC_IN[12]), .B(IR_IN[12]), .CI(\add_65/carry[12] ), 
        .CO(\add_65/carry[13] ), .S(N231) );
  FA_X1 \add_65/U1_13  ( .A(PC_IN[13]), .B(IR_IN[13]), .CI(\add_65/carry[13] ), 
        .CO(\add_65/carry[14] ), .S(N232) );
  FA_X1 \add_65/U1_14  ( .A(PC_IN[14]), .B(IR_IN[14]), .CI(\add_65/carry[14] ), 
        .CO(\add_65/carry[15] ), .S(N233) );
  FA_X1 \add_65/U1_15  ( .A(PC_IN[15]), .B(IR_IN[15]), .CI(\add_65/carry[15] ), 
        .CO(\add_65/carry[16] ), .S(N234) );
  FA_X1 \add_65/U1_16  ( .A(PC_IN[16]), .B(IR_IN[15]), .CI(\add_65/carry[16] ), 
        .CO(\add_65/carry[17] ), .S(N235) );
  FA_X1 \add_65/U1_17  ( .A(PC_IN[17]), .B(IR_IN[15]), .CI(\add_65/carry[17] ), 
        .CO(\add_65/carry[18] ), .S(N236) );
  FA_X1 \add_65/U1_18  ( .A(PC_IN[18]), .B(IR_IN[15]), .CI(\add_65/carry[18] ), 
        .CO(\add_65/carry[19] ), .S(N237) );
  FA_X1 \add_65/U1_19  ( .A(PC_IN[19]), .B(IR_IN[15]), .CI(\add_65/carry[19] ), 
        .CO(\add_65/carry[20] ), .S(N238) );
  FA_X1 \add_65/U1_20  ( .A(PC_IN[20]), .B(IR_IN[15]), .CI(\add_65/carry[20] ), 
        .CO(\add_65/carry[21] ), .S(N239) );
  FA_X1 \add_65/U1_21  ( .A(PC_IN[21]), .B(IR_IN[15]), .CI(\add_65/carry[21] ), 
        .CO(\add_65/carry[22] ), .S(N240) );
  FA_X1 \add_65/U1_22  ( .A(PC_IN[22]), .B(IR_IN[15]), .CI(\add_65/carry[22] ), 
        .CO(\add_65/carry[23] ), .S(N241) );
  FA_X1 \add_65/U1_23  ( .A(PC_IN[23]), .B(IR_IN[15]), .CI(\add_65/carry[23] ), 
        .CO(\add_65/carry[24] ), .S(N242) );
  FA_X1 \add_65/U1_24  ( .A(PC_IN[24]), .B(IR_IN[15]), .CI(\add_65/carry[24] ), 
        .CO(\add_65/carry[25] ), .S(N243) );
  FA_X1 \add_65/U1_25  ( .A(PC_IN[25]), .B(IR_IN[15]), .CI(\add_65/carry[25] ), 
        .CO(\add_65/carry[26] ), .S(N244) );
  FA_X1 \add_65/U1_26  ( .A(PC_IN[26]), .B(IR_IN[15]), .CI(\add_65/carry[26] ), 
        .CO(\add_65/carry[27] ), .S(N245) );
  FA_X1 \add_65/U1_27  ( .A(PC_IN[27]), .B(IR_IN[15]), .CI(\add_65/carry[27] ), 
        .CO(\add_65/carry[28] ), .S(N246) );
  FA_X1 \add_65/U1_28  ( .A(PC_IN[28]), .B(IR_IN[15]), .CI(\add_65/carry[28] ), 
        .CO(\add_65/carry[29] ), .S(N247) );
  FA_X1 \add_65/U1_29  ( .A(PC_IN[29]), .B(IR_IN[15]), .CI(\add_65/carry[29] ), 
        .CO(\add_65/carry[30] ), .S(N248) );
  FA_X1 \add_65/U1_30  ( .A(PC_IN[30]), .B(IR_IN[15]), .CI(\add_65/carry[30] ), 
        .CO(\add_65/carry[31] ), .S(N249) );
  FA_X1 \add_65/U1_31  ( .A(PC_IN[31]), .B(IR_IN[15]), .CI(\add_65/carry[31] ), 
        .S(N250) );
  FA_X1 \add_59/U1_1  ( .A(N114), .B(IR_IN[1]), .CI(\add_59/n1 ), .CO(
        \add_59/carry[2] ), .S(N82) );
  FA_X1 \add_59/U1_2  ( .A(PC_IN[2]), .B(IR_IN[2]), .CI(\add_59/carry[2] ), 
        .CO(\add_59/carry[3] ), .S(N83) );
  FA_X1 \add_59/U1_3  ( .A(PC_IN[3]), .B(IR_IN[3]), .CI(\add_59/carry[3] ), 
        .CO(\add_59/carry[4] ), .S(N84) );
  FA_X1 \add_59/U1_4  ( .A(PC_IN[4]), .B(IR_IN[4]), .CI(\add_59/carry[4] ), 
        .CO(\add_59/carry[5] ), .S(N85) );
  FA_X1 \add_59/U1_5  ( .A(PC_IN[5]), .B(IR_IN[5]), .CI(\add_59/carry[5] ), 
        .CO(\add_59/carry[6] ), .S(N86) );
  FA_X1 \add_59/U1_6  ( .A(PC_IN[6]), .B(IR_IN[6]), .CI(\add_59/carry[6] ), 
        .CO(\add_59/carry[7] ), .S(N87) );
  FA_X1 \add_59/U1_7  ( .A(PC_IN[7]), .B(IR_IN[7]), .CI(\add_59/carry[7] ), 
        .CO(\add_59/carry[8] ), .S(N88) );
  FA_X1 \add_59/U1_8  ( .A(PC_IN[8]), .B(IR_IN[8]), .CI(\add_59/carry[8] ), 
        .CO(\add_59/carry[9] ), .S(N89) );
  FA_X1 \add_59/U1_9  ( .A(PC_IN[9]), .B(IR_IN[9]), .CI(\add_59/carry[9] ), 
        .CO(\add_59/carry[10] ), .S(N90) );
  FA_X1 \add_59/U1_10  ( .A(PC_IN[10]), .B(IR_IN[10]), .CI(\add_59/carry[10] ), 
        .CO(\add_59/carry[11] ), .S(N91) );
  FA_X1 \add_59/U1_11  ( .A(PC_IN[11]), .B(IR_IN[11]), .CI(\add_59/carry[11] ), 
        .CO(\add_59/carry[12] ), .S(N92) );
  FA_X1 \add_59/U1_12  ( .A(PC_IN[12]), .B(IR_IN[12]), .CI(\add_59/carry[12] ), 
        .CO(\add_59/carry[13] ), .S(N93) );
  FA_X1 \add_59/U1_13  ( .A(PC_IN[13]), .B(IR_IN[13]), .CI(\add_59/carry[13] ), 
        .CO(\add_59/carry[14] ), .S(N94) );
  FA_X1 \add_59/U1_14  ( .A(PC_IN[14]), .B(IR_IN[14]), .CI(\add_59/carry[14] ), 
        .CO(\add_59/carry[15] ), .S(N95) );
  FA_X1 \add_59/U1_15  ( .A(PC_IN[15]), .B(IR_IN[15]), .CI(\add_59/carry[15] ), 
        .CO(\add_59/carry[16] ), .S(N96) );
  FA_X1 \add_59/U1_16  ( .A(PC_IN[16]), .B(IR_IN[16]), .CI(\add_59/carry[16] ), 
        .CO(\add_59/carry[17] ), .S(N97) );
  FA_X1 \add_59/U1_17  ( .A(PC_IN[17]), .B(IR_IN[17]), .CI(\add_59/carry[17] ), 
        .CO(\add_59/carry[18] ), .S(N98) );
  FA_X1 \add_59/U1_18  ( .A(PC_IN[18]), .B(IR_IN[18]), .CI(\add_59/carry[18] ), 
        .CO(\add_59/carry[19] ), .S(N99) );
  FA_X1 \add_59/U1_19  ( .A(PC_IN[19]), .B(IR_IN[19]), .CI(\add_59/carry[19] ), 
        .CO(\add_59/carry[20] ), .S(N100) );
  FA_X1 \add_59/U1_20  ( .A(PC_IN[20]), .B(IR_IN[20]), .CI(\add_59/carry[20] ), 
        .CO(\add_59/carry[21] ), .S(N101) );
  FA_X1 \add_59/U1_21  ( .A(PC_IN[21]), .B(IR_IN[21]), .CI(\add_59/carry[21] ), 
        .CO(\add_59/carry[22] ), .S(N102) );
  FA_X1 \add_59/U1_22  ( .A(PC_IN[22]), .B(IR_IN[22]), .CI(\add_59/carry[22] ), 
        .CO(\add_59/carry[23] ), .S(N103) );
  FA_X1 \add_59/U1_23  ( .A(PC_IN[23]), .B(IR_IN[23]), .CI(\add_59/carry[23] ), 
        .CO(\add_59/carry[24] ), .S(N104) );
  FA_X1 \add_59/U1_24  ( .A(PC_IN[24]), .B(IR_IN[24]), .CI(\add_59/carry[24] ), 
        .CO(\add_59/carry[25] ), .S(N105) );
  FA_X1 \add_59/U1_25  ( .A(PC_IN[25]), .B(IR_IN[25]), .CI(\add_59/carry[25] ), 
        .CO(\add_59/carry[26] ), .S(N106) );
  FA_X1 \add_59/U1_26  ( .A(PC_IN[26]), .B(IR_IN[25]), .CI(\add_59/carry[26] ), 
        .CO(\add_59/carry[27] ), .S(N107) );
  FA_X1 \add_59/U1_27  ( .A(PC_IN[27]), .B(IR_IN[25]), .CI(\add_59/carry[27] ), 
        .CO(\add_59/carry[28] ), .S(N108) );
  FA_X1 \add_59/U1_28  ( .A(PC_IN[28]), .B(IR_IN[25]), .CI(\add_59/carry[28] ), 
        .CO(\add_59/carry[29] ), .S(N109) );
  FA_X1 \add_59/U1_29  ( .A(PC_IN[29]), .B(IR_IN[25]), .CI(\add_59/carry[29] ), 
        .CO(\add_59/carry[30] ), .S(N110) );
  FA_X1 \add_59/U1_30  ( .A(PC_IN[30]), .B(IR_IN[25]), .CI(\add_59/carry[30] ), 
        .CO(\add_59/carry[31] ), .S(N111) );
  FA_X1 \add_59/U1_31  ( .A(PC_IN[31]), .B(IR_IN[25]), .CI(\add_59/carry[31] ), 
        .S(N112) );
  FA_X1 \add_53_aco/U1_1  ( .A(PC_FAIL[1]), .B(n6), .CI(\add_53_aco/n2 ), .CO(
        \add_53_aco/carry[2] ), .S(N47) );
  FA_X1 \add_53_aco/U1_2  ( .A(PC_FAIL[2]), .B(n8), .CI(\add_53_aco/carry[2] ), 
        .CO(\add_53_aco/carry[3] ), .S(N48) );
  FA_X1 \add_53_aco/U1_3  ( .A(PC_FAIL[3]), .B(n9), .CI(\add_53_aco/carry[3] ), 
        .CO(\add_53_aco/carry[4] ), .S(N49) );
  FA_X1 \add_53_aco/U1_4  ( .A(PC_FAIL[4]), .B(n10), .CI(\add_53_aco/carry[4] ), .CO(\add_53_aco/carry[5] ), .S(N50) );
  FA_X1 \add_53_aco/U1_5  ( .A(PC_FAIL[5]), .B(n7), .CI(\add_53_aco/carry[5] ), 
        .CO(\add_53_aco/carry[6] ), .S(N51) );
  FA_X1 \add_53_aco/U1_6  ( .A(PC_FAIL[6]), .B(n11), .CI(\add_53_aco/carry[6] ), .CO(\add_53_aco/carry[7] ), .S(N52) );
  FA_X1 \add_53_aco/U1_7  ( .A(PC_FAIL[7]), .B(n12), .CI(\add_53_aco/carry[7] ), .CO(\add_53_aco/carry[8] ), .S(N53) );
  FA_X1 \add_53_aco/U1_8  ( .A(PC_FAIL[8]), .B(n13), .CI(\add_53_aco/carry[8] ), .CO(\add_53_aco/carry[9] ), .S(N54) );
  FA_X1 \add_53_aco/U1_9  ( .A(PC_FAIL[9]), .B(n14), .CI(\add_53_aco/carry[9] ), .CO(\add_53_aco/carry[10] ), .S(N55) );
  FA_X1 \add_53_aco/U1_10  ( .A(PC_FAIL[10]), .B(n15), .CI(
        \add_53_aco/carry[10] ), .CO(\add_53_aco/carry[11] ), .S(N56) );
  FA_X1 \add_53_aco/U1_11  ( .A(PC_FAIL[11]), .B(n16), .CI(
        \add_53_aco/carry[11] ), .CO(\add_53_aco/carry[12] ), .S(N57) );
  FA_X1 \add_53_aco/U1_12  ( .A(PC_FAIL[12]), .B(n17), .CI(
        \add_53_aco/carry[12] ), .CO(\add_53_aco/carry[13] ), .S(N58) );
  FA_X1 \add_53_aco/U1_13  ( .A(PC_FAIL[13]), .B(n18), .CI(
        \add_53_aco/carry[13] ), .CO(\add_53_aco/carry[14] ), .S(N59) );
  FA_X1 \add_53_aco/U1_14  ( .A(PC_FAIL[14]), .B(n19), .CI(
        \add_53_aco/carry[14] ), .CO(\add_53_aco/carry[15] ), .S(N60) );
  FA_X1 \add_53_aco/U1_15  ( .A(PC_FAIL[15]), .B(n5), .CI(
        \add_53_aco/carry[15] ), .CO(\add_53_aco/carry[16] ), .S(N61) );
  FA_X1 \add_53_aco/U1_16  ( .A(PC_FAIL[16]), .B(n5), .CI(
        \add_53_aco/carry[16] ), .CO(\add_53_aco/carry[17] ), .S(N62) );
  FA_X1 \add_53_aco/U1_17  ( .A(PC_FAIL[17]), .B(n5), .CI(
        \add_53_aco/carry[17] ), .CO(\add_53_aco/carry[18] ), .S(N63) );
  FA_X1 \add_53_aco/U1_18  ( .A(PC_FAIL[18]), .B(n5), .CI(
        \add_53_aco/carry[18] ), .CO(\add_53_aco/carry[19] ), .S(N64) );
  FA_X1 \add_53_aco/U1_19  ( .A(PC_FAIL[19]), .B(n5), .CI(
        \add_53_aco/carry[19] ), .CO(\add_53_aco/carry[20] ), .S(N65) );
  FA_X1 \add_53_aco/U1_20  ( .A(PC_FAIL[20]), .B(n5), .CI(
        \add_53_aco/carry[20] ), .CO(\add_53_aco/carry[21] ), .S(N66) );
  FA_X1 \add_53_aco/U1_21  ( .A(PC_FAIL[21]), .B(n5), .CI(
        \add_53_aco/carry[21] ), .CO(\add_53_aco/carry[22] ), .S(N67) );
  FA_X1 \add_53_aco/U1_22  ( .A(PC_FAIL[22]), .B(n5), .CI(
        \add_53_aco/carry[22] ), .CO(\add_53_aco/carry[23] ), .S(N68) );
  FA_X1 \add_53_aco/U1_23  ( .A(PC_FAIL[23]), .B(n5), .CI(
        \add_53_aco/carry[23] ), .CO(\add_53_aco/carry[24] ), .S(N69) );
  FA_X1 \add_53_aco/U1_24  ( .A(PC_FAIL[24]), .B(n5), .CI(
        \add_53_aco/carry[24] ), .CO(\add_53_aco/carry[25] ), .S(N70) );
  FA_X1 \add_53_aco/U1_25  ( .A(PC_FAIL[25]), .B(n5), .CI(
        \add_53_aco/carry[25] ), .CO(\add_53_aco/carry[26] ), .S(N71) );
  FA_X1 \add_53_aco/U1_26  ( .A(PC_FAIL[26]), .B(n5), .CI(
        \add_53_aco/carry[26] ), .CO(\add_53_aco/carry[27] ), .S(N72) );
  FA_X1 \add_53_aco/U1_27  ( .A(PC_FAIL[27]), .B(n5), .CI(
        \add_53_aco/carry[27] ), .CO(\add_53_aco/carry[28] ), .S(N73) );
  FA_X1 \add_53_aco/U1_28  ( .A(PC_FAIL[28]), .B(n5), .CI(
        \add_53_aco/carry[28] ), .CO(\add_53_aco/carry[29] ), .S(N74) );
  FA_X1 \add_53_aco/U1_29  ( .A(PC_FAIL[29]), .B(n5), .CI(
        \add_53_aco/carry[29] ), .CO(\add_53_aco/carry[30] ), .S(N75) );
  FA_X1 \add_53_aco/U1_30  ( .A(PC_FAIL[30]), .B(n5), .CI(
        \add_53_aco/carry[30] ), .CO(\add_53_aco/carry[31] ), .S(N76) );
  FA_X1 \add_53_aco/U1_31  ( .A(PC_FAIL[31]), .B(n5), .CI(
        \add_53_aco/carry[31] ), .S(N77) );
  NAND2_X1 U3 ( .A1(n5320), .A2(n5455), .ZN(N323) );
  AOI21_X1 U4 ( .B1(n5451), .B2(RIGHT_PRE), .A(n5548), .ZN(n5400) );
  INV_X1 U5 ( .A(n5516), .ZN(n5319) );
  NAND2_X1 U6 ( .A1(n5515), .A2(n5319), .ZN(n5321) );
  NOR2_X2 U7 ( .A1(n5325), .A2(n5454), .ZN(N645) );
  INV_X2 U8 ( .A(n5321), .ZN(n5320) );
  NOR2_X2 U9 ( .A1(n5465), .A2(n5451), .ZN(N644) );
  INV_X2 U10 ( .A(n5465), .ZN(n5548) );
  NOR3_X2 U11 ( .A1(n5373), .A2(n5376), .A3(n5375), .ZN(n5429) );
  AOI211_X4 U12 ( .C1(n5449), .C2(n5448), .A(n5447), .B(n5446), .ZN(n5467) );
  BUF_X1 U13 ( .A(N356), .Z(n5323) );
  INV_X1 U14 ( .A(n5429), .ZN(n5405) );
  OAI221_X1 U15 ( .B1(n5324), .B2(n5515), .C1(n5324), .C2(n5455), .A(n5465), 
        .ZN(SEL) );
  BUF_X1 U16 ( .A(n5547), .Z(n5322) );
  NOR2_X1 U17 ( .A1(n5516), .A2(n5515), .ZN(n5547) );
  INV_X1 U18 ( .A(PC_FAIL[2]), .ZN(n5375) );
  INV_X1 U19 ( .A(PC_FAIL[5]), .ZN(n5430) );
  INV_X1 U20 ( .A(PC_FAIL[3]), .ZN(n5376) );
  INV_X1 U21 ( .A(RST), .ZN(n5324) );
  INV_X1 U22 ( .A(RST), .ZN(n5325) );
  INV_X1 U23 ( .A(IR_IN[28]), .ZN(n5326) );
  INV_X1 U24 ( .A(n5457), .ZN(n5461) );
  AND2_X2 U25 ( .A1(n5467), .A2(IR_FAIL[15]), .ZN(n5) );
  INV_X1 U26 ( .A(PC_FAIL[6]), .ZN(n5431) );
  NOR2_X1 U27 ( .A1(PC_FAIL[4]), .A2(n5374), .ZN(n5436) );
  NOR3_X1 U28 ( .A1(IR_IN[29]), .A2(IR_IN[30]), .A3(IR_IN[31]), .ZN(n5365) );
  NAND3_X1 U29 ( .A1(n5365), .A2(IR_IN[27]), .A3(n5326), .ZN(n5515) );
  INV_X1 U30 ( .A(WRONG_PRE), .ZN(n5453) );
  NAND2_X1 U31 ( .A1(RST), .A2(n5453), .ZN(n5516) );
  NAND2_X1 U32 ( .A1(PC_IN[3]), .A2(PC_IN[2]), .ZN(n5457) );
  INV_X1 U33 ( .A(PC_IN[4]), .ZN(n5456) );
  INV_X1 U34 ( .A(PC_IN[5]), .ZN(n5368) );
  NOR2_X1 U35 ( .A1(n5456), .A2(n5368), .ZN(n5343) );
  NAND2_X1 U36 ( .A1(n5461), .A2(n5343), .ZN(n5460) );
  INV_X1 U37 ( .A(n5460), .ZN(n5366) );
  NAND2_X1 U38 ( .A1(n5366), .A2(PC_IN[6]), .ZN(n5514) );
  INV_X1 U39 ( .A(n5514), .ZN(n5458) );
  AOI21_X1 U40 ( .B1(\CACHE_mem[31][1] ), .B2(n5458), .A(IR_IN[27]), .ZN(n5364) );
  NOR2_X1 U41 ( .A1(PC_IN[5]), .A2(n5456), .ZN(n5351) );
  AND2_X1 U42 ( .A1(\CACHE_mem[21][1] ), .A2(n5351), .ZN(n5327) );
  INV_X1 U43 ( .A(PC_IN[6]), .ZN(n5459) );
  AOI211_X1 U44 ( .C1(n5343), .C2(\CACHE_mem[29][1] ), .A(n5327), .B(n5459), 
        .ZN(n5334) );
  NOR2_X1 U45 ( .A1(PC_IN[4]), .A2(n5368), .ZN(n5350) );
  NOR2_X1 U46 ( .A1(PC_IN[4]), .A2(PC_IN[5]), .ZN(n5352) );
  AOI22_X1 U47 ( .A1(\CACHE_mem[25][1] ), .A2(n5350), .B1(\CACHE_mem[17][1] ), 
        .B2(n5352), .ZN(n5333) );
  INV_X1 U48 ( .A(\CACHE_mem[5][1] ), .ZN(n5330) );
  INV_X1 U49 ( .A(n5351), .ZN(n5329) );
  AOI22_X1 U50 ( .A1(n5343), .A2(\CACHE_mem[13][1] ), .B1(\CACHE_mem[9][1] ), 
        .B2(n5350), .ZN(n5328) );
  OAI211_X1 U51 ( .C1(n5330), .C2(n5329), .A(n5328), .B(n5459), .ZN(n5331) );
  AOI21_X1 U52 ( .B1(\CACHE_mem[1][1] ), .B2(n5352), .A(n5331), .ZN(n5332) );
  AOI211_X1 U53 ( .C1(n5334), .C2(n5333), .A(PC_IN[3]), .B(n5332), .ZN(n5362)
         );
  AOI22_X1 U54 ( .A1(n5343), .A2(\CACHE_mem[14][1] ), .B1(\CACHE_mem[10][1] ), 
        .B2(n5350), .ZN(n5336) );
  AOI22_X1 U55 ( .A1(\CACHE_mem[2][1] ), .A2(n5352), .B1(\CACHE_mem[6][1] ), 
        .B2(n5351), .ZN(n5335) );
  INV_X1 U56 ( .A(PC_IN[3]), .ZN(n5463) );
  AOI21_X1 U57 ( .B1(n5336), .B2(n5335), .A(n5463), .ZN(n5340) );
  AOI22_X1 U58 ( .A1(n5343), .A2(\CACHE_mem[12][1] ), .B1(\CACHE_mem[8][1] ), 
        .B2(n5350), .ZN(n5338) );
  AOI22_X1 U59 ( .A1(\CACHE_mem[0][1] ), .A2(n5352), .B1(\CACHE_mem[4][1] ), 
        .B2(n5351), .ZN(n5337) );
  AOI21_X1 U60 ( .B1(n5338), .B2(n5337), .A(PC_IN[3]), .ZN(n5339) );
  NOR2_X1 U61 ( .A1(n5340), .A2(n5339), .ZN(n5349) );
  AOI22_X1 U62 ( .A1(n5343), .A2(\CACHE_mem[30][1] ), .B1(\CACHE_mem[26][1] ), 
        .B2(n5350), .ZN(n5342) );
  AOI22_X1 U63 ( .A1(\CACHE_mem[18][1] ), .A2(n5352), .B1(\CACHE_mem[22][1] ), 
        .B2(n5351), .ZN(n5341) );
  AOI21_X1 U64 ( .B1(n5342), .B2(n5341), .A(n5463), .ZN(n5347) );
  AOI22_X1 U65 ( .A1(n5343), .A2(\CACHE_mem[28][1] ), .B1(\CACHE_mem[24][1] ), 
        .B2(n5350), .ZN(n5345) );
  AOI22_X1 U66 ( .A1(\CACHE_mem[20][1] ), .A2(n5351), .B1(\CACHE_mem[16][1] ), 
        .B2(n5352), .ZN(n5344) );
  AOI21_X1 U67 ( .B1(n5345), .B2(n5344), .A(PC_IN[3]), .ZN(n5346) );
  OAI21_X1 U68 ( .B1(n5347), .B2(n5346), .A(PC_IN[6]), .ZN(n5348) );
  OAI21_X1 U69 ( .B1(PC_IN[6]), .B2(n5349), .A(n5348), .ZN(n5361) );
  INV_X1 U70 ( .A(PC_IN[2]), .ZN(n5462) );
  AOI21_X1 U71 ( .B1(\CACHE_mem[23][1] ), .B2(n5351), .A(n5459), .ZN(n5359) );
  AOI22_X1 U72 ( .A1(\CACHE_mem[27][1] ), .A2(n5350), .B1(\CACHE_mem[19][1] ), 
        .B2(n5352), .ZN(n5358) );
  INV_X1 U73 ( .A(\CACHE_mem[11][1] ), .ZN(n5355) );
  INV_X1 U74 ( .A(n5350), .ZN(n5354) );
  AOI22_X1 U75 ( .A1(\CACHE_mem[3][1] ), .A2(n5352), .B1(\CACHE_mem[7][1] ), 
        .B2(n5351), .ZN(n5353) );
  OAI211_X1 U76 ( .C1(n5355), .C2(n5354), .A(n5353), .B(n5459), .ZN(n5356) );
  AOI22_X1 U77 ( .A1(n5461), .A2(n5356), .B1(n5366), .B2(\CACHE_mem[15][1] ), 
        .ZN(n5357) );
  AOI21_X1 U78 ( .B1(n5359), .B2(n5358), .A(n5357), .ZN(n5360) );
  AOI221_X1 U79 ( .B1(n5362), .B2(PC_IN[2]), .C1(n5361), .C2(n5462), .A(n5360), 
        .ZN(n5363) );
  NAND4_X1 U80 ( .A1(n5365), .A2(IR_IN[28]), .A3(n5364), .A4(n5363), .ZN(n5455) );
  OAI21_X1 U81 ( .B1(WRONG_PRE), .B2(n5515), .A(RST), .ZN(N356) );
  AND2_X1 U82 ( .A1(RST), .A2(N113), .ZN(N357) );
  AND2_X1 U83 ( .A1(RST), .A2(N114), .ZN(N358) );
  NAND2_X1 U84 ( .A1(n5461), .A2(PC_IN[4]), .ZN(n5367) );
  AOI211_X1 U85 ( .C1(n5368), .C2(n5367), .A(n5366), .B(n5325), .ZN(N362) );
  INV_X1 U86 ( .A(PC_IN[7]), .ZN(n5513) );
  NOR2_X1 U87 ( .A1(n5514), .A2(n5513), .ZN(n5512) );
  NAND2_X1 U88 ( .A1(n5512), .A2(PC_IN[8]), .ZN(n5511) );
  INV_X1 U89 ( .A(PC_IN[9]), .ZN(n5510) );
  NOR2_X1 U90 ( .A1(n5511), .A2(n5510), .ZN(n5509) );
  NAND2_X1 U91 ( .A1(n5509), .A2(PC_IN[10]), .ZN(n5508) );
  INV_X1 U92 ( .A(PC_IN[11]), .ZN(n5507) );
  NOR2_X1 U93 ( .A1(n5508), .A2(n5507), .ZN(n5506) );
  NAND2_X1 U94 ( .A1(n5506), .A2(PC_IN[12]), .ZN(n5505) );
  INV_X1 U95 ( .A(PC_IN[13]), .ZN(n5504) );
  NOR2_X1 U96 ( .A1(n5505), .A2(n5504), .ZN(n5503) );
  NAND2_X1 U97 ( .A1(n5503), .A2(PC_IN[14]), .ZN(n5502) );
  INV_X1 U98 ( .A(PC_IN[15]), .ZN(n5501) );
  NOR2_X1 U99 ( .A1(n5502), .A2(n5501), .ZN(n5500) );
  NAND2_X1 U100 ( .A1(n5500), .A2(PC_IN[16]), .ZN(n5499) );
  INV_X1 U101 ( .A(PC_IN[17]), .ZN(n5498) );
  NOR2_X1 U102 ( .A1(n5499), .A2(n5498), .ZN(n5497) );
  NAND2_X1 U103 ( .A1(n5497), .A2(PC_IN[18]), .ZN(n5496) );
  INV_X1 U104 ( .A(PC_IN[19]), .ZN(n5495) );
  NOR2_X1 U105 ( .A1(n5496), .A2(n5495), .ZN(n5494) );
  NAND2_X1 U106 ( .A1(n5494), .A2(PC_IN[20]), .ZN(n5493) );
  INV_X1 U107 ( .A(PC_IN[21]), .ZN(n5492) );
  NOR2_X1 U108 ( .A1(n5493), .A2(n5492), .ZN(n5491) );
  NAND2_X1 U109 ( .A1(n5491), .A2(PC_IN[22]), .ZN(n5490) );
  INV_X1 U110 ( .A(PC_IN[23]), .ZN(n5489) );
  NOR2_X1 U111 ( .A1(n5490), .A2(n5489), .ZN(n5488) );
  NAND2_X1 U112 ( .A1(n5488), .A2(PC_IN[24]), .ZN(n5487) );
  INV_X1 U113 ( .A(PC_IN[25]), .ZN(n5486) );
  NOR2_X1 U114 ( .A1(n5487), .A2(n5486), .ZN(n5485) );
  NAND2_X1 U115 ( .A1(n5485), .A2(PC_IN[26]), .ZN(n5484) );
  INV_X1 U116 ( .A(PC_IN[27]), .ZN(n5483) );
  NOR2_X1 U117 ( .A1(n5484), .A2(n5483), .ZN(n5482) );
  NAND2_X1 U118 ( .A1(n5482), .A2(PC_IN[28]), .ZN(n5481) );
  INV_X1 U119 ( .A(PC_IN[29]), .ZN(n5480) );
  NOR2_X1 U120 ( .A1(n5481), .A2(n5480), .ZN(n5479) );
  INV_X1 U121 ( .A(n5479), .ZN(n5370) );
  INV_X1 U122 ( .A(PC_IN[30]), .ZN(n5369) );
  NOR2_X1 U123 ( .A1(n5370), .A2(n5369), .ZN(n5372) );
  AOI211_X1 U124 ( .C1(n5370), .C2(n5369), .A(n5372), .B(n5324), .ZN(N387) );
  OAI21_X1 U125 ( .B1(PC_IN[31]), .B2(n5372), .A(RST), .ZN(n5371) );
  AOI21_X1 U126 ( .B1(PC_IN[31]), .B2(n5372), .A(n5371), .ZN(N388) );
  INV_X1 U127 ( .A(PC_FAIL[4]), .ZN(n5373) );
  NAND3_X1 U128 ( .A1(n5373), .A2(n5376), .A3(n5375), .ZN(n5413) );
  INV_X1 U129 ( .A(n5413), .ZN(n5434) );
  NAND3_X1 U130 ( .A1(n5373), .A2(n5376), .A3(PC_FAIL[2]), .ZN(n5411) );
  INV_X1 U131 ( .A(n5411), .ZN(n5428) );
  AOI22_X1 U132 ( .A1(n5434), .A2(\CACHE_mem[8][0] ), .B1(n5428), .B2(
        \CACHE_mem[9][0] ), .ZN(n5380) );
  NAND3_X1 U133 ( .A1(n5373), .A2(n5375), .A3(PC_FAIL[3]), .ZN(n5410) );
  INV_X1 U134 ( .A(n5410), .ZN(n5433) );
  NAND2_X1 U135 ( .A1(PC_FAIL[3]), .A2(PC_FAIL[2]), .ZN(n5374) );
  AOI22_X1 U136 ( .A1(n5433), .A2(\CACHE_mem[10][0] ), .B1(n5436), .B2(
        \CACHE_mem[11][0] ), .ZN(n5379) );
  NAND3_X1 U137 ( .A1(n5376), .A2(n5375), .A3(PC_FAIL[4]), .ZN(n5408) );
  INV_X1 U138 ( .A(n5408), .ZN(n5435) );
  NAND3_X1 U139 ( .A1(n5375), .A2(PC_FAIL[3]), .A3(PC_FAIL[4]), .ZN(n5406) );
  INV_X1 U140 ( .A(n5406), .ZN(n5438) );
  AOI22_X1 U141 ( .A1(n5435), .A2(\CACHE_mem[12][0] ), .B1(n5438), .B2(
        \CACHE_mem[14][0] ), .ZN(n5378) );
  NAND3_X1 U142 ( .A1(n5376), .A2(PC_FAIL[4]), .A3(PC_FAIL[2]), .ZN(n5407) );
  INV_X1 U143 ( .A(n5407), .ZN(n5437) );
  AOI22_X1 U144 ( .A1(n5429), .A2(\CACHE_mem[15][0] ), .B1(n5437), .B2(
        \CACHE_mem[13][0] ), .ZN(n5377) );
  NAND4_X1 U145 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n5386)
         );
  AOI22_X1 U146 ( .A1(n5428), .A2(\CACHE_mem[1][0] ), .B1(n5433), .B2(
        \CACHE_mem[2][0] ), .ZN(n5384) );
  AOI22_X1 U147 ( .A1(n5436), .A2(\CACHE_mem[3][0] ), .B1(n5438), .B2(
        \CACHE_mem[6][0] ), .ZN(n5383) );
  AOI22_X1 U148 ( .A1(n5429), .A2(\CACHE_mem[7][0] ), .B1(n5437), .B2(
        \CACHE_mem[5][0] ), .ZN(n5382) );
  AOI22_X1 U149 ( .A1(n5434), .A2(\CACHE_mem[0][0] ), .B1(n5435), .B2(
        \CACHE_mem[4][0] ), .ZN(n5381) );
  NAND4_X1 U150 ( .A1(n5384), .A2(n5383), .A3(n5382), .A4(n5381), .ZN(n5385)
         );
  AOI22_X1 U151 ( .A1(PC_FAIL[5]), .A2(n5386), .B1(n5385), .B2(n5430), .ZN(
        n5398) );
  AOI22_X1 U152 ( .A1(n5428), .A2(\CACHE_mem[17][0] ), .B1(n5433), .B2(
        \CACHE_mem[18][0] ), .ZN(n5390) );
  AOI22_X1 U153 ( .A1(n5436), .A2(\CACHE_mem[19][0] ), .B1(n5438), .B2(
        \CACHE_mem[22][0] ), .ZN(n5389) );
  AOI22_X1 U154 ( .A1(n5429), .A2(\CACHE_mem[23][0] ), .B1(n5437), .B2(
        \CACHE_mem[21][0] ), .ZN(n5388) );
  AOI22_X1 U155 ( .A1(n5434), .A2(\CACHE_mem[16][0] ), .B1(n5435), .B2(
        \CACHE_mem[20][0] ), .ZN(n5387) );
  NAND4_X1 U156 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n5396)
         );
  AOI22_X1 U157 ( .A1(n5434), .A2(\CACHE_mem[24][0] ), .B1(n5428), .B2(
        \CACHE_mem[25][0] ), .ZN(n5394) );
  AOI22_X1 U158 ( .A1(n5433), .A2(\CACHE_mem[26][0] ), .B1(n5436), .B2(
        \CACHE_mem[27][0] ), .ZN(n5393) );
  AOI22_X1 U159 ( .A1(n5435), .A2(\CACHE_mem[28][0] ), .B1(n5438), .B2(
        \CACHE_mem[30][0] ), .ZN(n5392) );
  AOI22_X1 U160 ( .A1(n5429), .A2(\CACHE_mem[31][0] ), .B1(n5437), .B2(
        \CACHE_mem[29][0] ), .ZN(n5391) );
  NAND4_X1 U161 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n5395)
         );
  OAI221_X1 U162 ( .B1(PC_FAIL[5]), .B2(n5396), .C1(n5430), .C2(n5395), .A(
        PC_FAIL[6]), .ZN(n5397) );
  OAI21_X1 U163 ( .B1(PC_FAIL[6]), .B2(n5398), .A(n5397), .ZN(n5451) );
  NAND2_X1 U164 ( .A1(RST), .A2(WRONG_PRE), .ZN(n5465) );
  NOR2_X1 U165 ( .A1(n5400), .A2(n5430), .ZN(n5402) );
  NAND2_X1 U166 ( .A1(PC_FAIL[6]), .A2(n5402), .ZN(n5399) );
  OAI21_X1 U167 ( .B1(n5405), .B2(n5399), .A(RST), .ZN(N612) );
  OAI21_X1 U168 ( .B1(n5406), .B2(n5399), .A(RST), .ZN(N613) );
  OAI21_X1 U169 ( .B1(n5407), .B2(n5399), .A(RST), .ZN(N614) );
  OAI21_X1 U170 ( .B1(n5408), .B2(n5399), .A(RST), .ZN(N615) );
  INV_X1 U171 ( .A(n5436), .ZN(n5409) );
  OAI21_X1 U172 ( .B1(n5409), .B2(n5399), .A(RST), .ZN(N616) );
  OAI21_X1 U173 ( .B1(n5410), .B2(n5399), .A(RST), .ZN(N617) );
  OAI21_X1 U174 ( .B1(n5411), .B2(n5399), .A(RST), .ZN(N618) );
  OAI21_X1 U175 ( .B1(n5413), .B2(n5399), .A(RST), .ZN(N619) );
  NOR2_X1 U176 ( .A1(PC_FAIL[5]), .A2(n5400), .ZN(n5404) );
  NAND2_X1 U177 ( .A1(PC_FAIL[6]), .A2(n5404), .ZN(n5401) );
  OAI21_X1 U178 ( .B1(n5405), .B2(n5401), .A(RST), .ZN(N620) );
  OAI21_X1 U179 ( .B1(n5406), .B2(n5401), .A(RST), .ZN(N621) );
  OAI21_X1 U180 ( .B1(n5407), .B2(n5401), .A(RST), .ZN(N622) );
  OAI21_X1 U181 ( .B1(n5408), .B2(n5401), .A(RST), .ZN(N623) );
  OAI21_X1 U182 ( .B1(n5409), .B2(n5401), .A(RST), .ZN(N624) );
  OAI21_X1 U183 ( .B1(n5410), .B2(n5401), .A(RST), .ZN(N625) );
  OAI21_X1 U184 ( .B1(n5411), .B2(n5401), .A(RST), .ZN(N626) );
  OAI21_X1 U185 ( .B1(n5413), .B2(n5401), .A(RST), .ZN(N627) );
  NAND2_X1 U186 ( .A1(n5402), .A2(n5431), .ZN(n5403) );
  OAI21_X1 U187 ( .B1(n5405), .B2(n5403), .A(RST), .ZN(N628) );
  OAI21_X1 U188 ( .B1(n5406), .B2(n5403), .A(RST), .ZN(N629) );
  OAI21_X1 U189 ( .B1(n5407), .B2(n5403), .A(RST), .ZN(N630) );
  OAI21_X1 U190 ( .B1(n5408), .B2(n5403), .A(RST), .ZN(N631) );
  OAI21_X1 U191 ( .B1(n5409), .B2(n5403), .A(RST), .ZN(N632) );
  OAI21_X1 U192 ( .B1(n5410), .B2(n5403), .A(RST), .ZN(N633) );
  OAI21_X1 U193 ( .B1(n5411), .B2(n5403), .A(RST), .ZN(N634) );
  OAI21_X1 U194 ( .B1(n5413), .B2(n5403), .A(RST), .ZN(N635) );
  NAND2_X1 U195 ( .A1(n5404), .A2(n5431), .ZN(n5412) );
  OAI21_X1 U196 ( .B1(n5405), .B2(n5412), .A(RST), .ZN(N636) );
  OAI21_X1 U197 ( .B1(n5406), .B2(n5412), .A(RST), .ZN(N637) );
  OAI21_X1 U198 ( .B1(n5407), .B2(n5412), .A(RST), .ZN(N638) );
  OAI21_X1 U199 ( .B1(n5408), .B2(n5412), .A(RST), .ZN(N639) );
  OAI21_X1 U200 ( .B1(n5409), .B2(n5412), .A(RST), .ZN(N640) );
  OAI21_X1 U201 ( .B1(n5410), .B2(n5412), .A(RST), .ZN(N641) );
  OAI21_X1 U202 ( .B1(n5411), .B2(n5412), .A(RST), .ZN(N642) );
  OAI21_X1 U203 ( .B1(n5413), .B2(n5412), .A(RST), .ZN(N643) );
  AOI22_X1 U204 ( .A1(n5428), .A2(\CACHE_mem[9][1] ), .B1(n5436), .B2(
        \CACHE_mem[11][1] ), .ZN(n5449) );
  NOR2_X1 U205 ( .A1(PC_FAIL[6]), .A2(n5430), .ZN(n5417) );
  AOI22_X1 U206 ( .A1(n5438), .A2(\CACHE_mem[14][1] ), .B1(n5437), .B2(
        \CACHE_mem[13][1] ), .ZN(n5416) );
  AOI22_X1 U207 ( .A1(n5429), .A2(\CACHE_mem[15][1] ), .B1(n5434), .B2(
        \CACHE_mem[8][1] ), .ZN(n5415) );
  AOI22_X1 U208 ( .A1(n5433), .A2(\CACHE_mem[10][1] ), .B1(n5435), .B2(
        \CACHE_mem[12][1] ), .ZN(n5414) );
  AND4_X1 U209 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n5448) );
  AOI211_X1 U210 ( .C1(n5438), .C2(\CACHE_mem[30][1] ), .A(n5430), .B(n5431), 
        .ZN(n5418) );
  INV_X1 U211 ( .A(n5418), .ZN(n5423) );
  AOI22_X1 U212 ( .A1(n5434), .A2(\CACHE_mem[24][1] ), .B1(n5435), .B2(
        \CACHE_mem[28][1] ), .ZN(n5421) );
  AOI22_X1 U213 ( .A1(n5428), .A2(\CACHE_mem[25][1] ), .B1(n5437), .B2(
        \CACHE_mem[29][1] ), .ZN(n5420) );
  AOI22_X1 U214 ( .A1(n5429), .A2(\CACHE_mem[31][1] ), .B1(n5436), .B2(
        \CACHE_mem[27][1] ), .ZN(n5419) );
  NAND3_X1 U215 ( .A1(n5421), .A2(n5420), .A3(n5419), .ZN(n5422) );
  AOI211_X1 U216 ( .C1(n5433), .C2(\CACHE_mem[26][1] ), .A(n5423), .B(n5422), 
        .ZN(n5447) );
  AOI22_X1 U217 ( .A1(n5434), .A2(\CACHE_mem[16][1] ), .B1(n5436), .B2(
        \CACHE_mem[19][1] ), .ZN(n5424) );
  NAND3_X1 U218 ( .A1(PC_FAIL[6]), .A2(n5424), .A3(n5430), .ZN(n5445) );
  AOI22_X1 U219 ( .A1(n5428), .A2(\CACHE_mem[17][1] ), .B1(n5433), .B2(
        \CACHE_mem[18][1] ), .ZN(n5427) );
  AOI22_X1 U220 ( .A1(n5435), .A2(\CACHE_mem[20][1] ), .B1(n5438), .B2(
        \CACHE_mem[22][1] ), .ZN(n5426) );
  AOI22_X1 U221 ( .A1(n5429), .A2(\CACHE_mem[23][1] ), .B1(n5437), .B2(
        \CACHE_mem[21][1] ), .ZN(n5425) );
  NAND3_X1 U222 ( .A1(n5427), .A2(n5426), .A3(n5425), .ZN(n5444) );
  AOI22_X1 U223 ( .A1(n5429), .A2(\CACHE_mem[7][1] ), .B1(n5428), .B2(
        \CACHE_mem[1][1] ), .ZN(n5432) );
  NAND3_X1 U224 ( .A1(n5432), .A2(n5431), .A3(n5430), .ZN(n5443) );
  AOI22_X1 U225 ( .A1(n5434), .A2(\CACHE_mem[0][1] ), .B1(n5433), .B2(
        \CACHE_mem[2][1] ), .ZN(n5441) );
  AOI22_X1 U226 ( .A1(n5436), .A2(\CACHE_mem[3][1] ), .B1(n5435), .B2(
        \CACHE_mem[4][1] ), .ZN(n5440) );
  AOI22_X1 U227 ( .A1(n5438), .A2(\CACHE_mem[6][1] ), .B1(n5437), .B2(
        \CACHE_mem[5][1] ), .ZN(n5439) );
  NAND3_X1 U228 ( .A1(n5441), .A2(n5440), .A3(n5439), .ZN(n5442) );
  OAI22_X1 U229 ( .A1(n5445), .A2(n5444), .B1(n5443), .B2(n5442), .ZN(n5446)
         );
  NOR2_X1 U230 ( .A1(n5467), .A2(n5453), .ZN(n5450) );
  XNOR2_X1 U231 ( .A(n5451), .B(n5450), .ZN(n5452) );
  AOI21_X1 U232 ( .B1(n5467), .B2(n5453), .A(n5452), .ZN(n5454) );
  NOR2_X1 U233 ( .A1(n5455), .A2(n5321), .ZN(TAKEN) );
  AND3_X1 U234 ( .A1(n5467), .A2(IR_FAIL[0]), .A3(PC_FAIL[0]), .ZN(
        \add_53_aco/n2 ) );
  AND2_X1 U235 ( .A1(N113), .A2(IR_IN[0]), .ZN(\add_59/n1 ) );
  AND2_X1 U236 ( .A1(n5467), .A2(IR_FAIL[4]), .ZN(n10) );
  AND2_X1 U237 ( .A1(n5467), .A2(IR_FAIL[6]), .ZN(n11) );
  AND2_X1 U238 ( .A1(n5467), .A2(IR_FAIL[7]), .ZN(n12) );
  AND2_X1 U239 ( .A1(n5467), .A2(IR_FAIL[8]), .ZN(n13) );
  AND2_X1 U240 ( .A1(n5467), .A2(IR_FAIL[9]), .ZN(n14) );
  AND2_X1 U241 ( .A1(n5467), .A2(IR_FAIL[10]), .ZN(n15) );
  AND2_X1 U242 ( .A1(n5467), .A2(IR_FAIL[11]), .ZN(n16) );
  AND2_X1 U243 ( .A1(n5467), .A2(IR_FAIL[12]), .ZN(n17) );
  AND2_X1 U244 ( .A1(n5467), .A2(IR_FAIL[13]), .ZN(n18) );
  AND2_X1 U245 ( .A1(n5467), .A2(IR_FAIL[14]), .ZN(n19) );
  AOI221_X1 U246 ( .B1(n5461), .B2(PC_IN[4]), .C1(n5457), .C2(n5456), .A(n5325), .ZN(n286) );
  AOI211_X1 U247 ( .C1(n5460), .C2(n5459), .A(n5458), .B(n5324), .ZN(n291) );
  AOI211_X1 U248 ( .C1(n5463), .C2(n5462), .A(n5461), .B(n5324), .ZN(n59) );
  AND2_X1 U249 ( .A1(n5467), .A2(IR_FAIL[1]), .ZN(n6) );
  NOR2_X1 U250 ( .A1(N113), .A2(IR_IN[0]), .ZN(n5466) );
  AOI21_X1 U251 ( .B1(IR_FAIL[0]), .B2(n5467), .A(PC_FAIL[0]), .ZN(n5464) );
  OAI33_X1 U252 ( .A1(n5516), .A2(\add_59/n1 ), .A3(n5466), .B1(n5465), .B2(
        n5464), .B3(\add_53_aco/n2 ), .ZN(n60) );
  NOR2_X1 U253 ( .A1(PC_IN[2]), .A2(n5324), .ZN(n62) );
  AND2_X1 U254 ( .A1(n5467), .A2(IR_FAIL[5]), .ZN(n7) );
  AND2_X1 U255 ( .A1(n5467), .A2(IR_FAIL[2]), .ZN(n8) );
  AND2_X1 U256 ( .A1(n5467), .A2(IR_FAIL[3]), .ZN(n9) );
  OAI211_X1 U257 ( .C1(n5491), .C2(PC_IN[22]), .A(n5490), .B(RST), .ZN(n5468)
         );
  INV_X1 U258 ( .A(n5468), .ZN(n292) );
  OAI211_X1 U259 ( .C1(n5494), .C2(PC_IN[20]), .A(n5493), .B(RST), .ZN(n5469)
         );
  INV_X1 U260 ( .A(n5469), .ZN(n290) );
  OAI211_X1 U261 ( .C1(n5500), .C2(PC_IN[16]), .A(n5499), .B(RST), .ZN(n5470)
         );
  INV_X1 U262 ( .A(n5470), .ZN(n289) );
  OAI211_X1 U263 ( .C1(n5485), .C2(PC_IN[26]), .A(n5484), .B(RST), .ZN(n5471)
         );
  INV_X1 U264 ( .A(n5471), .ZN(n288) );
  OAI211_X1 U265 ( .C1(n5488), .C2(PC_IN[24]), .A(n5487), .B(RST), .ZN(n5472)
         );
  INV_X1 U266 ( .A(n5472), .ZN(n287) );
  OAI211_X1 U267 ( .C1(n5509), .C2(PC_IN[10]), .A(n5508), .B(RST), .ZN(n5473)
         );
  INV_X1 U268 ( .A(n5473), .ZN(n285) );
  OAI211_X1 U269 ( .C1(n5506), .C2(PC_IN[12]), .A(n5505), .B(RST), .ZN(n5474)
         );
  INV_X1 U270 ( .A(n5474), .ZN(n284) );
  OAI211_X1 U271 ( .C1(n5497), .C2(PC_IN[18]), .A(n5496), .B(RST), .ZN(n5475)
         );
  INV_X1 U272 ( .A(n5475), .ZN(n283) );
  OAI211_X1 U273 ( .C1(n5482), .C2(PC_IN[28]), .A(n5481), .B(RST), .ZN(n5476)
         );
  INV_X1 U274 ( .A(n5476), .ZN(n282) );
  OAI211_X1 U275 ( .C1(n5503), .C2(PC_IN[14]), .A(n5502), .B(RST), .ZN(n5477)
         );
  INV_X1 U276 ( .A(n5477), .ZN(n281) );
  OAI211_X1 U277 ( .C1(n5512), .C2(PC_IN[8]), .A(n5511), .B(RST), .ZN(n5478)
         );
  INV_X1 U278 ( .A(n5478), .ZN(n280) );
  AOI211_X1 U279 ( .C1(n5481), .C2(n5480), .A(n5479), .B(n5324), .ZN(n58) );
  AOI211_X1 U280 ( .C1(n5484), .C2(n5483), .A(n5482), .B(n5324), .ZN(n57) );
  AOI211_X1 U281 ( .C1(n5487), .C2(n5486), .A(n5485), .B(n5324), .ZN(n56) );
  AOI211_X1 U282 ( .C1(n5490), .C2(n5489), .A(n5488), .B(n5324), .ZN(n55) );
  AOI211_X1 U283 ( .C1(n5493), .C2(n5492), .A(n5491), .B(n5324), .ZN(n54) );
  AOI211_X1 U284 ( .C1(n5496), .C2(n5495), .A(n5494), .B(n5325), .ZN(n53) );
  AOI211_X1 U285 ( .C1(n5499), .C2(n5498), .A(n5497), .B(n5325), .ZN(n52) );
  AOI211_X1 U286 ( .C1(n5502), .C2(n5501), .A(n5500), .B(n5325), .ZN(n51) );
  AOI211_X1 U287 ( .C1(n5505), .C2(n5504), .A(n5503), .B(n5325), .ZN(n50) );
  AOI211_X1 U288 ( .C1(n5508), .C2(n5507), .A(n5506), .B(n5325), .ZN(n49) );
  AOI211_X1 U289 ( .C1(n5511), .C2(n5510), .A(n5509), .B(n5325), .ZN(n48) );
  AOI211_X1 U290 ( .C1(n5514), .C2(n5513), .A(n5512), .B(n5324), .ZN(n47) );
  AOI222_X1 U291 ( .A1(n5548), .A2(N47), .B1(n5320), .B2(N220), .C1(n5547), 
        .C2(N82), .ZN(n5517) );
  INV_X1 U292 ( .A(n5517), .ZN(n46) );
  AOI222_X1 U293 ( .A1(n5548), .A2(N48), .B1(n5320), .B2(N221), .C1(n5322), 
        .C2(N83), .ZN(n5518) );
  INV_X1 U294 ( .A(n5518), .ZN(n45) );
  AOI222_X1 U295 ( .A1(n5548), .A2(N49), .B1(n5320), .B2(N222), .C1(n5547), 
        .C2(N84), .ZN(n5519) );
  INV_X1 U296 ( .A(n5519), .ZN(n44) );
  AOI222_X1 U297 ( .A1(n5548), .A2(N50), .B1(n5320), .B2(N223), .C1(n5322), 
        .C2(N85), .ZN(n5520) );
  INV_X1 U298 ( .A(n5520), .ZN(n43) );
  AOI222_X1 U299 ( .A1(n5548), .A2(N51), .B1(n5320), .B2(N224), .C1(n5547), 
        .C2(N86), .ZN(n5521) );
  INV_X1 U300 ( .A(n5521), .ZN(n42) );
  AOI222_X1 U301 ( .A1(n5548), .A2(N52), .B1(n5320), .B2(N225), .C1(n5322), 
        .C2(N87), .ZN(n5522) );
  INV_X1 U302 ( .A(n5522), .ZN(n41) );
  AOI222_X1 U303 ( .A1(n5548), .A2(N53), .B1(n5320), .B2(N226), .C1(n5547), 
        .C2(N88), .ZN(n5523) );
  INV_X1 U304 ( .A(n5523), .ZN(n40) );
  AOI222_X1 U305 ( .A1(n5548), .A2(N54), .B1(n5320), .B2(N227), .C1(n5547), 
        .C2(N89), .ZN(n5524) );
  INV_X1 U306 ( .A(n5524), .ZN(n39) );
  AOI222_X1 U307 ( .A1(n5548), .A2(N55), .B1(n5320), .B2(N228), .C1(n5547), 
        .C2(N90), .ZN(n5525) );
  INV_X1 U308 ( .A(n5525), .ZN(n38) );
  AOI222_X1 U309 ( .A1(n5548), .A2(N56), .B1(n5320), .B2(N229), .C1(n5547), 
        .C2(N91), .ZN(n5526) );
  INV_X1 U310 ( .A(n5526), .ZN(n37) );
  AOI222_X1 U311 ( .A1(n5548), .A2(N57), .B1(n5320), .B2(N230), .C1(n5547), 
        .C2(N92), .ZN(n5527) );
  INV_X1 U312 ( .A(n5527), .ZN(n36) );
  AOI222_X1 U313 ( .A1(n5548), .A2(N58), .B1(n5320), .B2(N231), .C1(n5547), 
        .C2(N93), .ZN(n5528) );
  INV_X1 U314 ( .A(n5528), .ZN(n35) );
  AOI222_X1 U315 ( .A1(n5548), .A2(N59), .B1(n5320), .B2(N232), .C1(n5322), 
        .C2(N94), .ZN(n5529) );
  INV_X1 U316 ( .A(n5529), .ZN(n34) );
  AOI222_X1 U317 ( .A1(n5548), .A2(N60), .B1(n5320), .B2(N233), .C1(n5322), 
        .C2(N95), .ZN(n5530) );
  INV_X1 U318 ( .A(n5530), .ZN(n33) );
  AOI222_X1 U319 ( .A1(n5548), .A2(N61), .B1(n5320), .B2(N234), .C1(n5322), 
        .C2(N96), .ZN(n5531) );
  INV_X1 U320 ( .A(n5531), .ZN(n32) );
  AOI222_X1 U321 ( .A1(n5548), .A2(N62), .B1(n5320), .B2(N235), .C1(n5322), 
        .C2(N97), .ZN(n5532) );
  INV_X1 U322 ( .A(n5532), .ZN(n31) );
  AOI222_X1 U323 ( .A1(n5548), .A2(N63), .B1(n5320), .B2(N236), .C1(n5322), 
        .C2(N98), .ZN(n5533) );
  INV_X1 U324 ( .A(n5533), .ZN(n30) );
  AOI222_X1 U325 ( .A1(n5548), .A2(N64), .B1(n5320), .B2(N237), .C1(n5322), 
        .C2(N99), .ZN(n5534) );
  INV_X1 U326 ( .A(n5534), .ZN(n29) );
  AOI222_X1 U327 ( .A1(n5548), .A2(N65), .B1(n5320), .B2(N238), .C1(n5322), 
        .C2(N100), .ZN(n5535) );
  INV_X1 U328 ( .A(n5535), .ZN(n28) );
  AOI222_X1 U329 ( .A1(n5548), .A2(N66), .B1(n5320), .B2(N239), .C1(n5547), 
        .C2(N101), .ZN(n5536) );
  INV_X1 U330 ( .A(n5536), .ZN(n27) );
  AOI222_X1 U331 ( .A1(n5548), .A2(N67), .B1(n5320), .B2(N240), .C1(n5322), 
        .C2(N102), .ZN(n5537) );
  INV_X1 U332 ( .A(n5537), .ZN(n26) );
  AOI222_X1 U333 ( .A1(n5548), .A2(N68), .B1(n5320), .B2(N241), .C1(n5547), 
        .C2(N103), .ZN(n5538) );
  INV_X1 U334 ( .A(n5538), .ZN(n25) );
  AOI222_X1 U335 ( .A1(n5548), .A2(N69), .B1(n5320), .B2(N242), .C1(n5322), 
        .C2(N104), .ZN(n5539) );
  INV_X1 U336 ( .A(n5539), .ZN(n24) );
  AOI222_X1 U337 ( .A1(n5548), .A2(N70), .B1(n5320), .B2(N243), .C1(n5547), 
        .C2(N105), .ZN(n5540) );
  INV_X1 U338 ( .A(n5540), .ZN(n23) );
  AOI222_X1 U339 ( .A1(n5548), .A2(N71), .B1(n5320), .B2(N244), .C1(n5322), 
        .C2(N106), .ZN(n5541) );
  INV_X1 U340 ( .A(n5541), .ZN(n22) );
  AOI222_X1 U341 ( .A1(n5548), .A2(N72), .B1(n5320), .B2(N245), .C1(n5322), 
        .C2(N107), .ZN(n5542) );
  INV_X1 U342 ( .A(n5542), .ZN(n21) );
  AOI222_X1 U343 ( .A1(n5548), .A2(N73), .B1(n5320), .B2(N246), .C1(n5322), 
        .C2(N108), .ZN(n5543) );
  INV_X1 U344 ( .A(n5543), .ZN(n20) );
  AOI222_X1 U345 ( .A1(n5548), .A2(N74), .B1(n5320), .B2(N247), .C1(n5322), 
        .C2(N109), .ZN(n5544) );
  INV_X1 U346 ( .A(n5544), .ZN(n4) );
  AOI222_X1 U347 ( .A1(n5548), .A2(N75), .B1(n5320), .B2(N248), .C1(n5322), 
        .C2(N110), .ZN(n5545) );
  INV_X1 U348 ( .A(n5545), .ZN(n3) );
  AOI222_X1 U349 ( .A1(n5548), .A2(N76), .B1(n5320), .B2(N249), .C1(n5322), 
        .C2(N111), .ZN(n5546) );
  INV_X1 U350 ( .A(n5546), .ZN(n2) );
  AOI222_X1 U351 ( .A1(n5548), .A2(N77), .B1(n5320), .B2(N250), .C1(n5322), 
        .C2(N112), .ZN(n5549) );
  INV_X1 U352 ( .A(n5549), .ZN(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_IF_ID ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module DLX_syn ( Clk, Rst, IRAM_DATA_OUT, DRAM_DATA_OUT, DRAM_DATA_IN, 
        DRAM_ADDRESS, DRAM_ENABLE, DRAM_RW, DRAM_SEL, IRAM_ADDRESS );
  input [31:0] IRAM_DATA_OUT;
  input [31:0] DRAM_DATA_OUT;
  output [31:0] DRAM_DATA_IN;
  output [11:0] DRAM_ADDRESS;
  output [2:0] DRAM_SEL;
  output [7:0] IRAM_ADDRESS;
  input Clk, Rst;
  output DRAM_ENABLE, DRAM_RW;
  wire   IR_CU_31, IR_CU_28, IR_CU_27, IR_CU_26, BR_EN_i, \WB_MUX_SEL_i[1] ,
         RF_WE_i, \CU_I/aluOpcode_i[4] , \CU_I/aluOpcode_i[3] ,
         \CU_I/aluOpcode_i[2] , \CU_I/aluOpcode_i[1] , \CU_I/aluOpcode_i[0] ,
         \CU_I/cw2[1] , \CU_I/cw[10] , \CU_I/cw[9] , \CU_I/cw[7] ,
         \CU_I/cw[6] , \CU_I/cw[4] , \CU_I/cw[3] , \CU_I/cw[1] , \CU_I/cw[0] ,
         \DataP/LMD_out[31] , \DataP/LMD_out[30] , \DataP/LMD_out[29] ,
         \DataP/LMD_out[28] , \DataP/LMD_out[27] , \DataP/LMD_out[26] ,
         \DataP/LMD_out[25] , \DataP/LMD_out[24] , \DataP/LMD_out[23] ,
         \DataP/LMD_out[22] , \DataP/LMD_out[21] , \DataP/LMD_out[20] ,
         \DataP/LMD_out[19] , \DataP/LMD_out[18] , \DataP/LMD_out[17] ,
         \DataP/LMD_out[16] , \DataP/LMD_out[15] , \DataP/LMD_out[14] ,
         \DataP/LMD_out[13] , \DataP/LMD_out[12] , \DataP/LMD_out[11] ,
         \DataP/LMD_out[10] , \DataP/LMD_out[9] , \DataP/LMD_out[8] ,
         \DataP/LMD_out[7] , \DataP/LMD_out[6] , \DataP/LMD_out[5] ,
         \DataP/LMD_out[4] , \DataP/LMD_out[3] , \DataP/LMD_out[2] ,
         \DataP/LMD_out[1] , \DataP/LMD_out[0] , \DataP/link_addr_W[31] ,
         \DataP/link_addr_W[30] , \DataP/link_addr_W[29] ,
         \DataP/link_addr_W[28] , \DataP/link_addr_W[27] ,
         \DataP/link_addr_W[26] , \DataP/link_addr_W[25] ,
         \DataP/link_addr_W[24] , \DataP/link_addr_W[23] ,
         \DataP/link_addr_W[22] , \DataP/link_addr_W[21] ,
         \DataP/link_addr_W[20] , \DataP/link_addr_W[19] ,
         \DataP/link_addr_W[18] , \DataP/link_addr_W[17] ,
         \DataP/link_addr_W[16] , \DataP/link_addr_W[15] ,
         \DataP/link_addr_W[14] , \DataP/link_addr_W[13] ,
         \DataP/link_addr_W[12] , \DataP/link_addr_W[11] ,
         \DataP/link_addr_W[10] , \DataP/link_addr_W[9] ,
         \DataP/link_addr_W[8] , \DataP/link_addr_W[7] ,
         \DataP/link_addr_W[6] , \DataP/link_addr_W[5] ,
         \DataP/link_addr_W[4] , \DataP/link_addr_W[3] ,
         \DataP/link_addr_W[2] , \DataP/link_addr_W[1] ,
         \DataP/link_addr_W[0] , \DataP/FWD_MUX_BR_S[1] ,
         \DataP/FWD_MUX_BR_S[0] , \DataP/alu_b_in[31] , \DataP/alu_b_in[30] ,
         \DataP/alu_b_in[29] , \DataP/alu_b_in[28] , \DataP/alu_b_in[27] ,
         \DataP/alu_b_in[26] , \DataP/alu_b_in[25] , \DataP/alu_b_in[24] ,
         \DataP/alu_b_in[23] , \DataP/alu_b_in[22] , \DataP/alu_b_in[21] ,
         \DataP/alu_b_in[20] , \DataP/alu_b_in[19] , \DataP/alu_b_in[18] ,
         \DataP/alu_b_in[17] , \DataP/alu_b_in[16] , \DataP/alu_b_in[15] ,
         \DataP/alu_b_in[13] , \DataP/alu_b_in[12] , \DataP/alu_b_in[10] ,
         \DataP/alu_b_in[9] , \DataP/alu_b_in[8] , \DataP/alu_b_in[7] ,
         \DataP/alu_b_in[6] , \DataP/alu_b_in[5] , \DataP/alu_b_in[3] ,
         \DataP/alu_b_in[2] , \DataP/alu_b_in[0] , \DataP/alu_a_in[31] ,
         \DataP/alu_a_in[30] , \DataP/alu_a_in[29] , \DataP/alu_a_in[28] ,
         \DataP/alu_a_in[27] , \DataP/alu_a_in[26] , \DataP/alu_a_in[25] ,
         \DataP/alu_a_in[24] , \DataP/alu_a_in[23] , \DataP/alu_a_in[22] ,
         \DataP/alu_a_in[21] , \DataP/alu_a_in[20] , \DataP/alu_a_in[19] ,
         \DataP/alu_a_in[18] , \DataP/alu_a_in[17] , \DataP/alu_a_in[16] ,
         \DataP/alu_a_in[15] , \DataP/alu_a_in[14] , \DataP/alu_a_in[13] ,
         \DataP/alu_a_in[12] , \DataP/alu_a_in[11] , \DataP/alu_a_in[10] ,
         \DataP/alu_a_in[9] , \DataP/alu_a_in[8] , \DataP/alu_a_in[7] ,
         \DataP/alu_a_in[6] , \DataP/alu_a_in[5] , \DataP/alu_a_in[4] ,
         \DataP/alu_a_in[3] , \DataP/alu_a_in[2] , \DataP/alu_a_in[1] ,
         \DataP/alu_a_in[0] , \DataP/alu_out_W[0] , \DataP/alu_out_W[1] ,
         \DataP/alu_out_W[2] , \DataP/alu_out_W[3] , \DataP/alu_out_W[4] ,
         \DataP/alu_out_W[5] , \DataP/alu_out_W[6] , \DataP/alu_out_W[7] ,
         \DataP/alu_out_W[8] , \DataP/alu_out_W[9] , \DataP/alu_out_W[10] ,
         \DataP/alu_out_W[11] , \DataP/alu_out_W[12] , \DataP/alu_out_W[13] ,
         \DataP/alu_out_W[14] , \DataP/alu_out_W[15] , \DataP/alu_out_W[16] ,
         \DataP/alu_out_W[17] , \DataP/alu_out_W[18] , \DataP/alu_out_W[19] ,
         \DataP/alu_out_W[20] , \DataP/alu_out_W[21] , \DataP/alu_out_W[22] ,
         \DataP/alu_out_W[23] , \DataP/alu_out_W[24] , \DataP/alu_out_W[25] ,
         \DataP/alu_out_W[26] , \DataP/alu_out_W[27] , \DataP/alu_out_W[28] ,
         \DataP/alu_out_W[29] , \DataP/alu_out_W[30] , \DataP/alu_out_W[31] ,
         \DataP/alu_out_M[12] , \DataP/alu_out_M[13] , \DataP/alu_out_M[14] ,
         \DataP/alu_out_M[15] , \DataP/alu_out_M[16] , \DataP/alu_out_M[17] ,
         \DataP/alu_out_M[18] , \DataP/alu_out_M[19] , \DataP/alu_out_M[20] ,
         \DataP/alu_out_M[21] , \DataP/alu_out_M[22] , \DataP/alu_out_M[23] ,
         \DataP/alu_out_M[24] , \DataP/alu_out_M[25] , \DataP/alu_out_M[26] ,
         \DataP/alu_out_M[27] , \DataP/alu_out_M[28] , \DataP/alu_out_M[29] ,
         \DataP/alu_out_M[30] , \DataP/alu_out_M[31] , \DataP/opcode_W[0] ,
         \DataP/opcode_W[1] , \DataP/opcode_W[2] , \DataP/opcode_W[3] ,
         \DataP/opcode_W[4] , \DataP/opcode_W[5] , \DataP/opcode_M[0] ,
         \DataP/opcode_M[1] , \DataP/opcode_M[3] , \DataP/opcode_M[4] ,
         \DataP/opcode_M[5] , \DataP/dest_M[0] , \DataP/dest_M[1] ,
         \DataP/dest_M[2] , \DataP/dest_M[3] , \DataP/dest_M[4] , \DataP/pr_E ,
         \DataP/opcode_E[0] , \DataP/opcode_E[3] , \DataP/opcode_E[4] ,
         \DataP/Rs2[4] , \DataP/Rs2[3] , \DataP/Rs2[2] , \DataP/Rs2[1] ,
         \DataP/Rs2[0] , \DataP/Rs1[1] , \DataP/Rs1[2] , \DataP/IMM_s[31] ,
         \DataP/IMM_s[24] , \DataP/IMM_s[23] , \DataP/IMM_s[22] ,
         \DataP/IMM_s[21] , \DataP/IMM_s[20] , \DataP/IMM_s[19] ,
         \DataP/IMM_s[18] , \DataP/IMM_s[17] , \DataP/IMM_s[16] ,
         \DataP/B_s[0] , \DataP/B_s[1] , \DataP/B_s[2] , \DataP/B_s[3] ,
         \DataP/B_s[4] , \DataP/B_s[5] , \DataP/B_s[6] , \DataP/B_s[7] ,
         \DataP/B_s[8] , \DataP/B_s[9] , \DataP/B_s[10] , \DataP/B_s[11] ,
         \DataP/B_s[12] , \DataP/B_s[13] , \DataP/B_s[14] , \DataP/B_s[15] ,
         \DataP/B_s[16] , \DataP/B_s[17] , \DataP/B_s[18] , \DataP/B_s[19] ,
         \DataP/B_s[20] , \DataP/B_s[21] , \DataP/B_s[22] , \DataP/B_s[23] ,
         \DataP/B_s[24] , \DataP/B_s[25] , \DataP/B_s[26] , \DataP/B_s[27] ,
         \DataP/B_s[28] , \DataP/B_s[29] , \DataP/B_s[30] , \DataP/B_s[31] ,
         \DataP/A_s[0] , \DataP/A_s[1] , \DataP/A_s[2] , \DataP/A_s[3] ,
         \DataP/A_s[4] , \DataP/A_s[5] , \DataP/A_s[6] , \DataP/A_s[7] ,
         \DataP/A_s[8] , \DataP/A_s[9] , \DataP/A_s[10] , \DataP/A_s[11] ,
         \DataP/A_s[12] , \DataP/A_s[13] , \DataP/A_s[14] , \DataP/A_s[15] ,
         \DataP/A_s[16] , \DataP/A_s[17] , \DataP/A_s[18] , \DataP/A_s[19] ,
         \DataP/A_s[20] , \DataP/A_s[21] , \DataP/A_s[22] , \DataP/A_s[23] ,
         \DataP/A_s[24] , \DataP/A_s[25] , \DataP/A_s[26] , \DataP/A_s[27] ,
         \DataP/A_s[28] , \DataP/A_s[29] , \DataP/A_s[30] , \DataP/A_s[31] ,
         \DataP/imm_out[31] , \DataP/imm_out[24] , \DataP/imm_out[23] ,
         \DataP/imm_out[22] , \DataP/imm_out[21] , \DataP/imm_out[20] ,
         \DataP/imm_out[19] , \DataP/imm_out[18] , \DataP/imm_out[17] ,
         \DataP/imm_out[16] , \DataP/b_out[31] , \DataP/b_out[30] ,
         \DataP/b_out[29] , \DataP/b_out[28] , \DataP/b_out[27] ,
         \DataP/b_out[26] , \DataP/b_out[25] , \DataP/b_out[24] ,
         \DataP/b_out[23] , \DataP/b_out[22] , \DataP/b_out[21] ,
         \DataP/b_out[20] , \DataP/b_out[19] , \DataP/b_out[18] ,
         \DataP/b_out[17] , \DataP/b_out[16] , \DataP/b_out[15] ,
         \DataP/b_out[14] , \DataP/b_out[13] , \DataP/b_out[12] ,
         \DataP/b_out[11] , \DataP/b_out[10] , \DataP/b_out[9] ,
         \DataP/b_out[8] , \DataP/b_out[7] , \DataP/b_out[6] ,
         \DataP/b_out[5] , \DataP/b_out[4] , \DataP/b_out[3] ,
         \DataP/b_out[2] , \DataP/b_out[1] , \DataP/b_out[0] ,
         \DataP/a_out[31] , \DataP/a_out[30] , \DataP/a_out[29] ,
         \DataP/a_out[28] , \DataP/a_out[27] , \DataP/a_out[26] ,
         \DataP/a_out[25] , \DataP/a_out[24] , \DataP/a_out[23] ,
         \DataP/a_out[22] , \DataP/a_out[21] , \DataP/a_out[20] ,
         \DataP/a_out[19] , \DataP/a_out[18] , \DataP/a_out[17] ,
         \DataP/a_out[16] , \DataP/a_out[15] , \DataP/a_out[14] ,
         \DataP/a_out[13] , \DataP/a_out[12] , \DataP/a_out[11] ,
         \DataP/a_out[10] , \DataP/a_out[9] , \DataP/a_out[8] ,
         \DataP/a_out[7] , \DataP/a_out[6] , \DataP/a_out[5] ,
         \DataP/a_out[4] , \DataP/a_out[3] , \DataP/a_out[2] ,
         \DataP/a_out[1] , \DataP/a_out[0] , \DataP/WB[31] , \DataP/WB[30] ,
         \DataP/WB[29] , \DataP/WB[28] , \DataP/WB[27] , \DataP/WB[26] ,
         \DataP/WB[25] , \DataP/WB[24] , \DataP/WB[23] , \DataP/WB[22] ,
         \DataP/WB[21] , \DataP/WB[20] , \DataP/WB[19] , \DataP/WB[18] ,
         \DataP/WB[17] , \DataP/WB[16] , \DataP/WB[15] , \DataP/WB[14] ,
         \DataP/WB[13] , \DataP/WB[12] , \DataP/WB[11] , \DataP/WB[10] ,
         \DataP/WB[9] , \DataP/WB[8] , \DataP/WB[7] , \DataP/WB[6] ,
         \DataP/WB[5] , \DataP/WB[4] , \DataP/WB[3] , \DataP/WB[2] ,
         \DataP/WB[1] , \DataP/WB[0] , \DataP/add_D[0] , \DataP/add_D[1] ,
         \DataP/add_D[2] , \DataP/add_D[3] , \DataP/add_D[4] ,
         \DataP/dest_D[4] , \DataP/dest_D[3] , \DataP/dest_D[2] ,
         \DataP/dest_D[1] , \DataP/dest_D[0] , \DataP/add_S2[0] ,
         \DataP/add_S2[1] , \DataP/add_S2[2] , \DataP/add_S2[3] ,
         \DataP/add_S2[4] , \DataP/prediction , \DataP/npc_mux_sel ,
         \DataP/link_addr_F[31] , \DataP/link_addr_F[30] ,
         \DataP/link_addr_F[29] , \DataP/link_addr_F[28] ,
         \DataP/link_addr_F[27] , \DataP/link_addr_F[26] ,
         \DataP/link_addr_F[25] , \DataP/link_addr_F[24] ,
         \DataP/link_addr_F[23] , \DataP/link_addr_F[22] ,
         \DataP/link_addr_F[21] , \DataP/link_addr_F[20] ,
         \DataP/link_addr_F[19] , \DataP/link_addr_F[18] ,
         \DataP/link_addr_F[17] , \DataP/link_addr_F[16] ,
         \DataP/link_addr_F[15] , \DataP/link_addr_F[14] ,
         \DataP/link_addr_F[13] , \DataP/link_addr_F[12] ,
         \DataP/link_addr_F[11] , \DataP/link_addr_F[10] ,
         \DataP/link_addr_F[9] , \DataP/link_addr_F[8] ,
         \DataP/link_addr_F[7] , \DataP/link_addr_F[6] ,
         \DataP/link_addr_F[5] , \DataP/link_addr_F[4] ,
         \DataP/link_addr_F[3] , \DataP/link_addr_F[2] ,
         \DataP/link_addr_F[1] , \DataP/link_addr_F[0] , \DataP/npc_pre[31] ,
         \DataP/npc_pre[30] , \DataP/npc_pre[29] , \DataP/npc_pre[28] ,
         \DataP/npc_pre[27] , \DataP/npc_pre[26] , \DataP/npc_pre[25] ,
         \DataP/npc_pre[24] , \DataP/npc_pre[23] , \DataP/npc_pre[22] ,
         \DataP/npc_pre[21] , \DataP/npc_pre[20] , \DataP/npc_pre[19] ,
         \DataP/npc_pre[18] , \DataP/npc_pre[17] , \DataP/npc_pre[16] ,
         \DataP/npc_pre[15] , \DataP/npc_pre[14] , \DataP/npc_pre[13] ,
         \DataP/npc_pre[12] , \DataP/npc_pre[11] , \DataP/npc_pre[10] ,
         \DataP/npc_pre[9] , \DataP/npc_pre[8] , \DataP/npc_pre[7] ,
         \DataP/npc_pre[6] , \DataP/npc_pre[5] , \DataP/npc_pre[4] ,
         \DataP/npc_pre[3] , \DataP/npc_pre[2] , \DataP/npc_pre[1] ,
         \DataP/npc_pre[0] , \DataP/right_br , \DataP/wrong_br ,
         \DataP/ir_E[15] , \DataP/ir_E[14] , \DataP/ir_E[13] ,
         \DataP/ir_E[12] , \DataP/ir_E[11] , \DataP/ir_E[10] , \DataP/ir_E[9] ,
         \DataP/ir_E[8] , \DataP/ir_E[7] , \DataP/ir_E[6] , \DataP/ir_E[5] ,
         \DataP/ir_E[4] , \DataP/ir_E[3] , \DataP/ir_E[2] , \DataP/ir_E[1] ,
         \DataP/ir_E[0] , \DataP/npc_M[31] , \DataP/npc_M[30] ,
         \DataP/npc_M[29] , \DataP/npc_M[28] , \DataP/npc_M[27] ,
         \DataP/npc_M[26] , \DataP/npc_M[25] , \DataP/npc_M[24] ,
         \DataP/npc_M[23] , \DataP/npc_M[22] , \DataP/npc_M[21] ,
         \DataP/npc_M[20] , \DataP/npc_M[19] , \DataP/npc_M[18] ,
         \DataP/npc_M[17] , \DataP/npc_M[16] , \DataP/npc_M[15] ,
         \DataP/npc_M[14] , \DataP/npc_M[13] , \DataP/npc_M[12] ,
         \DataP/npc_M[11] , \DataP/npc_M[10] , \DataP/npc_M[9] ,
         \DataP/npc_M[8] , \DataP/npc_M[7] , \DataP/npc_M[6] ,
         \DataP/npc_M[5] , \DataP/npc_M[4] , \DataP/npc_M[3] ,
         \DataP/npc_M[2] , \DataP/npc_M[1] , \DataP/npc_M[0] ,
         \DataP/pc_out_0 , \DataP/pc_out_1 , \DataP/pc_out[10] ,
         \DataP/pc_out[11] , \DataP/pc_out[12] , \DataP/pc_out[13] ,
         \DataP/pc_out[14] , \DataP/pc_out[15] , \DataP/pc_out[16] ,
         \DataP/pc_out[17] , \DataP/pc_out[18] , \DataP/pc_out[19] ,
         \DataP/pc_out[20] , \DataP/pc_out[21] , \DataP/pc_out[22] ,
         \DataP/pc_out[23] , \DataP/pc_out[24] , \DataP/pc_out[25] ,
         \DataP/pc_out[26] , \DataP/pc_out[27] , \DataP/pc_out[28] ,
         \DataP/pc_out[29] , \DataP/pc_out[30] , \DataP/pc_out[31] ,
         \DataP/npc[0] , \DataP/npc[1] , \DataP/npc[2] , \DataP/npc[3] ,
         \DataP/npc[4] , \DataP/npc[5] , \DataP/npc[6] , \DataP/npc[7] ,
         \DataP/npc[8] , \DataP/npc[9] , \DataP/npc[10] , \DataP/npc[11] ,
         \DataP/npc[12] , \DataP/npc[13] , \DataP/npc[14] , \DataP/npc[15] ,
         \DataP/npc[16] , \DataP/npc[17] , \DataP/npc[18] , \DataP/npc[19] ,
         \DataP/npc[20] , \DataP/npc[21] , \DataP/npc[22] , \DataP/npc[23] ,
         \DataP/npc[24] , \DataP/npc[25] , \DataP/npc[26] , \DataP/npc[27] ,
         \DataP/npc[28] , \DataP/npc[29] , \DataP/npc[30] , \DataP/npc[31] ,
         \DataP/IR1[11] , \DataP/IR1[12] , \DataP/IR1[13] , \DataP/IR1[14] ,
         \DataP/IR1[15] , \DataP/IR1[21] , \DataP/IR1[22] , \DataP/IR1[23] ,
         \DataP/IR1[24] , \DataP/IR1[25] , \DataP/PC_reg/N33 ,
         \DataP/PC_reg/N32 , \DataP/PC_reg/N31 , \DataP/PC_reg/N30 ,
         \DataP/PC_reg/N29 , \DataP/PC_reg/N28 , \DataP/PC_reg/N27 ,
         \DataP/PC_reg/N26 , \DataP/PC_reg/N25 , \DataP/PC_reg/N24 ,
         \DataP/PC_reg/N23 , \DataP/PC_reg/N22 , \DataP/PC_reg/N21 ,
         \DataP/PC_reg/N20 , \DataP/PC_reg/N19 , \DataP/PC_reg/N18 ,
         \DataP/PC_reg/N17 , \DataP/PC_reg/N16 , \DataP/PC_reg/N15 ,
         \DataP/PC_reg/N14 , \DataP/PC_reg/N13 , \DataP/PC_reg/N12 ,
         \DataP/PC_reg/N11 , \DataP/PC_reg/N10 , \DataP/PC_reg/N9 ,
         \DataP/PC_reg/N8 , \DataP/PC_reg/N7 , \DataP/PC_reg/N6 ,
         \DataP/PC_reg/N5 , \DataP/PC_reg/N4 , \DataP/PC_reg/N3 ,
         \DataP/PC_reg/N2 , \DataP/NPC_add/N32 , \DataP/NPC_add/N31 ,
         \DataP/NPC_add/N30 , \DataP/NPC_add/N29 , \DataP/NPC_add/N28 ,
         \DataP/NPC_add/N27 , \DataP/NPC_add/N26 , \DataP/NPC_add/N25 ,
         \DataP/NPC_add/N24 , \DataP/NPC_add/N23 , \DataP/NPC_add/N22 ,
         \DataP/NPC_add/N21 , \DataP/NPC_add/N20 , \DataP/NPC_add/N19 ,
         \DataP/NPC_add/N18 , \DataP/NPC_add/N17 , \DataP/NPC_add/N16 ,
         \DataP/NPC_add/N15 , \DataP/NPC_add/N14 , \DataP/NPC_add/N13 ,
         \DataP/NPC_add/N12 , \DataP/NPC_add/N11 , \DataP/NPC_add/N10 ,
         \DataP/NPC_add/N9 , \DataP/NPC_add/N8 , \DataP/NPC_add/N7 ,
         \DataP/NPC_add/N6 , \DataP/NPC_add/N5 , \DataP/NPC_add/N4 ,
         \DataP/NPC_add/N3 , \DataP/NPC_add/N2 , \DataP/NPC_add/N1 ,
         \DataP/NPC_add/N0 , \DataP/IF_IDs/net834167 ,
         \DataP/FORWARDING_BR/N12 , \DataP/ALU_C/shifter/N107 ,
         \DataP/ALU_C/shifter/N106 , \DataP/ALU_C/shifter/N105 ,
         \DataP/ALU_C/shifter/N104 , \DataP/ALU_C/shifter/N103 ,
         \DataP/ALU_C/shifter/N102 , \DataP/ALU_C/shifter/N101 ,
         \DataP/ALU_C/shifter/N100 , \DataP/ALU_C/shifter/N99 ,
         \DataP/ALU_C/shifter/N98 , \DataP/ALU_C/shifter/N97 ,
         \DataP/ALU_C/shifter/N96 , \DataP/ALU_C/shifter/N95 ,
         \DataP/ALU_C/shifter/N94 , \DataP/ALU_C/shifter/N93 ,
         \DataP/ALU_C/shifter/N92 , \DataP/ALU_C/shifter/N89 ,
         \DataP/ALU_C/shifter/N83 , \DataP/ALU_C/shifter/N82 ,
         \DataP/ALU_C/shifter/N81 , \DataP/ALU_C/shifter/N80 ,
         \DataP/ALU_C/shifter/N79 , \DataP/ALU_C/shifter/N78 ,
         \DataP/ALU_C/shifter/N77 , \DataP/ALU_C/shifter/N76 ,
         \DataP/ALU_C/shifter/N75 , \DataP/ALU_C/shifter/N74 ,
         \DataP/ALU_C/shifter/N73 , \DataP/ALU_C/shifter/N72 ,
         \DataP/ALU_C/shifter/N71 , \DataP/ALU_C/shifter/N70 ,
         \DataP/ALU_C/shifter/N69 , \DataP/ALU_C/shifter/N68 ,
         \DataP/ALU_C/shifter/N67 , \DataP/ALU_C/shifter/N66 ,
         \DataP/ALU_C/shifter/N65 , \DataP/ALU_C/shifter/N64 ,
         \DataP/ALU_C/shifter/N63 , \DataP/ALU_C/shifter/N62 ,
         \DataP/ALU_C/shifter/N61 , \DataP/ALU_C/shifter/N60 ,
         \DataP/ALU_C/shifter/N51 , \DataP/ALU_C/shifter/N50 ,
         \DataP/ALU_C/shifter/N49 , \DataP/ALU_C/shifter/N48 ,
         \DataP/ALU_C/shifter/N47 , \DataP/ALU_C/shifter/N46 ,
         \DataP/ALU_C/shifter/N43 , \DataP/ALU_C/shifter/N42 ,
         \DataP/ALU_C/shifter/N40 , \DataP/ALU_C/shifter/N39 ,
         \DataP/ALU_C/shifter/N38 , \DataP/ALU_C/shifter/N37 ,
         \DataP/ALU_C/shifter/N36 , \DataP/ALU_C/shifter/N34 ,
         \DataP/ALU_C/shifter/N33 , \DataP/ALU_C/shifter/N32 ,
         \DataP/ALU_C/shifter/N31 , \DataP/ALU_C/shifter/N30 ,
         \DataP/ALU_C/shifter/N29 , \DataP/ALU_C/shifter/N28 ,
         \DataP/ALU_C/shifter/N19 , \DataP/ALU_C/comp/N24 , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n296, n297, n299, n300, n301, n303, n304, n308, n309,
         n311, n313, n317, n319, n322, n323, n326, n330, n332, n333, n337,
         n340, n341, n345, n350, n353, n354, n355, n356, n357, n358, n399,
         n432, n443, n476, n477, n478, n479, n480, n482, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n497, n504, n510,
         n514, n515, n516, n520, n521, n523, n524, n528, n529, n530, n536,
         n538, n540, n606, n1357, n1371, n1448, \sra_131/SH[4] ,
         \sra_131/SH[1] , \lt_x_135/B[4] , \lt_x_134/B[5] , \lt_x_134/B[4] ,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023;
  wire   [10:0] IR_CU;
  wire   [4:0] ALU_OPCODE_i;

  register_file_N32_addBit5 \DataP/Reg_F  ( .RESET(Rst), .RE(1'b1), .WE(
        RF_WE_i), .ADD_WR({\DataP/add_D[4] , \DataP/add_D[3] , n1955, n1892, 
        n1852}), .ADD_RDA({n494, n493, n492, n491, n490}), .ADD_RDB({
        \DataP/add_S2[4] , \DataP/add_S2[3] , \DataP/add_S2[2] , 
        \DataP/add_S2[1] , \DataP/add_S2[0] }), .DATAIN({\DataP/WB[31] , 
        \DataP/WB[30] , \DataP/WB[29] , \DataP/WB[28] , \DataP/WB[27] , 
        \DataP/WB[26] , \DataP/WB[25] , \DataP/WB[24] , \DataP/WB[23] , 
        \DataP/WB[22] , \DataP/WB[21] , \DataP/WB[20] , \DataP/WB[19] , 
        \DataP/WB[18] , \DataP/WB[17] , \DataP/WB[16] , \DataP/WB[15] , 
        \DataP/WB[14] , \DataP/WB[13] , \DataP/WB[12] , \DataP/WB[11] , 
        \DataP/WB[10] , \DataP/WB[9] , \DataP/WB[8] , \DataP/WB[7] , 
        \DataP/WB[6] , \DataP/WB[5] , \DataP/WB[4] , \DataP/WB[3] , 
        \DataP/WB[2] , \DataP/WB[1] , \DataP/WB[0] }), .OUTA({
        \DataP/a_out[31] , \DataP/a_out[30] , \DataP/a_out[29] , 
        \DataP/a_out[28] , \DataP/a_out[27] , \DataP/a_out[26] , 
        \DataP/a_out[25] , \DataP/a_out[24] , \DataP/a_out[23] , 
        \DataP/a_out[22] , \DataP/a_out[21] , \DataP/a_out[20] , 
        \DataP/a_out[19] , \DataP/a_out[18] , \DataP/a_out[17] , 
        \DataP/a_out[16] , \DataP/a_out[15] , \DataP/a_out[14] , 
        \DataP/a_out[13] , \DataP/a_out[12] , \DataP/a_out[11] , 
        \DataP/a_out[10] , \DataP/a_out[9] , \DataP/a_out[8] , 
        \DataP/a_out[7] , \DataP/a_out[6] , \DataP/a_out[5] , \DataP/a_out[4] , 
        \DataP/a_out[3] , \DataP/a_out[2] , \DataP/a_out[1] , \DataP/a_out[0] }), .OUTB({\DataP/b_out[31] , \DataP/b_out[30] , \DataP/b_out[29] , 
        \DataP/b_out[28] , \DataP/b_out[27] , \DataP/b_out[26] , 
        \DataP/b_out[25] , \DataP/b_out[24] , \DataP/b_out[23] , 
        \DataP/b_out[22] , \DataP/b_out[21] , \DataP/b_out[20] , 
        \DataP/b_out[19] , \DataP/b_out[18] , \DataP/b_out[17] , 
        \DataP/b_out[16] , \DataP/b_out[15] , \DataP/b_out[14] , 
        \DataP/b_out[13] , \DataP/b_out[12] , \DataP/b_out[11] , 
        \DataP/b_out[10] , \DataP/b_out[9] , \DataP/b_out[8] , 
        \DataP/b_out[7] , \DataP/b_out[6] , \DataP/b_out[5] , \DataP/b_out[4] , 
        \DataP/b_out[3] , \DataP/b_out[2] , \DataP/b_out[1] , \DataP/b_out[0] }) );
  branch_predictor \DataP/BR_pred  ( .RST(Rst), .PC_IN({\DataP/pc_out[31] , 
        \DataP/pc_out[30] , \DataP/pc_out[29] , \DataP/pc_out[28] , 
        \DataP/pc_out[27] , \DataP/pc_out[26] , \DataP/pc_out[25] , 
        \DataP/pc_out[24] , \DataP/pc_out[23] , \DataP/pc_out[22] , 
        \DataP/pc_out[21] , \DataP/pc_out[20] , \DataP/pc_out[19] , 
        \DataP/pc_out[18] , \DataP/pc_out[17] , \DataP/pc_out[16] , 
        \DataP/pc_out[15] , \DataP/pc_out[14] , \DataP/pc_out[13] , 
        \DataP/pc_out[12] , \DataP/pc_out[11] , \DataP/pc_out[10] , 
        IRAM_ADDRESS, \DataP/pc_out_1 , \DataP/pc_out_0 }), .PC_FAIL({
        \DataP/npc_M[31] , \DataP/npc_M[30] , \DataP/npc_M[29] , 
        \DataP/npc_M[28] , \DataP/npc_M[27] , \DataP/npc_M[26] , 
        \DataP/npc_M[25] , \DataP/npc_M[24] , \DataP/npc_M[23] , 
        \DataP/npc_M[22] , \DataP/npc_M[21] , \DataP/npc_M[20] , 
        \DataP/npc_M[19] , \DataP/npc_M[18] , \DataP/npc_M[17] , 
        \DataP/npc_M[16] , \DataP/npc_M[15] , \DataP/npc_M[14] , 
        \DataP/npc_M[13] , \DataP/npc_M[12] , \DataP/npc_M[11] , 
        \DataP/npc_M[10] , \DataP/npc_M[9] , \DataP/npc_M[8] , 
        \DataP/npc_M[7] , \DataP/npc_M[6] , \DataP/npc_M[5] , \DataP/npc_M[4] , 
        \DataP/npc_M[3] , \DataP/npc_M[2] , \DataP/npc_M[1] , \DataP/npc_M[0] }), .IR_IN({IRAM_DATA_OUT[31:27], 1'b0, IRAM_DATA_OUT[25:0]}), .IR_FAIL({
        \DataP/ir_E[15] , \DataP/ir_E[14] , \DataP/ir_E[13] , \DataP/ir_E[12] , 
        \DataP/ir_E[11] , \DataP/ir_E[10] , \DataP/ir_E[9] , \DataP/ir_E[8] , 
        \DataP/ir_E[7] , \DataP/ir_E[6] , \DataP/ir_E[5] , \DataP/ir_E[4] , 
        \DataP/ir_E[3] , \DataP/ir_E[2] , \DataP/ir_E[1] , \DataP/ir_E[0] }), 
        .WRONG_PRE(\DataP/wrong_br ), .RIGHT_PRE(\DataP/right_br ), .NPC_OUT({
        \DataP/npc_pre[31] , \DataP/npc_pre[30] , \DataP/npc_pre[29] , 
        \DataP/npc_pre[28] , \DataP/npc_pre[27] , \DataP/npc_pre[26] , 
        \DataP/npc_pre[25] , \DataP/npc_pre[24] , \DataP/npc_pre[23] , 
        \DataP/npc_pre[22] , \DataP/npc_pre[21] , \DataP/npc_pre[20] , 
        \DataP/npc_pre[19] , \DataP/npc_pre[18] , \DataP/npc_pre[17] , 
        \DataP/npc_pre[16] , \DataP/npc_pre[15] , \DataP/npc_pre[14] , 
        \DataP/npc_pre[13] , \DataP/npc_pre[12] , \DataP/npc_pre[11] , 
        \DataP/npc_pre[10] , \DataP/npc_pre[9] , \DataP/npc_pre[8] , 
        \DataP/npc_pre[7] , \DataP/npc_pre[6] , \DataP/npc_pre[5] , 
        \DataP/npc_pre[4] , \DataP/npc_pre[3] , \DataP/npc_pre[2] , 
        \DataP/npc_pre[1] , \DataP/npc_pre[0] }), .LINK_ADD({
        \DataP/link_addr_F[31] , \DataP/link_addr_F[30] , 
        \DataP/link_addr_F[29] , \DataP/link_addr_F[28] , 
        \DataP/link_addr_F[27] , \DataP/link_addr_F[26] , 
        \DataP/link_addr_F[25] , \DataP/link_addr_F[24] , 
        \DataP/link_addr_F[23] , \DataP/link_addr_F[22] , 
        \DataP/link_addr_F[21] , \DataP/link_addr_F[20] , 
        \DataP/link_addr_F[19] , \DataP/link_addr_F[18] , 
        \DataP/link_addr_F[17] , \DataP/link_addr_F[16] , 
        \DataP/link_addr_F[15] , \DataP/link_addr_F[14] , 
        \DataP/link_addr_F[13] , \DataP/link_addr_F[12] , 
        \DataP/link_addr_F[11] , \DataP/link_addr_F[10] , 
        \DataP/link_addr_F[9] , \DataP/link_addr_F[8] , \DataP/link_addr_F[7] , 
        \DataP/link_addr_F[6] , \DataP/link_addr_F[5] , \DataP/link_addr_F[4] , 
        \DataP/link_addr_F[3] , \DataP/link_addr_F[2] , \DataP/link_addr_F[1] , 
        \DataP/link_addr_F[0] }), .SEL(\DataP/npc_mux_sel ), .TAKEN(
        \DataP/prediction ) );
  SNPS_CLOCK_GATE_HIGH_IF_ID \DataP/IF_IDs/clk_gate_PR_OUT_reg  ( .CLK(Clk), 
        .EN(n1448), .ENCLK(\DataP/IF_IDs/net834167 ), .TE(1'b0) );
  DLH_X1 \DataP/NPC_add/outPC_reg[0]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N1 ), .Q(\DataP/npc[0] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[1]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N2 ), .Q(\DataP/npc[1] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[2]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N3 ), .Q(\DataP/npc[2] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[3]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N4 ), .Q(\DataP/npc[3] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[4]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N5 ), .Q(\DataP/npc[4] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[5]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N6 ), .Q(\DataP/npc[5] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[6]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N7 ), .Q(\DataP/npc[6] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[7]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N8 ), .Q(\DataP/npc[7] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[8]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N9 ), .Q(\DataP/npc[8] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[9]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N10 ), .Q(\DataP/npc[9] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[10]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N11 ), .Q(\DataP/npc[10] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[11]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N12 ), .Q(\DataP/npc[11] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[12]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N13 ), .Q(\DataP/npc[12] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[13]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N14 ), .Q(\DataP/npc[13] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[14]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N15 ), .Q(\DataP/npc[14] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[15]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N16 ), .Q(\DataP/npc[15] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[16]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N17 ), .Q(\DataP/npc[16] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[17]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N18 ), .Q(\DataP/npc[17] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[18]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N19 ), .Q(\DataP/npc[18] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[19]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N20 ), .Q(\DataP/npc[19] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[20]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N21 ), .Q(\DataP/npc[20] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[21]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N22 ), .Q(\DataP/npc[21] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[22]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N23 ), .Q(\DataP/npc[22] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[23]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N24 ), .Q(\DataP/npc[23] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[24]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N25 ), .Q(\DataP/npc[24] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[25]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N26 ), .Q(\DataP/npc[25] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[26]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N27 ), .Q(\DataP/npc[26] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[27]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N28 ), .Q(\DataP/npc[27] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[28]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N29 ), .Q(\DataP/npc[28] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[29]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N30 ), .Q(\DataP/npc[29] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[30]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N31 ), .Q(\DataP/npc[30] ) );
  DLH_X1 \DataP/NPC_add/outPC_reg[31]  ( .G(\DataP/NPC_add/N0 ), .D(
        \DataP/NPC_add/N32 ), .Q(\DataP/npc[31] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[0]  ( .D(DRAM_DATA_OUT[0]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[0] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[1]  ( .D(DRAM_DATA_OUT[1]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[1] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[2]  ( .D(DRAM_DATA_OUT[2]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[2] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[3]  ( .D(DRAM_DATA_OUT[3]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[3] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[4]  ( .D(DRAM_DATA_OUT[4]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[4] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[5]  ( .D(DRAM_DATA_OUT[5]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[5] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[6]  ( .D(DRAM_DATA_OUT[6]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[6] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[7]  ( .D(DRAM_DATA_OUT[7]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[7] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[8]  ( .D(DRAM_DATA_OUT[8]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[8] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[9]  ( .D(DRAM_DATA_OUT[9]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[9] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[10]  ( .D(DRAM_DATA_OUT[10]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[10] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[11]  ( .D(DRAM_DATA_OUT[11]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[11] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[12]  ( .D(DRAM_DATA_OUT[12]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[12] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[13]  ( .D(DRAM_DATA_OUT[13]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[13] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[14]  ( .D(DRAM_DATA_OUT[14]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[14] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[15]  ( .D(DRAM_DATA_OUT[15]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[15] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[16]  ( .D(DRAM_DATA_OUT[16]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[16] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[17]  ( .D(DRAM_DATA_OUT[17]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[17] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[18]  ( .D(DRAM_DATA_OUT[18]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[18] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[19]  ( .D(DRAM_DATA_OUT[19]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[19] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[20]  ( .D(DRAM_DATA_OUT[20]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[20] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[21]  ( .D(DRAM_DATA_OUT[21]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[21] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[22]  ( .D(DRAM_DATA_OUT[22]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[22] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[23]  ( .D(DRAM_DATA_OUT[23]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[23] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[24]  ( .D(DRAM_DATA_OUT[24]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[24] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[25]  ( .D(DRAM_DATA_OUT[25]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[25] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[26]  ( .D(DRAM_DATA_OUT[26]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[26] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[27]  ( .D(DRAM_DATA_OUT[27]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[27] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[28]  ( .D(DRAM_DATA_OUT[28]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[28] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[29]  ( .D(DRAM_DATA_OUT[29]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[29] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[30]  ( .D(DRAM_DATA_OUT[30]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[30] ) );
  DFFR_X1 \DataP/MEM_WB_s/LMD_OUT_reg[31]  ( .D(DRAM_DATA_OUT[31]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/LMD_out[31] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[31]  ( .D(\DataP/alu_out_M[31] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[31] ), .QN(n2267) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[31]  ( .D(\DataP/link_addr_F[31] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n293) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[31]  ( .D(n293), .CK(Clk), .SN(Rst), .Q(
        n292) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[31]  ( .D(n292), .CK(Clk), .SN(Rst), 
        .Q(n291) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[31]  ( .D(n291), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[31] ) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[0]  ( .D(\DataP/b_out[0] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[0] ), .QN(n290) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[0]  ( .D(n290), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[0]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[1]  ( .D(\DataP/b_out[1] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[1] ), .QN(n289) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[1]  ( .D(n289), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[1]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[2]  ( .D(\DataP/b_out[2] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[2] ), .QN(n288) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[2]  ( .D(n288), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[2]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[3]  ( .D(\DataP/b_out[3] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[3] ), .QN(n287) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[3]  ( .D(n287), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[3]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[4]  ( .D(\DataP/b_out[4] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[4] ), .QN(n286) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[4]  ( .D(n286), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[4]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[5]  ( .D(\DataP/b_out[5] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[5] ), .QN(n285) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[5]  ( .D(n285), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[5]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[6]  ( .D(\DataP/b_out[6] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[6] ), .QN(n284) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[6]  ( .D(n284), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[6]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[7]  ( .D(\DataP/b_out[7] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[7] ), .QN(n283) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[7]  ( .D(n283), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[7]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[8]  ( .D(\DataP/b_out[8] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[8] ), .QN(n282) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[8]  ( .D(n282), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[8]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[9]  ( .D(\DataP/b_out[9] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[9] ), .QN(n281) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[9]  ( .D(n281), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[9]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[10]  ( .D(\DataP/b_out[10] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[10] ), .QN(n280) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[10]  ( .D(n280), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[10]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[11]  ( .D(\DataP/b_out[11] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[11] ), .QN(n279) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[11]  ( .D(n279), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[11]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[12]  ( .D(\DataP/b_out[12] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[12] ), .QN(n278) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[12]  ( .D(n278), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[12]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[13]  ( .D(\DataP/b_out[13] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[13] ), .QN(n277) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[13]  ( .D(n277), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[13]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[14]  ( .D(\DataP/b_out[14] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[14] ), .QN(n276) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[14]  ( .D(n276), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[14]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[15]  ( .D(\DataP/b_out[15] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[15] ), .QN(n275) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[15]  ( .D(n275), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[15]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[16]  ( .D(\DataP/b_out[16] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[16] ), .QN(n274) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[16]  ( .D(n274), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[16]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[17]  ( .D(\DataP/b_out[17] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[17] ), .QN(n273) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[17]  ( .D(n273), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[17]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[18]  ( .D(\DataP/b_out[18] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[18] ), .QN(n272) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[18]  ( .D(n272), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[18]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[19]  ( .D(\DataP/b_out[19] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[19] ), .QN(n271) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[19]  ( .D(n271), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[19]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[20]  ( .D(\DataP/b_out[20] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[20] ), .QN(n270) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[20]  ( .D(n270), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[20]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[21]  ( .D(\DataP/b_out[21] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[21] ), .QN(n269) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[21]  ( .D(n269), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[21]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[22]  ( .D(\DataP/b_out[22] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[22] ), .QN(n268) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[22]  ( .D(n268), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[22]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[23]  ( .D(\DataP/b_out[23] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[23] ), .QN(n267) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[23]  ( .D(n267), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[23]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[24]  ( .D(\DataP/b_out[24] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[24] ), .QN(n266) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[24]  ( .D(n266), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[24]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[25]  ( .D(\DataP/b_out[25] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[25] ), .QN(n265) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[25]  ( .D(n265), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[25]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[26]  ( .D(\DataP/b_out[26] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[26] ), .QN(n264) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[26]  ( .D(n264), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[26]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[27]  ( .D(\DataP/b_out[27] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[27] ), .QN(n263) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[27]  ( .D(n263), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[27]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[28]  ( .D(\DataP/b_out[28] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[28] ), .QN(n262) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[28]  ( .D(n262), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[28]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[29]  ( .D(\DataP/b_out[29] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[29] ), .QN(n261) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[29]  ( .D(n261), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[29]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[30]  ( .D(\DataP/b_out[30] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[30] ), .QN(n260) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[30]  ( .D(n260), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[30]) );
  DFFR_X1 \DataP/ID_EXs/B_OUT_reg[31]  ( .D(\DataP/b_out[31] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/B_s[31] ), .QN(n259) );
  DFFS_X1 \DataP/EX_MEM_s/B_OUT_reg[31]  ( .D(n259), .CK(Clk), .SN(Rst), .QN(
        DRAM_DATA_IN[31]) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[0]  ( .D(\DataP/a_out[0] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[0] ), .QN(n2214) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[1]  ( .D(\DataP/a_out[1] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[1] ), .QN(n2215) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[2]  ( .D(\DataP/a_out[2] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[2] ), .QN(n2213) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[3]  ( .D(\DataP/a_out[3] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[3] ), .QN(n2212) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[4]  ( .D(\DataP/a_out[4] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[4] ), .QN(n2221) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[5]  ( .D(\DataP/a_out[5] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[5] ), .QN(n2198) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[6]  ( .D(\DataP/a_out[6] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[6] ), .QN(n2216) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[7]  ( .D(\DataP/a_out[7] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[7] ), .QN(n2205) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[8]  ( .D(\DataP/a_out[8] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[8] ), .QN(n2220) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[9]  ( .D(\DataP/a_out[9] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[9] ), .QN(n2190) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[10]  ( .D(\DataP/a_out[10] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[10] ), .QN(n2211) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[11]  ( .D(\DataP/a_out[11] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[11] ), .QN(n2204) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[12]  ( .D(\DataP/a_out[12] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[12] ), .QN(n2197) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[13]  ( .D(\DataP/a_out[13] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[13] ), .QN(n2210) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[14]  ( .D(\DataP/a_out[14] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[14] ), .QN(n2203) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[15]  ( .D(\DataP/a_out[15] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[15] ), .QN(n2196) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[16]  ( .D(\DataP/a_out[16] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[16] ), .QN(n2219) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[17]  ( .D(\DataP/a_out[17] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[17] ), .QN(n2195) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[18]  ( .D(\DataP/a_out[18] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[18] ), .QN(n2209) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[19]  ( .D(\DataP/a_out[19] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[19] ), .QN(n2202) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[20]  ( .D(\DataP/a_out[20] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[20] ), .QN(n2208) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[21]  ( .D(\DataP/a_out[21] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[21] ), .QN(n2201) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[22]  ( .D(\DataP/a_out[22] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[22] ), .QN(n2218) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[23]  ( .D(\DataP/a_out[23] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[23] ), .QN(n2194) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[24]  ( .D(\DataP/a_out[24] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[24] ), .QN(n2217) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[25]  ( .D(\DataP/a_out[25] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[25] ), .QN(n2207) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[26]  ( .D(\DataP/a_out[26] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[26] ), .QN(n2200) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[27]  ( .D(\DataP/a_out[27] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[27] ), .QN(n2193) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[28]  ( .D(\DataP/a_out[28] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[28] ), .QN(n2206) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[29]  ( .D(\DataP/a_out[29] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[29] ), .QN(n2199) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[30]  ( .D(\DataP/a_out[30] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[30] ), .QN(n2192) );
  DFFR_X1 \DataP/ID_EXs/A_OUT_reg[31]  ( .D(\DataP/a_out[31] ), .CK(Clk), .RN(
        Rst), .Q(\DataP/A_s[31] ), .QN(n2191) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[0]  ( .D(n296), .CK(Clk), .SN(Rst), .Q(
        n2234), .QN(DRAM_ADDRESS[0]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[0]  ( .D(DRAM_ADDRESS[0]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[0] ), .QN(n2272) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[7]  ( .D(n350), .CK(Clk), .SN(Rst), .Q(
        n2230), .QN(DRAM_ADDRESS[7]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[7]  ( .D(DRAM_ADDRESS[7]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[7] ), .QN(n2275) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[15]  ( .D(\DataP/alu_out_M[15] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[15] ), .QN(n2247) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[19]  ( .D(\DataP/alu_out_M[19] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[19] ), .QN(n2253) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[23]  ( .D(\DataP/alu_out_M[23] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[23] ), .QN(n2249) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[27]  ( .D(n301), .CK(Clk), .SN(Rst), .Q(
        n2165), .QN(\DataP/alu_out_M[27] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[27]  ( .D(\DataP/alu_out_M[27] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[27] ), .QN(n2250) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[30]  ( .D(\DataP/alu_out_M[30] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[30] ), .QN(n2266) );
  DFFS_X1 \DataP/ID_EXs/PR_OUT_reg  ( .D(n258), .CK(Clk), .SN(Rst), .QN(
        \DataP/pr_E ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[30]  ( .D(\DataP/link_addr_F[30] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n257) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[30]  ( .D(n257), .CK(Clk), .SN(Rst), .Q(
        n256) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[30]  ( .D(n256), .CK(Clk), .SN(Rst), 
        .Q(n255) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[30]  ( .D(n255), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[30] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[29]  ( .D(\DataP/link_addr_F[29] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n254) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[29]  ( .D(n254), .CK(Clk), .SN(Rst), .Q(
        n253) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[29]  ( .D(n253), .CK(Clk), .SN(Rst), 
        .Q(n252) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[29]  ( .D(n252), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[29] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[28]  ( .D(\DataP/link_addr_F[28] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n251) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[28]  ( .D(n251), .CK(Clk), .SN(Rst), .Q(
        n250) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[28]  ( .D(n250), .CK(Clk), .SN(Rst), 
        .Q(n249) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[28]  ( .D(n249), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[28] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[27]  ( .D(\DataP/link_addr_F[27] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n248) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[27]  ( .D(n248), .CK(Clk), .SN(Rst), .Q(
        n247) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[27]  ( .D(n247), .CK(Clk), .SN(Rst), 
        .Q(n246) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[27]  ( .D(n246), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[27] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[26]  ( .D(\DataP/link_addr_F[26] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n245) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[26]  ( .D(n245), .CK(Clk), .SN(Rst), .Q(
        n244) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[26]  ( .D(n244), .CK(Clk), .SN(Rst), 
        .Q(n243) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[26]  ( .D(n243), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[26] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[25]  ( .D(\DataP/link_addr_F[25] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n242) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[25]  ( .D(n242), .CK(Clk), .SN(Rst), .Q(
        n241) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[25]  ( .D(n241), .CK(Clk), .SN(Rst), 
        .Q(n240) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[25]  ( .D(n240), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[25] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[24]  ( .D(\DataP/link_addr_F[24] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n239) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[24]  ( .D(n239), .CK(Clk), .SN(Rst), .Q(
        n238) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[24]  ( .D(n238), .CK(Clk), .SN(Rst), 
        .Q(n237) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[24]  ( .D(n237), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[24] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[23]  ( .D(\DataP/link_addr_F[23] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n236) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[23]  ( .D(n236), .CK(Clk), .SN(Rst), .Q(
        n235) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[23]  ( .D(n235), .CK(Clk), .SN(Rst), 
        .Q(n234) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[23]  ( .D(n234), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[23] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[22]  ( .D(\DataP/link_addr_F[22] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n233) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[22]  ( .D(n233), .CK(Clk), .SN(Rst), .Q(
        n232) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[22]  ( .D(n232), .CK(Clk), .SN(Rst), 
        .Q(n231) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[22]  ( .D(n231), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[22] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[21]  ( .D(\DataP/link_addr_F[21] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n230) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[21]  ( .D(n230), .CK(Clk), .SN(Rst), .Q(
        n229) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[21]  ( .D(n229), .CK(Clk), .SN(Rst), 
        .Q(n228) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[21]  ( .D(n228), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[21] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[20]  ( .D(\DataP/link_addr_F[20] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n227) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[20]  ( .D(n227), .CK(Clk), .SN(Rst), .Q(
        n226) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[20]  ( .D(n226), .CK(Clk), .SN(Rst), 
        .Q(n225) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[20]  ( .D(n225), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[20] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[19]  ( .D(\DataP/link_addr_F[19] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n224) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[19]  ( .D(n224), .CK(Clk), .SN(Rst), .Q(
        n223) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[19]  ( .D(n223), .CK(Clk), .SN(Rst), 
        .Q(n222) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[19]  ( .D(n222), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[19] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[18]  ( .D(\DataP/link_addr_F[18] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n221) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[18]  ( .D(n221), .CK(Clk), .SN(Rst), .Q(
        n220) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[18]  ( .D(n220), .CK(Clk), .SN(Rst), 
        .Q(n219) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[18]  ( .D(n219), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[18] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[17]  ( .D(\DataP/link_addr_F[17] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n218) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[17]  ( .D(n218), .CK(Clk), .SN(Rst), .Q(
        n217) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[17]  ( .D(n217), .CK(Clk), .SN(Rst), 
        .Q(n216) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[17]  ( .D(n216), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[17] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[16]  ( .D(\DataP/link_addr_F[16] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n215) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[16]  ( .D(n215), .CK(Clk), .SN(Rst), .Q(
        n214) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[16]  ( .D(n214), .CK(Clk), .SN(Rst), 
        .Q(n213) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[16]  ( .D(n213), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[16] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[15]  ( .D(\DataP/link_addr_F[15] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n212) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[15]  ( .D(n212), .CK(Clk), .SN(Rst), .Q(
        n211) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[15]  ( .D(n211), .CK(Clk), .SN(Rst), 
        .Q(n210) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[15]  ( .D(n210), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[15] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[14]  ( .D(\DataP/link_addr_F[14] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n209) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[14]  ( .D(n209), .CK(Clk), .SN(Rst), .Q(
        n208) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[14]  ( .D(n208), .CK(Clk), .SN(Rst), 
        .Q(n207) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[14]  ( .D(n207), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[14] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[13]  ( .D(\DataP/link_addr_F[13] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n206) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[13]  ( .D(n206), .CK(Clk), .SN(Rst), .Q(
        n205) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[13]  ( .D(n205), .CK(Clk), .SN(Rst), 
        .Q(n204) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[13]  ( .D(n204), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[13] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[12]  ( .D(\DataP/link_addr_F[12] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n203) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[12]  ( .D(n203), .CK(Clk), .SN(Rst), .Q(
        n202) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[12]  ( .D(n202), .CK(Clk), .SN(Rst), 
        .Q(n201) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[12]  ( .D(n201), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[12] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[11]  ( .D(\DataP/link_addr_F[11] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n200) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[11]  ( .D(n200), .CK(Clk), .SN(Rst), .Q(
        n199) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[11]  ( .D(n199), .CK(Clk), .SN(Rst), 
        .Q(n198) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[11]  ( .D(n198), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[11] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[10]  ( .D(\DataP/link_addr_F[10] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n197) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[10]  ( .D(n197), .CK(Clk), .SN(Rst), .Q(
        n196) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[10]  ( .D(n196), .CK(Clk), .SN(Rst), 
        .Q(n195) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[10]  ( .D(n195), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[10] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[9]  ( .D(\DataP/link_addr_F[9] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n194) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[9]  ( .D(n194), .CK(Clk), .SN(Rst), .Q(
        n193) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[9]  ( .D(n193), .CK(Clk), .SN(Rst), 
        .Q(n192) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[9]  ( .D(n192), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[9] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[8]  ( .D(\DataP/link_addr_F[8] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n191) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[8]  ( .D(n191), .CK(Clk), .SN(Rst), .Q(
        n190) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[8]  ( .D(n190), .CK(Clk), .SN(Rst), 
        .Q(n189) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[8]  ( .D(n189), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[8] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[7]  ( .D(\DataP/link_addr_F[7] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n188) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[7]  ( .D(n188), .CK(Clk), .SN(Rst), .Q(
        n187) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[7]  ( .D(n187), .CK(Clk), .SN(Rst), 
        .Q(n186) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[7]  ( .D(n186), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[7] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[6]  ( .D(\DataP/link_addr_F[6] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n185) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[6]  ( .D(n185), .CK(Clk), .SN(Rst), .Q(
        n184) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[6]  ( .D(n184), .CK(Clk), .SN(Rst), 
        .Q(n183) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[6]  ( .D(n183), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[6] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[5]  ( .D(\DataP/link_addr_F[5] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n182) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[5]  ( .D(n182), .CK(Clk), .SN(Rst), .Q(
        n181) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[5]  ( .D(n181), .CK(Clk), .SN(Rst), 
        .Q(n180) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[5]  ( .D(n180), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[5] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[4]  ( .D(\DataP/link_addr_F[4] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n179) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[4]  ( .D(n179), .CK(Clk), .SN(Rst), .Q(
        n178) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[4]  ( .D(n178), .CK(Clk), .SN(Rst), 
        .Q(n177) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[4]  ( .D(n177), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[4] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[3]  ( .D(\DataP/link_addr_F[3] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n176) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[3]  ( .D(n176), .CK(Clk), .SN(Rst), .Q(
        n175) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[3]  ( .D(n175), .CK(Clk), .SN(Rst), 
        .Q(n174) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[3]  ( .D(n174), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[3] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[2]  ( .D(\DataP/link_addr_F[2] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n173) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[2]  ( .D(n173), .CK(Clk), .SN(Rst), .Q(
        n172) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[2]  ( .D(n172), .CK(Clk), .SN(Rst), 
        .Q(n171) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[2]  ( .D(n171), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[2] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[1]  ( .D(\DataP/link_addr_F[1] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n170) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[1]  ( .D(n170), .CK(Clk), .SN(Rst), .Q(
        n169) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[1]  ( .D(n169), .CK(Clk), .SN(Rst), 
        .Q(n168) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[1]  ( .D(n168), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[1] ) );
  DFFR_X1 \DataP/IF_IDs/NPC_L_OUT_reg[0]  ( .D(\DataP/link_addr_F[0] ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n167) );
  DFFS_X1 \DataP/ID_EXs/NPC_L_OUT_reg[0]  ( .D(n167), .CK(Clk), .SN(Rst), .Q(
        n166) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_L_OUT_reg[0]  ( .D(n166), .CK(Clk), .SN(Rst), 
        .Q(n165) );
  DFFS_X1 \DataP/MEM_WB_s/NPC_L_OUT_reg[0]  ( .D(n165), .CK(Clk), .SN(Rst), 
        .QN(\DataP/link_addr_W[0] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[0]  ( .D(IRAM_DATA_OUT[0]), .CK(Clk), .RN(
        n164), .Q(IR_CU[0]), .QN(n476) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[0]  ( .D(n476), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[0] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[1]  ( .D(IRAM_DATA_OUT[1]), .CK(Clk), .RN(
        n164), .Q(IR_CU[1]), .QN(n477) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[1]  ( .D(n477), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[1] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[2]  ( .D(IRAM_DATA_OUT[2]), .CK(Clk), .RN(
        n164), .Q(n2128), .QN(n478) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[2]  ( .D(n478), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[2] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[3]  ( .D(IRAM_DATA_OUT[3]), .CK(Clk), .RN(
        n164), .Q(n2135), .QN(n479) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[3]  ( .D(n479), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[3] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[4]  ( .D(IRAM_DATA_OUT[4]), .CK(Clk), .RN(
        n164), .Q(IR_CU[4]), .QN(n480) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[4]  ( .D(n480), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[4] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[5]  ( .D(IRAM_DATA_OUT[5]), .CK(Clk), .RN(
        n164), .Q(IR_CU[5]), .QN(n482) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[5]  ( .D(n482), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[5] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[6]  ( .D(IRAM_DATA_OUT[6]), .CK(Clk), .RN(
        n164), .Q(IR_CU[6]), .QN(n163) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[6]  ( .D(n163), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[6] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[7]  ( .D(IRAM_DATA_OUT[7]), .CK(Clk), .RN(
        n164), .Q(IR_CU[7]), .QN(n162) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[7]  ( .D(n162), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[7] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[8]  ( .D(IRAM_DATA_OUT[8]), .CK(Clk), .RN(
        n164), .Q(IR_CU[8]), .QN(n161) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[8]  ( .D(n161), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[8] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[9]  ( .D(IRAM_DATA_OUT[9]), .CK(Clk), .RN(
        n164), .Q(IR_CU[9]), .QN(n160) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[9]  ( .D(n160), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[9] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[10]  ( .D(IRAM_DATA_OUT[10]), .CK(Clk), 
        .RN(n164), .QN(n484) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[10]  ( .D(n484), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[10] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[11]  ( .D(IRAM_DATA_OUT[11]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[11] ), .QN(n159) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[11]  ( .D(n159), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[11] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[12]  ( .D(IRAM_DATA_OUT[12]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[12] ), .QN(n158) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[12]  ( .D(n158), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[12] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[13]  ( .D(IRAM_DATA_OUT[13]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[13] ), .QN(n157) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[13]  ( .D(n157), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[13] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[14]  ( .D(IRAM_DATA_OUT[14]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[14] ), .QN(n156) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[14]  ( .D(n156), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[14] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[15]  ( .D(IRAM_DATA_OUT[15]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[15] ), .QN(n155) );
  DFFS_X1 \DataP/ID_EXs/IR_OUT_reg[15]  ( .D(n155), .CK(Clk), .SN(Rst), .QN(
        \DataP/ir_E[15] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[16]  ( .D(IRAM_DATA_OUT[16]), .CK(Clk), 
        .RN(n164), .QN(n485) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[17]  ( .D(IRAM_DATA_OUT[17]), .CK(Clk), 
        .RN(n164), .QN(n486) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[18]  ( .D(IRAM_DATA_OUT[18]), .CK(Clk), 
        .RN(n164), .QN(n487) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[19]  ( .D(IRAM_DATA_OUT[19]), .CK(Clk), 
        .RN(n164), .QN(n488) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[20]  ( .D(IRAM_DATA_OUT[20]), .CK(Clk), 
        .RN(n164), .QN(n489) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[21]  ( .D(IRAM_DATA_OUT[21]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[21] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[22]  ( .D(IRAM_DATA_OUT[22]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[22] ), .QN(n153) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[23]  ( .D(IRAM_DATA_OUT[23]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[23] ), .QN(n152) );
  DFFS_X1 \DataP/ID_EXs/RS1_OUT_reg[2]  ( .D(n152), .CK(Clk), .SN(Rst), .Q(
        n2156), .QN(\DataP/Rs1[2] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[24]  ( .D(IRAM_DATA_OUT[24]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[24] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[25]  ( .D(IRAM_DATA_OUT[25]), .CK(Clk), 
        .RN(n164), .Q(\DataP/IR1[25] ) );
  DFFR_X1 \DataP/ID_EXs/RS1_OUT_reg[4]  ( .D(\DataP/IR1[25] ), .CK(Clk), .RN(
        Rst), .QN(n524) );
  DFFS_X1 \DataP/IF_IDs/IR_OUT_reg[26]  ( .D(IRAM_DATA_OUT[26]), .CK(Clk), 
        .SN(n164), .Q(IR_CU_26), .QN(n497) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[0]  ( .D(n150), .CK(Clk), .SN(Rst), 
        .Q(n2162), .QN(\DataP/opcode_W[0] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[27]  ( .D(IRAM_DATA_OUT[27]), .CK(Clk), 
        .RN(n164), .Q(IR_CU_27), .QN(n504) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[1]  ( .D(n520), .CK(Clk), .SN(Rst), 
        .Q(n2576), .QN(\DataP/opcode_M[1] ) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[2]  ( .D(n510), .CK(Clk), .SN(Rst), .Q(
        n521), .QN(n2574) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[29]  ( .D(IRAM_DATA_OUT[29]), .CK(Clk), 
        .RN(n164), .Q(n2141), .QN(n514) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[3]  ( .D(n514), .CK(Clk), .SN(Rst), .Q(
        n149), .QN(\DataP/opcode_E[3] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[3]  ( .D(n149), .CK(Clk), .SN(Rst), 
        .Q(n148), .QN(\DataP/opcode_M[3] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[3]  ( .D(n148), .CK(Clk), .SN(Rst), 
        .Q(n2159), .QN(\DataP/opcode_W[3] ) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[4]  ( .D(n515), .CK(Clk), .SN(Rst), .Q(
        n147), .QN(\DataP/opcode_E[4] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[4]  ( .D(n146), .CK(Clk), .SN(Rst), 
        .Q(n2151), .QN(\DataP/opcode_W[4] ) );
  DFFR_X1 \DataP/IF_IDs/IR_OUT_reg[31]  ( .D(IRAM_DATA_OUT[31]), .CK(Clk), 
        .RN(n164), .Q(IR_CU_31), .QN(n516) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[5]  ( .D(n516), .CK(Clk), .SN(Rst), .Q(
        n145) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[5]  ( .D(n145), .CK(Clk), .SN(Rst), 
        .Q(n2161), .QN(\DataP/opcode_M[5] ) );
  DLH_X1 \DataP/FORWARDING_BR/SEL_reg[1]  ( .G(\DataP/FORWARDING_BR/N12 ), .D(
        n3710), .Q(\DataP/FWD_MUX_BR_S[1] ) );
  SDFFR_X1 \CU_I/cw1_reg[8]  ( .D(n144), .SI(n606), .SE(n504), .CK(Clk), .RN(
        Rst), .Q(BR_EN_i) );
  DFFR_X1 \CU_I/aluOpcode1_reg[3]  ( .D(\CU_I/aluOpcode_i[3] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[3]), .QN(n2146) );
  DFFR_X1 \CU_I/cw1_reg[10]  ( .D(\CU_I/cw[10] ), .CK(Clk), .RN(Rst), .Q(n2155), .QN(n432) );
  DFFS_X1 \CU_I/cw2_reg[7]  ( .D(n143), .CK(Clk), .SN(Rst), .QN(DRAM_RW) );
  DFFR_X1 \DataP/ID_EXs/RS2_OUT_reg[2]  ( .D(\DataP/add_S2[2] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/Rs2[2] ) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[4]  ( .D(n142), .CK(Clk), .SN(Rst), .Q(
        n2569), .QN(\DataP/dest_M[4] ) );
  DFFR_X1 \DataP/MEM_WB_s/RD_OUT_reg[4]  ( .D(\DataP/dest_M[4] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/add_D[4] ), .QN(n540) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[3]  ( .D(n141), .CK(Clk), .SN(Rst), .Q(
        n2570), .QN(\DataP/dest_M[3] ) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[2]  ( .D(n140), .CK(Clk), .SN(Rst), .Q(
        n530), .QN(\DataP/dest_M[2] ) );
  DFFS_X1 \DataP/EX_MEM_s/RD_OUT_reg[1]  ( .D(n139), .CK(Clk), .SN(Rst), .Q(
        n529), .QN(\DataP/dest_M[1] ) );
  DFFR_X1 \DataP/MEM_WB_s/RD_OUT_reg[0]  ( .D(\DataP/dest_M[0] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/add_D[0] ), .QN(n536) );
  DLH_X1 \DataP/FORWARDING_BR/SEL_reg[0]  ( .G(\DataP/FORWARDING_BR/N12 ), .D(
        n2469), .Q(\DataP/FWD_MUX_BR_S[0] ) );
  DFFR_X1 \CU_I/aluOpcode1_reg[0]  ( .D(\CU_I/aluOpcode_i[0] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[0]), .QN(n2150) );
  DFFR_X1 \CU_I/aluOpcode1_reg[4]  ( .D(\CU_I/aluOpcode_i[4] ), .CK(Clk), .RN(
        Rst), .Q(n2134), .QN(n443) );
  DFFR_X1 \CU_I/aluOpcode1_reg[2]  ( .D(\CU_I/aluOpcode_i[2] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[2]), .QN(n2144) );
  DFFR_X1 \CU_I/aluOpcode1_reg[1]  ( .D(\CU_I/aluOpcode_i[1] ), .CK(Clk), .RN(
        Rst), .Q(ALU_OPCODE_i[1]), .QN(n2132) );
  DFFS_X1 \CU_I/cw1_reg[5]  ( .D(n1357), .CK(Clk), .SN(Rst), .Q(n137) );
  DFFS_X1 \CU_I/cw2_reg[5]  ( .D(n137), .CK(Clk), .SN(Rst), .QN(DRAM_SEL[2])
         );
  DFFS_X1 \CU_I/cw2_reg[0]  ( .D(n136), .CK(Clk), .SN(Rst), .Q(n135) );
  DFFS_X1 \CU_I/cw3_reg[0]  ( .D(n135), .CK(Clk), .SN(Rst), .QN(RF_WE_i) );
  DFFS_X1 \CU_I/cw1_reg[2]  ( .D(n1371), .CK(Clk), .SN(Rst), .Q(n134) );
  DFFS_X1 \CU_I/cw2_reg[2]  ( .D(n134), .CK(Clk), .SN(Rst), .Q(n133) );
  DFFS_X1 \CU_I/cw3_reg[2]  ( .D(n133), .CK(Clk), .SN(Rst), .QN(
        \WB_MUX_SEL_i[1] ) );
  DFFS_X1 \CU_I/cw2_reg[4]  ( .D(n132), .CK(Clk), .SN(Rst), .QN(DRAM_SEL[1])
         );
  DFFS_X1 \CU_I/cw2_reg[3]  ( .D(n131), .CK(Clk), .SN(Rst), .QN(DRAM_SEL[0])
         );
  DFFS_X1 \CU_I/cw2_reg[6]  ( .D(n130), .CK(Clk), .SN(Rst), .QN(DRAM_ENABLE)
         );
  DFFR_X1 \CU_I/cw1_reg[9]  ( .D(\CU_I/cw[9] ), .CK(Clk), .RN(Rst), .Q(n2189), 
        .QN(n399) );
  DFFS_X1 \CU_I/cw2_reg[1]  ( .D(n129), .CK(Clk), .SN(Rst), .QN(\CU_I/cw2[1] )
         );
  DFFR_X1 \CU_I/cw3_reg[1]  ( .D(\CU_I/cw2[1] ), .CK(Clk), .RN(Rst), .QN(n294)
         );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[31]  ( .D(\DataP/imm_out[31] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[31] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[24]  ( .D(\DataP/imm_out[24] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[24] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[23]  ( .D(\DataP/imm_out[23] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[23] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[22]  ( .D(\DataP/imm_out[22] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[22] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[21]  ( .D(\DataP/imm_out[21] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[21] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[20]  ( .D(\DataP/imm_out[20] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[20] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[19]  ( .D(\DataP/imm_out[19] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[19] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[18]  ( .D(\DataP/imm_out[18] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[18] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[17]  ( .D(\DataP/imm_out[17] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[17] ) );
  DFFR_X1 \DataP/ID_EXs/IMM_OUT_reg[16]  ( .D(\DataP/imm_out[16] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/IMM_s[16] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[0]  ( .D(\DataP/npc[0] ), .CK(Clk), .RN(
        n126), .SN(n127), .QN(n128) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[0]  ( .D(n128), .CK(Clk), .SN(Rst), .Q(
        n125) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[0]  ( .D(n125), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[0] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[1]  ( .D(\DataP/npc[1] ), .CK(Clk), .RN(
        n122), .SN(n123), .QN(n124) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[1]  ( .D(n124), .CK(Clk), .SN(Rst), .Q(
        n121) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[1]  ( .D(n121), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[1] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[1]  ( .D(n358), .CK(Clk), .SN(Rst), .Q(
        n2233), .QN(DRAM_ADDRESS[1]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[1]  ( .D(DRAM_ADDRESS[1]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[1] ), .QN(n2273) );
  DFF_X1 \DataP/PC_reg/O_reg[1]  ( .D(\DataP/PC_reg/N3 ), .CK(Clk), .Q(
        \DataP/pc_out_1 ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[2]  ( .D(\DataP/npc[2] ), .CK(Clk), .RN(
        n118), .SN(n119), .QN(n120) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[2]  ( .D(n120), .CK(Clk), .SN(Rst), .Q(
        n117) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[2]  ( .D(n117), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[2] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[2]  ( .D(n357), .CK(Clk), .SN(Rst), .Q(
        n2232), .QN(DRAM_ADDRESS[2]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[2]  ( .D(DRAM_ADDRESS[2]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[2] ), .QN(n2276) );
  DFF_X1 \DataP/PC_reg/O_reg[2]  ( .D(\DataP/PC_reg/N4 ), .CK(Clk), .Q(
        IRAM_ADDRESS[0]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[3]  ( .D(\DataP/npc[3] ), .CK(Clk), .RN(
        n114), .SN(n115), .QN(n116) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[3]  ( .D(n116), .CK(Clk), .SN(Rst), .Q(
        n113) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[3]  ( .D(n113), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[3] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[3]  ( .D(n356), .CK(Clk), .SN(Rst), .Q(
        n2231), .QN(DRAM_ADDRESS[3]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[3]  ( .D(DRAM_ADDRESS[3]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[3] ), .QN(n2277) );
  DFF_X1 \DataP/PC_reg/O_reg[3]  ( .D(\DataP/PC_reg/N5 ), .CK(Clk), .Q(
        IRAM_ADDRESS[1]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[4]  ( .D(\DataP/npc[4] ), .CK(Clk), .RN(
        n110), .SN(n111), .QN(n112) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[4]  ( .D(n112), .CK(Clk), .SN(Rst), .Q(
        n109) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[4]  ( .D(n109), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[4] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[4]  ( .D(n355), .CK(Clk), .SN(Rst), .Q(
        n2229), .QN(DRAM_ADDRESS[4]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[4]  ( .D(DRAM_ADDRESS[4]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[4] ), .QN(n2274) );
  DFF_X1 \DataP/PC_reg/O_reg[4]  ( .D(\DataP/PC_reg/N6 ), .CK(Clk), .Q(
        IRAM_ADDRESS[2]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[5]  ( .D(\DataP/npc[5] ), .CK(Clk), .RN(
        n106), .SN(n107), .QN(n108) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[5]  ( .D(n108), .CK(Clk), .SN(Rst), .Q(
        n105) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[5]  ( .D(n105), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[5] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[5]  ( .D(n354), .CK(Clk), .SN(Rst), .Q(
        n2227), .QN(DRAM_ADDRESS[5]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[5]  ( .D(DRAM_ADDRESS[5]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[5] ), .QN(n2270) );
  DFF_X1 \DataP/PC_reg/O_reg[5]  ( .D(\DataP/PC_reg/N7 ), .CK(Clk), .Q(
        IRAM_ADDRESS[3]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[6]  ( .D(\DataP/npc[6] ), .CK(Clk), .RN(
        n102), .SN(n103), .QN(n104) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[6]  ( .D(n104), .CK(Clk), .SN(Rst), .Q(
        n101) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[6]  ( .D(n101), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[6] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[6]  ( .D(n353), .CK(Clk), .SN(Rst), .Q(
        n2182), .QN(DRAM_ADDRESS[6]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[6]  ( .D(DRAM_ADDRESS[6]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[6] ), .QN(n2268) );
  DFF_X1 \DataP/PC_reg/O_reg[6]  ( .D(\DataP/PC_reg/N8 ), .CK(Clk), .Q(
        IRAM_ADDRESS[4]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[7]  ( .D(\DataP/npc[7] ), .CK(Clk), .RN(
        n98), .SN(n99), .QN(n100) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[7]  ( .D(n100), .CK(Clk), .SN(Rst), .Q(n97) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[7]  ( .D(n97), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[7] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[8]  ( .D(\DataP/npc[8] ), .CK(Clk), .RN(
        n94), .SN(n95), .QN(n96) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[8]  ( .D(n96), .CK(Clk), .SN(Rst), .Q(n93)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[8]  ( .D(n93), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[8] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[8]  ( .D(n345), .CK(Clk), .SN(Rst), .QN(
        DRAM_ADDRESS[8]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[8]  ( .D(DRAM_ADDRESS[8]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[8] ), .QN(n2271) );
  DFF_X1 \DataP/PC_reg/O_reg[8]  ( .D(\DataP/PC_reg/N10 ), .CK(Clk), .Q(
        IRAM_ADDRESS[6]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[9]  ( .D(\DataP/npc[9] ), .CK(Clk), .RN(
        n90), .SN(n91), .QN(n92) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[9]  ( .D(n92), .CK(Clk), .SN(Rst), .Q(n89)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[9]  ( .D(n89), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[9] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[9]  ( .D(n341), .CK(Clk), .SN(Rst), .Q(
        n2228), .QN(DRAM_ADDRESS[9]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[9]  ( .D(DRAM_ADDRESS[9]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[9] ), .QN(n2269) );
  DFF_X1 \DataP/PC_reg/O_reg[9]  ( .D(\DataP/PC_reg/N11 ), .CK(Clk), .Q(
        IRAM_ADDRESS[7]) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[10]  ( .D(\DataP/npc[10] ), .CK(Clk), 
        .RN(n86), .SN(n87), .QN(n88) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[10]  ( .D(n88), .CK(Clk), .SN(Rst), .Q(n85) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[10]  ( .D(n85), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[10] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[10]  ( .D(n340), .CK(Clk), .SN(Rst), 
        .QN(DRAM_ADDRESS[10]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[10]  ( .D(DRAM_ADDRESS[10]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[10] ), .QN(n2257) );
  DFF_X1 \DataP/PC_reg/O_reg[10]  ( .D(\DataP/PC_reg/N12 ), .CK(Clk), .Q(
        \DataP/pc_out[10] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[11]  ( .D(\DataP/npc[11] ), .CK(Clk), 
        .RN(n82), .SN(n83), .QN(n84) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[11]  ( .D(n84), .CK(Clk), .SN(Rst), .Q(n81) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[11]  ( .D(n81), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[11] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[11]  ( .D(n2137), .CK(Clk), .SN(Rst), 
        .Q(n2164), .QN(DRAM_ADDRESS[11]) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[11]  ( .D(DRAM_ADDRESS[11]), .CK(Clk), 
        .RN(Rst), .Q(\DataP/alu_out_W[11] ), .QN(n2251) );
  DFF_X1 \DataP/PC_reg/O_reg[11]  ( .D(\DataP/PC_reg/N13 ), .CK(Clk), .Q(
        \DataP/pc_out[11] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[12]  ( .D(\DataP/npc[12] ), .CK(Clk), 
        .RN(n78), .SN(n79), .QN(n80) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[12]  ( .D(n80), .CK(Clk), .SN(Rst), .Q(n77) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[12]  ( .D(n77), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[12] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[12]  ( .D(n337), .CK(Clk), .SN(Rst), .Q(
        n2177), .QN(\DataP/alu_out_M[12] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[12]  ( .D(\DataP/alu_out_M[12] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[12] ), .QN(n2246) );
  DFF_X1 \DataP/PC_reg/O_reg[12]  ( .D(\DataP/PC_reg/N14 ), .CK(Clk), .Q(
        \DataP/pc_out[12] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[13]  ( .D(\DataP/npc[13] ), .CK(Clk), 
        .RN(n74), .SN(n75), .QN(n76) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[13]  ( .D(n76), .CK(Clk), .SN(Rst), .Q(n73) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[13]  ( .D(n73), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[13] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[13]  ( .D(n333), .CK(Clk), .SN(Rst), .Q(
        n2176), .QN(\DataP/alu_out_M[13] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[13]  ( .D(\DataP/alu_out_M[13] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[13] ), .QN(n2258) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[14]  ( .D(\DataP/npc[14] ), .CK(Clk), 
        .RN(n70), .SN(n71), .QN(n72) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[14]  ( .D(n72), .CK(Clk), .SN(Rst), .Q(n69) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[14]  ( .D(n69), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[14] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[14]  ( .D(n332), .CK(Clk), .SN(Rst), .Q(
        n2171), .QN(\DataP/alu_out_M[14] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[14]  ( .D(\DataP/alu_out_M[14] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[14] ), .QN(n2252) );
  DFF_X1 \DataP/PC_reg/O_reg[14]  ( .D(\DataP/PC_reg/N16 ), .CK(Clk), .Q(
        \DataP/pc_out[14] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[15]  ( .D(\DataP/npc[15] ), .CK(Clk), 
        .RN(n66), .SN(n67), .QN(n68) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[15]  ( .D(n68), .CK(Clk), .SN(Rst), .Q(n65) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[15]  ( .D(n65), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[15] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[16]  ( .D(\DataP/npc[16] ), .CK(Clk), 
        .RN(n62), .SN(n63), .QN(n64) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[16]  ( .D(n64), .CK(Clk), .SN(Rst), .Q(n61) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[16]  ( .D(n61), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[16] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[16]  ( .D(n326), .CK(Clk), .SN(Rst), .Q(
        n2167), .QN(\DataP/alu_out_M[16] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[16]  ( .D(\DataP/alu_out_M[16] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[16] ), .QN(n2263) );
  DFF_X1 \DataP/PC_reg/O_reg[16]  ( .D(\DataP/PC_reg/N18 ), .CK(Clk), .Q(
        \DataP/pc_out[16] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[17]  ( .D(\DataP/npc[17] ), .CK(Clk), 
        .RN(n58), .SN(n59), .QN(n60) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[17]  ( .D(n60), .CK(Clk), .SN(Rst), .Q(n57) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[17]  ( .D(n57), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[17] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[17]  ( .D(\DataP/alu_out_M[17] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[17] ), .QN(n2248) );
  DFF_X1 \DataP/PC_reg/O_reg[17]  ( .D(\DataP/PC_reg/N19 ), .CK(Clk), .Q(
        \DataP/pc_out[17] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[18]  ( .D(\DataP/npc[18] ), .CK(Clk), 
        .RN(n54), .SN(n55), .QN(n56) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[18]  ( .D(n56), .CK(Clk), .SN(Rst), .Q(n53) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[18]  ( .D(n53), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[18] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[18]  ( .D(n322), .CK(Clk), .SN(Rst), 
        .QN(\DataP/alu_out_M[18] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[18]  ( .D(\DataP/alu_out_M[18] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[18] ), .QN(n2259) );
  DFF_X1 \DataP/PC_reg/O_reg[18]  ( .D(\DataP/PC_reg/N20 ), .CK(Clk), .Q(
        \DataP/pc_out[18] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[19]  ( .D(\DataP/npc[19] ), .CK(Clk), 
        .RN(n50), .SN(n51), .QN(n52) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[19]  ( .D(n52), .CK(Clk), .SN(Rst), .Q(n49) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[19]  ( .D(n49), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[19] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[20]  ( .D(\DataP/npc[20] ), .CK(Clk), 
        .RN(n46), .SN(n47), .QN(n48) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[20]  ( .D(n48), .CK(Clk), .SN(Rst), .Q(n45) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[20]  ( .D(n45), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[20] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[20]  ( .D(n317), .CK(Clk), .SN(Rst), .Q(
        n2173), .QN(\DataP/alu_out_M[20] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[20]  ( .D(\DataP/alu_out_M[20] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[20] ), .QN(n2260) );
  DFF_X1 \DataP/PC_reg/O_reg[20]  ( .D(\DataP/PC_reg/N22 ), .CK(Clk), .Q(
        \DataP/pc_out[20] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[21]  ( .D(\DataP/npc[21] ), .CK(Clk), 
        .RN(n42), .SN(n43), .QN(n44) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[21]  ( .D(n44), .CK(Clk), .SN(Rst), .Q(n41) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[21]  ( .D(n41), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[21] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[21]  ( .D(n313), .CK(Clk), .SN(Rst), .Q(
        n2172), .QN(\DataP/alu_out_M[21] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[21]  ( .D(\DataP/alu_out_M[21] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[21] ), .QN(n2254) );
  DFF_X1 \DataP/PC_reg/O_reg[21]  ( .D(\DataP/PC_reg/N23 ), .CK(Clk), .Q(
        \DataP/pc_out[21] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[22]  ( .D(\DataP/npc[22] ), .CK(Clk), 
        .RN(n38), .SN(n39), .QN(n40) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[22]  ( .D(n40), .CK(Clk), .SN(Rst), .Q(n37) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[22]  ( .D(n37), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[22] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[22]  ( .D(\DataP/alu_out_M[22] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[22] ), .QN(n2264) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[23]  ( .D(\DataP/npc[23] ), .CK(Clk), 
        .RN(n34), .SN(n35), .QN(n36) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[23]  ( .D(n36), .CK(Clk), .SN(Rst), .Q(n33) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[23]  ( .D(n33), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[23] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[24]  ( .D(\DataP/npc[24] ), .CK(Clk), 
        .RN(n30), .SN(n31), .QN(n32) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[24]  ( .D(n32), .CK(Clk), .SN(Rst), .Q(n29) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[24]  ( .D(n29), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[24] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[24]  ( .D(n308), .CK(Clk), .SN(Rst), .Q(
        n2179), .QN(\DataP/alu_out_M[24] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[24]  ( .D(\DataP/alu_out_M[24] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[24] ), .QN(n2265) );
  DFF_X1 \DataP/PC_reg/O_reg[24]  ( .D(\DataP/PC_reg/N26 ), .CK(Clk), .Q(
        \DataP/pc_out[24] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[25]  ( .D(\DataP/npc[25] ), .CK(Clk), 
        .RN(n26), .SN(n27), .QN(n28) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[25]  ( .D(n28), .CK(Clk), .SN(Rst), .Q(n25) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[25]  ( .D(n25), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[25] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[25]  ( .D(n304), .CK(Clk), .SN(Rst), .Q(
        n2175), .QN(\DataP/alu_out_M[25] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[25]  ( .D(\DataP/alu_out_M[25] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[25] ), .QN(n2261) );
  DFF_X1 \DataP/PC_reg/O_reg[25]  ( .D(\DataP/PC_reg/N27 ), .CK(Clk), .Q(
        \DataP/pc_out[25] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[26]  ( .D(\DataP/npc[26] ), .CK(Clk), 
        .RN(n22), .SN(n23), .QN(n24) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[26]  ( .D(n24), .CK(Clk), .SN(Rst), .Q(n21) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[26]  ( .D(n21), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[26] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[26]  ( .D(\DataP/alu_out_M[26] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[26] ), .QN(n2255) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[27]  ( .D(\DataP/npc[27] ), .CK(Clk), 
        .RN(n18), .SN(n19), .QN(n20) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[27]  ( .D(n20), .CK(Clk), .SN(Rst), .Q(n17) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[27]  ( .D(n17), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[27] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[28]  ( .D(\DataP/npc[28] ), .CK(Clk), 
        .RN(n14), .SN(n15), .QN(n16) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[28]  ( .D(n16), .CK(Clk), .SN(Rst), .Q(n13) );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[28]  ( .D(n13), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[28] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[28]  ( .D(\DataP/alu_out_M[28] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[28] ), .QN(n2262) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[29]  ( .D(\DataP/npc[29] ), .CK(Clk), 
        .RN(n10), .SN(n11), .QN(n12) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[29]  ( .D(n12), .CK(Clk), .SN(Rst), .Q(n9)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[29]  ( .D(n9), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[29] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[29]  ( .D(n299), .CK(Clk), .SN(Rst), 
        .QN(\DataP/alu_out_M[29] ) );
  DFFR_X1 \DataP/MEM_WB_s/ALU_OUT_reg[29]  ( .D(\DataP/alu_out_M[29] ), .CK(
        Clk), .RN(Rst), .Q(\DataP/alu_out_W[29] ), .QN(n2256) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[30]  ( .D(\DataP/npc[30] ), .CK(Clk), 
        .RN(n6), .SN(n7), .QN(n8) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[30]  ( .D(n8), .CK(Clk), .SN(Rst), .Q(n5)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[30]  ( .D(n5), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[30] ) );
  DFFRS_X1 \DataP/IF_IDs/NPC_OUT_reg[31]  ( .D(\DataP/npc[31] ), .CK(Clk), 
        .RN(n2), .SN(n3), .QN(n4) );
  DFFS_X1 \DataP/ID_EXs/NPC_OUT_reg[31]  ( .D(n4), .CK(Clk), .SN(Rst), .Q(n1)
         );
  DFFS_X1 \DataP/EX_MEM_s/NPC_OUT_reg[31]  ( .D(n1), .CK(Clk), .SN(Rst), .QN(
        \DataP/npc_M[31] ) );
  DFF_X1 \DataP/PC_reg/O_reg[27]  ( .D(\DataP/PC_reg/N29 ), .CK(Clk), .Q(
        \DataP/pc_out[27] ) );
  DFF_X1 \DataP/PC_reg/O_reg[23]  ( .D(\DataP/PC_reg/N25 ), .CK(Clk), .Q(
        \DataP/pc_out[23] ) );
  DFF_X1 \DataP/PC_reg/O_reg[7]  ( .D(\DataP/PC_reg/N9 ), .CK(Clk), .Q(
        IRAM_ADDRESS[5]) );
  DFF_X1 \DataP/PC_reg/O_reg[0]  ( .D(\DataP/PC_reg/N2 ), .CK(Clk), .Q(
        \DataP/pc_out_0 ) );
  AOI21_X1 \sra_131/*cell*849188  ( .B1(n2065), .B2(n2929), .A(n2981), .ZN(
        n2930) );
  AOI21_X1 \sra_131/*cell*849192  ( .B1(n2065), .B2(n2925), .A(n2981), .ZN(
        n2926) );
  AOI22_X1 \sra_131/*cell*849318  ( .A1(n2713), .A2(n2857), .B1(n2860), .B2(
        n2988), .ZN(n2869) );
  AOI22_X1 \sra_131/*cell*849321  ( .A1(n2713), .A2(n2855), .B1(n2858), .B2(
        n2988), .ZN(n2866) );
  AOI22_X1 \sra_131/*cell*849322  ( .A1(n2986), .A2(\DataP/alu_a_in[21] ), 
        .B1(\DataP/alu_a_in[20] ), .B2(n2985), .ZN(n2858) );
  AOI22_X1 \sra_131/*cell*849327  ( .A1(n2986), .A2(\DataP/alu_a_in[25] ), 
        .B1(\DataP/alu_a_in[24] ), .B2(n2985), .ZN(n2856) );
  AOI22_X1 \sra_131/*cell*849328  ( .A1(n2986), .A2(\DataP/alu_a_in[27] ), 
        .B1(\DataP/alu_a_in[26] ), .B2(n2985), .ZN(n2853) );
  AOI22_X1 \sra_131/*cell*849329  ( .A1(n2839), .A2(n2852), .B1(n2854), .B2(
        n2988), .ZN(n2865) );
  AOI22_X1 \sra_131/*cell*849331  ( .A1(n2986), .A2(\DataP/alu_a_in[29] ), 
        .B1(\DataP/alu_a_in[28] ), .B2(n2985), .ZN(n2854) );
  AOI22_X1 \sra_131/*cell*849332  ( .A1(n2986), .A2(\DataP/alu_a_in[31] ), 
        .B1(\DataP/alu_a_in[30] ), .B2(n2985), .ZN(n2852) );
  AOI22_X1 \ashr_130/*cell*849337  ( .A1(n1915), .A2(n2835), .B1(n2834), .B2(
        n2845), .ZN(n2837) );
  AOI22_X1 \ashr_130/*cell*849339  ( .A1(n1915), .A2(n2831), .B1(n2830), .B2(
        n2064), .ZN(n2833) );
  AOI22_X1 \ashr_130/*cell*849345  ( .A1(n2841), .A2(n2821), .B1(n2820), .B2(
        n1930), .ZN(n2822) );
  AOI22_X1 \ashr_130/*cell*849348  ( .A1(n2841), .A2(n2816), .B1(n2815), .B2(
        n1930), .ZN(n2817) );
  AOI22_X1 \ashr_130/*cell*849350  ( .A1(n1915), .A2(n2812), .B1(n2811), .B2(
        n2127), .ZN(n2814) );
  AOI22_X1 \ashr_130/*cell*849351  ( .A1(n2842), .A2(n2810), .B1(n2809), .B2(
        n1930), .ZN(n2811) );
  AOI22_X1 \ashr_130/*cell*849356  ( .A1(\sra_131/SH[1] ), .A2(n2804), .B1(
        n2803), .B2(n1916), .ZN(n2825) );
  NOR2_X1 \ashr_130/*cell*849357  ( .A1(\lt_x_134/B[4] ), .A2(n2802), .ZN(
        \DataP/ALU_C/shifter/N81 ) );
  NOR2_X1 \ashr_130/*cell*849358  ( .A1(\lt_x_134/B[4] ), .A2(n2801), .ZN(
        \DataP/ALU_C/shifter/N80 ) );
  AOI22_X1 \ashr_130/*cell*849361  ( .A1(n2842), .A2(n2820), .B1(n2797), .B2(
        n1930), .ZN(n2798) );
  AOI22_X1 \ashr_130/*cell*849362  ( .A1(\sra_131/SH[1] ), .A2(n2796), .B1(
        n2795), .B2(n1916), .ZN(n2797) );
  AOI22_X1 \ashr_130/*cell*849363  ( .A1(\sra_131/SH[1] ), .A2(n2794), .B1(
        n2793), .B2(n1916), .ZN(n2820) );
  AND2_X1 \ashr_130/*cell*849364  ( .A1(n2792), .A2(n2847), .ZN(
        \DataP/ALU_C/shifter/N79 ) );
  NOR2_X1 \ashr_130/*cell*849365  ( .A1(\lt_x_135/B[4] ), .A2(n2791), .ZN(
        \DataP/ALU_C/shifter/N78 ) );
  AND2_X1 \ashr_130/*cell*849366  ( .A1(n2790), .A2(n2847), .ZN(
        \DataP/ALU_C/shifter/N77 ) );
  AND2_X1 \ashr_130/*cell*849367  ( .A1(n2789), .A2(n2065), .ZN(
        \DataP/ALU_C/shifter/N76 ) );
  AND2_X1 \ashr_130/*cell*849368  ( .A1(n2836), .A2(n2847), .ZN(
        \DataP/ALU_C/shifter/N75 ) );
  AOI22_X1 \ashr_130/*cell*849419  ( .A1(\sra_131/SH[1] ), .A2(n2747), .B1(
        n2746), .B2(n1916), .ZN(n2763) );
  AOI22_X1 \ashr_130/*cell*849420  ( .A1(n1915), .A2(n2779), .B1(n2818), .B2(
        n2845), .ZN(n2748) );
  AOI22_X1 \ashr_130/*cell*849421  ( .A1(n2842), .A2(n2764), .B1(n2771), .B2(
        n1930), .ZN(n2818) );
  AOI22_X1 \ashr_130/*cell*849422  ( .A1(n2839), .A2(n2745), .B1(n2744), .B2(
        n1916), .ZN(n2771) );
  AOI22_X1 \ashr_130/*cell*849423  ( .A1(n2839), .A2(n2743), .B1(n2742), .B2(
        n1916), .ZN(n2764) );
  AOI22_X1 \ashr_130/*cell*849424  ( .A1(n2842), .A2(n2762), .B1(n2765), .B2(
        n1930), .ZN(n2779) );
  AOI22_X1 \ashr_130/*cell*849425  ( .A1(n2839), .A2(n2741), .B1(n2740), .B2(
        n1916), .ZN(n2765) );
  AOI22_X1 \ashr_130/*cell*849426  ( .A1(n2839), .A2(n2739), .B1(n2738), .B2(
        n1916), .ZN(n2762) );
  OAI21_X1 \ashr_130/*cell*849427  ( .B1(n2847), .B2(n2791), .A(n2737), .ZN(
        \DataP/ALU_C/shifter/N62 ) );
  NAND2_X1 \ashr_130/*cell*849428  ( .A1(n2065), .A2(n2736), .ZN(n2737) );
  AOI22_X1 \ashr_130/*cell*849429  ( .A1(n1915), .A2(n2777), .B1(n2812), .B2(
        n2845), .ZN(n2736) );
  AOI22_X1 \ashr_130/*cell*849430  ( .A1(n2842), .A2(n2735), .B1(n2734), .B2(
        n1930), .ZN(n2812) );
  AOI22_X1 \ashr_130/*cell*849431  ( .A1(n2842), .A2(n2733), .B1(n2732), .B2(
        n1930), .ZN(n2777) );
  NAND3_X1 \ashr_130/*cell*849432  ( .A1(n2064), .A2(n1930), .A3(n2776), .ZN(
        n2791) );
  MUX2_X1 \ashr_130/*cell*849434  ( .A(n2731), .B(n2790), .S(\lt_x_135/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N61 ) );
  NOR2_X1 \ashr_130/*cell*849435  ( .A1(n1915), .A2(n2769), .ZN(n2790) );
  AOI22_X1 \ashr_130/*cell*849436  ( .A1(n2842), .A2(n2784), .B1(n2756), .B2(
        n2844), .ZN(n2769) );
  AOI22_X1 \ashr_130/*cell*849437  ( .A1(n2839), .A2(n2746), .B1(n2739), .B2(
        n1916), .ZN(n2756) );
  AOI22_X1 \ashr_130/*cell*849438  ( .A1(n1914), .A2(\DataP/alu_a_in[28] ), 
        .B1(\DataP/alu_a_in[27] ), .B2(n1931), .ZN(n2739) );
  AOI22_X1 \ashr_130/*cell*849439  ( .A1(n1914), .A2(\DataP/alu_a_in[30] ), 
        .B1(\DataP/alu_a_in[29] ), .B2(n1931), .ZN(n2746) );
  NOR2_X1 \ashr_130/*cell*849440  ( .A1(n2840), .A2(n2747), .ZN(n2784) );
  NAND2_X1 \ashr_130/*cell*849441  ( .A1(\DataP/alu_a_in[31] ), .A2(n1931), 
        .ZN(n2747) );
  AOI22_X1 \ashr_130/*cell*849442  ( .A1(n1915), .A2(n2768), .B1(n2807), .B2(
        n2845), .ZN(n2731) );
  AOI22_X1 \ashr_130/*cell*849443  ( .A1(n2842), .A2(n2757), .B1(n2826), .B2(
        n1930), .ZN(n2807) );
  AOI22_X1 \ashr_130/*cell*849444  ( .A1(n2839), .A2(n2744), .B1(n2770), .B2(
        n1916), .ZN(n2826) );
  AOI22_X1 \ashr_130/*cell*849445  ( .A1(n1914), .A2(\DataP/alu_a_in[12] ), 
        .B1(\DataP/alu_a_in[11] ), .B2(n1931), .ZN(n2770) );
  AOI22_X1 \ashr_130/*cell*849446  ( .A1(n1914), .A2(\DataP/alu_a_in[14] ), 
        .B1(\DataP/alu_a_in[13] ), .B2(n1931), .ZN(n2744) );
  AOI22_X1 \ashr_130/*cell*849447  ( .A1(n2839), .A2(n2742), .B1(n2745), .B2(
        n1916), .ZN(n2757) );
  AOI22_X1 \ashr_130/*cell*849448  ( .A1(n1914), .A2(\DataP/alu_a_in[16] ), 
        .B1(n1841), .B2(n1931), .ZN(n2745) );
  AOI22_X1 \ashr_130/*cell*849449  ( .A1(n1914), .A2(\DataP/alu_a_in[18] ), 
        .B1(\DataP/alu_a_in[17] ), .B2(n1931), .ZN(n2742) );
  AOI22_X1 \ashr_130/*cell*849450  ( .A1(n2842), .A2(n2755), .B1(n2758), .B2(
        n2844), .ZN(n2768) );
  AOI22_X1 \ashr_130/*cell*849451  ( .A1(n2839), .A2(n2740), .B1(n2743), .B2(
        n1916), .ZN(n2758) );
  AOI22_X1 \ashr_130/*cell*849452  ( .A1(n1914), .A2(\DataP/alu_a_in[20] ), 
        .B1(n1553), .B2(n1931), .ZN(n2743) );
  AOI22_X1 \ashr_130/*cell*849453  ( .A1(n1914), .A2(\DataP/alu_a_in[22] ), 
        .B1(\DataP/alu_a_in[21] ), .B2(n1931), .ZN(n2740) );
  AOI22_X1 \ashr_130/*cell*849454  ( .A1(n2839), .A2(n2738), .B1(n2741), .B2(
        n1916), .ZN(n2755) );
  AOI22_X1 \ashr_130/*cell*849455  ( .A1(n1914), .A2(\DataP/alu_a_in[24] ), 
        .B1(\DataP/alu_a_in[23] ), .B2(n1931), .ZN(n2741) );
  AOI22_X1 \ashr_130/*cell*849456  ( .A1(n1914), .A2(\DataP/alu_a_in[26] ), 
        .B1(\DataP/alu_a_in[25] ), .B2(n1931), .ZN(n2738) );
  MUX2_X1 \ashr_130/*cell*849457  ( .A(n2730), .B(n2789), .S(\lt_x_135/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N60 ) );
  NOR2_X1 \ashr_130/*cell*849458  ( .A1(n1915), .A2(n2767), .ZN(n2789) );
  AOI22_X1 \ashr_130/*cell*849459  ( .A1(n2842), .A2(n2781), .B1(n2750), .B2(
        n2844), .ZN(n2767) );
  AOI22_X1 \ashr_130/*cell*849460  ( .A1(n2839), .A2(n2729), .B1(n2728), .B2(
        n1916), .ZN(n2750) );
  NOR2_X1 \ashr_130/*cell*849461  ( .A1(n2840), .A2(n2727), .ZN(n2781) );
  AOI22_X1 \ashr_130/*cell*849462  ( .A1(n1915), .A2(n2766), .B1(n2799), .B2(
        n2845), .ZN(n2730) );
  AOI22_X1 \ashr_130/*cell*849463  ( .A1(n2842), .A2(n2751), .B1(n2821), .B2(
        n2844), .ZN(n2799) );
  AOI22_X1 \ashr_130/*cell*849464  ( .A1(n2840), .A2(n2726), .B1(n2725), .B2(
        n1916), .ZN(n2821) );
  AOI22_X1 \ashr_130/*cell*849465  ( .A1(n2839), .A2(n2724), .B1(n2723), .B2(
        n1916), .ZN(n2751) );
  AOI22_X1 \ashr_130/*cell*849466  ( .A1(n2843), .A2(n2749), .B1(n2752), .B2(
        n2844), .ZN(n2766) );
  AOI22_X1 \ashr_130/*cell*849467  ( .A1(n2840), .A2(n2722), .B1(n2721), .B2(
        n1916), .ZN(n2752) );
  AOI22_X1 \ashr_130/*cell*849468  ( .A1(n2840), .A2(n2720), .B1(n2719), .B2(
        n1916), .ZN(n2749) );
  MUX2_X1 \ashr_130/*cell*849469  ( .A(n2718), .B(n2761), .S(\lt_x_135/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N50 ) );
  AOI22_X1 \ashr_130/*cell*849470  ( .A1(n1915), .A2(n2787), .B1(n2831), .B2(
        n2845), .ZN(n2761) );
  AOI22_X1 \ashr_130/*cell*849471  ( .A1(n2843), .A2(n2732), .B1(n2735), .B2(
        n2844), .ZN(n2831) );
  AOI22_X1 \ashr_130/*cell*849472  ( .A1(n2840), .A2(n2721), .B1(n2724), .B2(
        n1916), .ZN(n2735) );
  AOI22_X1 \ashr_130/*cell*849473  ( .A1(n1914), .A2(\DataP/alu_a_in[17] ), 
        .B1(\DataP/alu_a_in[16] ), .B2(n1931), .ZN(n2724) );
  AOI22_X1 \ashr_130/*cell*849474  ( .A1(n1914), .A2(\DataP/alu_a_in[19] ), 
        .B1(\DataP/alu_a_in[18] ), .B2(n1931), .ZN(n2721) );
  AOI22_X1 \ashr_130/*cell*849475  ( .A1(n2840), .A2(n2719), .B1(n2722), .B2(
        n1916), .ZN(n2732) );
  AOI22_X1 \ashr_130/*cell*849476  ( .A1(n1914), .A2(\DataP/alu_a_in[21] ), 
        .B1(\DataP/alu_a_in[20] ), .B2(n1931), .ZN(n2722) );
  AOI22_X1 \ashr_130/*cell*849477  ( .A1(n1914), .A2(\DataP/alu_a_in[23] ), 
        .B1(\DataP/alu_a_in[22] ), .B2(n1931), .ZN(n2719) );
  AOI22_X1 \ashr_130/*cell*849478  ( .A1(n2843), .A2(n2776), .B1(n2733), .B2(
        n2844), .ZN(n2787) );
  AOI22_X1 \ashr_130/*cell*849479  ( .A1(n2840), .A2(n2728), .B1(n2720), .B2(
        n1916), .ZN(n2733) );
  AOI22_X1 \ashr_130/*cell*849480  ( .A1(n1914), .A2(\DataP/alu_a_in[25] ), 
        .B1(\DataP/alu_a_in[24] ), .B2(n1931), .ZN(n2720) );
  AOI22_X1 \ashr_130/*cell*849481  ( .A1(n1914), .A2(\DataP/alu_a_in[27] ), 
        .B1(\DataP/alu_a_in[26] ), .B2(n1931), .ZN(n2728) );
  AOI22_X1 \ashr_130/*cell*849482  ( .A1(n2840), .A2(n2727), .B1(n2729), .B2(
        n1916), .ZN(n2776) );
  AOI22_X1 \ashr_130/*cell*849483  ( .A1(n1914), .A2(\DataP/alu_a_in[29] ), 
        .B1(\DataP/alu_a_in[28] ), .B2(n1931), .ZN(n2729) );
  AOI22_X1 \ashr_130/*cell*849484  ( .A1(n1914), .A2(\DataP/alu_a_in[31] ), 
        .B1(\DataP/alu_a_in[30] ), .B2(n1931), .ZN(n2727) );
  AOI22_X1 \ashr_130/*cell*849485  ( .A1(n2846), .A2(n2830), .B1(n2717), .B2(
        n2064), .ZN(n2718) );
  AOI21_X1 \ashr_130/*cell*849487  ( .B1(n2841), .B2(n2809), .A(n2716), .ZN(
        n2717) );
  AOI221_X1 \ashr_130/*cell*849488  ( .B1(n2795), .B2(n2839), .C1(n2715), .C2(
        n1916), .A(n2841), .ZN(n2716) );
  AOI22_X1 \ashr_130/*cell*849489  ( .A1(n1914), .A2(\DataP/alu_a_in[1] ), 
        .B1(n1605), .B2(n1931), .ZN(n2715) );
  AOI22_X1 \ashr_130/*cell*849490  ( .A1(n1914), .A2(\DataP/alu_a_in[3] ), 
        .B1(\DataP/alu_a_in[2] ), .B2(n1931), .ZN(n2795) );
  AOI22_X1 \ashr_130/*cell*849491  ( .A1(n2840), .A2(n2793), .B1(n2796), .B2(
        n1916), .ZN(n2809) );
  AOI22_X1 \ashr_130/*cell*849492  ( .A1(n1914), .A2(\DataP/alu_a_in[5] ), 
        .B1(\DataP/alu_a_in[4] ), .B2(n1931), .ZN(n2796) );
  AOI22_X1 \ashr_130/*cell*849493  ( .A1(n1914), .A2(\DataP/alu_a_in[7] ), 
        .B1(\DataP/alu_a_in[6] ), .B2(n1931), .ZN(n2793) );
  AOI22_X1 \ashr_130/*cell*849494  ( .A1(n2842), .A2(n2734), .B1(n2810), .B2(
        n1930), .ZN(n2830) );
  AOI22_X1 \ashr_130/*cell*849496  ( .A1(n2840), .A2(n2725), .B1(n2794), .B2(
        n1916), .ZN(n2810) );
  AOI22_X1 \ashr_130/*cell*849497  ( .A1(n1914), .A2(\DataP/alu_a_in[9] ), 
        .B1(\DataP/alu_a_in[8] ), .B2(n1931), .ZN(n2794) );
  AOI22_X1 \ashr_130/*cell*849498  ( .A1(n1914), .A2(\DataP/alu_a_in[11] ), 
        .B1(\DataP/alu_a_in[10] ), .B2(n1931), .ZN(n2725) );
  AOI22_X1 \ashr_130/*cell*849499  ( .A1(n2839), .A2(n2723), .B1(n2726), .B2(
        n1916), .ZN(n2734) );
  AOI22_X1 \ashr_130/*cell*849501  ( .A1(n1914), .A2(\DataP/alu_a_in[13] ), 
        .B1(\DataP/alu_a_in[12] ), .B2(n1931), .ZN(n2726) );
  AOI22_X1 \ashr_130/*cell*849502  ( .A1(n1914), .A2(\DataP/alu_a_in[15] ), 
        .B1(\DataP/alu_a_in[14] ), .B2(n1931), .ZN(n2723) );
  MUX2_X1 \ash_129/*cell*849520  ( .A(n2689), .B(n2688), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N49 ) );
  AOI22_X1 \ash_129/*cell*849521  ( .A1(n2846), .A2(n2687), .B1(n2686), .B2(
        n2064), .ZN(n2689) );
  AOI22_X1 \ash_129/*cell*849522  ( .A1(n2714), .A2(n2685), .B1(n2684), .B2(
        n1930), .ZN(n2686) );
  AOI22_X1 \ash_129/*cell*849523  ( .A1(n2713), .A2(n2683), .B1(n2682), .B2(
        n1916), .ZN(n2684) );
  AOI22_X1 \ash_129/*cell*849524  ( .A1(n2709), .A2(\DataP/alu_a_in[30] ), 
        .B1(\DataP/alu_a_in[31] ), .B2(n2711), .ZN(n2682) );
  MUX2_X1 \ash_129/*cell*849525  ( .A(n2681), .B(n2680), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N48 ) );
  AOI22_X1 \ash_129/*cell*849526  ( .A1(n1915), .A2(n2679), .B1(n2678), .B2(
        n2845), .ZN(n2681) );
  AOI22_X1 \ash_129/*cell*849527  ( .A1(n2714), .A2(n2677), .B1(n2676), .B2(
        n2989), .ZN(n2678) );
  AOI22_X1 \ash_129/*cell*849528  ( .A1(n2713), .A2(n2675), .B1(n2674), .B2(
        n1916), .ZN(n2676) );
  AOI22_X1 \ash_129/*cell*849529  ( .A1(n2709), .A2(\DataP/alu_a_in[29] ), 
        .B1(\DataP/alu_a_in[30] ), .B2(n2710), .ZN(n2674) );
  MUX2_X1 \ash_129/*cell*849532  ( .A(n2672), .B(n2671), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N47 ) );
  AOI22_X1 \ash_129/*cell*849533  ( .A1(n1915), .A2(n2670), .B1(n2669), .B2(
        n2064), .ZN(n2672) );
  AOI22_X1 \ash_129/*cell*849534  ( .A1(n2714), .A2(n2668), .B1(n2667), .B2(
        n1913), .ZN(n2669) );
  AOI22_X1 \ash_129/*cell*849535  ( .A1(n2713), .A2(n2666), .B1(n2683), .B2(
        n1916), .ZN(n2667) );
  AOI22_X1 \ash_129/*cell*849536  ( .A1(n2709), .A2(\DataP/alu_a_in[28] ), 
        .B1(\DataP/alu_a_in[29] ), .B2(n2711), .ZN(n2683) );
  MUX2_X1 \ash_129/*cell*849537  ( .A(n2665), .B(n2664), .S(\lt_x_135/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N46 ) );
  AOI22_X1 \ash_129/*cell*849538  ( .A1(n1915), .A2(n2663), .B1(n2662), .B2(
        n2064), .ZN(n2665) );
  AOI22_X1 \ash_129/*cell*849539  ( .A1(n2714), .A2(n2661), .B1(n2660), .B2(
        n1930), .ZN(n2662) );
  AOI22_X1 \ash_129/*cell*849540  ( .A1(n2713), .A2(n2659), .B1(n2675), .B2(
        n1916), .ZN(n2660) );
  AOI22_X1 \ash_129/*cell*849541  ( .A1(n2709), .A2(\DataP/alu_a_in[27] ), 
        .B1(\DataP/alu_a_in[28] ), .B2(n2711), .ZN(n2675) );
  AOI22_X1 \ash_129/*cell*849545  ( .A1(n2713), .A2(n2655), .B1(n2666), .B2(
        n1916), .ZN(n2685) );
  AOI22_X1 \ash_129/*cell*849546  ( .A1(n2709), .A2(\DataP/alu_a_in[26] ), 
        .B1(\DataP/alu_a_in[27] ), .B2(n2711), .ZN(n2666) );
  AOI22_X1 \ash_129/*cell*849550  ( .A1(n2713), .A2(n2651), .B1(n2659), .B2(
        n1916), .ZN(n2677) );
  AOI22_X1 \ash_129/*cell*849551  ( .A1(n2709), .A2(\DataP/alu_a_in[25] ), 
        .B1(\DataP/alu_a_in[26] ), .B2(n2711), .ZN(n2659) );
  MUX2_X1 \ash_129/*cell*849552  ( .A(n2650), .B(n2696), .S(\lt_x_135/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N43 ) );
  AOI22_X1 \ash_129/*cell*849553  ( .A1(n1915), .A2(n2649), .B1(n2648), .B2(
        n2845), .ZN(n2696) );
  AOI22_X1 \ash_129/*cell*849554  ( .A1(n1915), .A2(n2647), .B1(n2646), .B2(
        n2845), .ZN(n2650) );
  AOI22_X1 \ash_129/*cell*849555  ( .A1(n2842), .A2(n2645), .B1(n2668), .B2(
        n1913), .ZN(n2646) );
  AOI22_X1 \ash_129/*cell*849556  ( .A1(n2713), .A2(n2644), .B1(n2655), .B2(
        n1916), .ZN(n2668) );
  AOI22_X1 \ash_129/*cell*849557  ( .A1(n2709), .A2(\DataP/alu_a_in[24] ), 
        .B1(\DataP/alu_a_in[25] ), .B2(n2710), .ZN(n2655) );
  MUX2_X1 \ash_129/*cell*849558  ( .A(n2643), .B(n2695), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N42 ) );
  AOI22_X1 \ash_129/*cell*849559  ( .A1(n1915), .A2(n2642), .B1(n2641), .B2(
        n2127), .ZN(n2695) );
  AOI22_X1 \ash_129/*cell*849560  ( .A1(n1915), .A2(n2640), .B1(n2639), .B2(
        n2845), .ZN(n2643) );
  AOI22_X1 \ash_129/*cell*849561  ( .A1(n2842), .A2(n2638), .B1(n2661), .B2(
        n1913), .ZN(n2639) );
  AOI22_X1 \ash_129/*cell*849562  ( .A1(n2713), .A2(n2637), .B1(n2651), .B2(
        n1916), .ZN(n2661) );
  AOI22_X1 \ash_129/*cell*849563  ( .A1(n2709), .A2(\DataP/alu_a_in[23] ), 
        .B1(\DataP/alu_a_in[24] ), .B2(n2710), .ZN(n2651) );
  NOR2_X1 \ash_129/*cell*849565  ( .A1(n1915), .A2(n2636), .ZN(n2694) );
  AOI22_X1 \ash_129/*cell*849567  ( .A1(n2842), .A2(n2634), .B1(n2656), .B2(
        n1913), .ZN(n2687) );
  AOI22_X1 \ash_129/*cell*849568  ( .A1(n2713), .A2(n2633), .B1(n2644), .B2(
        n1916), .ZN(n2656) );
  AOI22_X1 \ash_129/*cell*849569  ( .A1(n2709), .A2(\DataP/alu_a_in[22] ), 
        .B1(\DataP/alu_a_in[23] ), .B2(n2711), .ZN(n2644) );
  MUX2_X1 \ash_129/*cell*849570  ( .A(n2632), .B(n2693), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N40 ) );
  NOR2_X1 \ash_129/*cell*849571  ( .A1(n1915), .A2(n2631), .ZN(n2693) );
  AOI22_X1 \ash_129/*cell*849572  ( .A1(n1915), .A2(n2630), .B1(n2679), .B2(
        n2127), .ZN(n2632) );
  AOI22_X1 \ash_129/*cell*849573  ( .A1(n2842), .A2(n2629), .B1(n2652), .B2(
        n1913), .ZN(n2679) );
  AOI22_X1 \ash_129/*cell*849574  ( .A1(n2839), .A2(n2628), .B1(n2637), .B2(
        n1916), .ZN(n2652) );
  AOI22_X1 \ash_129/*cell*849575  ( .A1(n2709), .A2(\DataP/alu_a_in[21] ), 
        .B1(\DataP/alu_a_in[22] ), .B2(n2710), .ZN(n2637) );
  NOR2_X1 \ash_129/*cell*849577  ( .A1(n1915), .A2(n2627), .ZN(n2692) );
  AOI22_X1 \ash_129/*cell*849579  ( .A1(n2842), .A2(n2625), .B1(n2645), .B2(
        n1913), .ZN(n2670) );
  AOI22_X1 \ash_129/*cell*849580  ( .A1(\sra_131/SH[1] ), .A2(n2624), .B1(
        n2633), .B2(n1916), .ZN(n2645) );
  AOI22_X1 \ash_129/*cell*849581  ( .A1(n2709), .A2(\DataP/alu_a_in[20] ), 
        .B1(\DataP/alu_a_in[21] ), .B2(n2710), .ZN(n2633) );
  MUX2_X1 \ash_129/*cell*849582  ( .A(n2623), .B(n2691), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N38 ) );
  NOR2_X1 \ash_129/*cell*849583  ( .A1(n1915), .A2(n2622), .ZN(n2691) );
  AOI22_X1 \ash_129/*cell*849584  ( .A1(n1915), .A2(n2621), .B1(n2663), .B2(
        n2330), .ZN(n2623) );
  AOI22_X1 \ash_129/*cell*849585  ( .A1(n2842), .A2(n2620), .B1(n2638), .B2(
        n1913), .ZN(n2663) );
  AOI22_X1 \ash_129/*cell*849586  ( .A1(n2839), .A2(n2619), .B1(n2628), .B2(
        n1916), .ZN(n2638) );
  AOI22_X1 \ash_129/*cell*849587  ( .A1(n2709), .A2(\DataP/alu_a_in[19] ), 
        .B1(\DataP/alu_a_in[20] ), .B2(n2710), .ZN(n2628) );
  NOR2_X1 \ash_129/*cell*849588  ( .A1(\lt_x_135/B[4] ), .A2(n2703), .ZN(
        \DataP/ALU_C/shifter/N19 ) );
  MUX2_X1 \ash_129/*cell*849590  ( .A(n2617), .B(n2690), .S(\lt_x_134/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N37 ) );
  NOR2_X1 \ash_129/*cell*849591  ( .A1(n1915), .A2(n2616), .ZN(n2690) );
  AOI22_X1 \ash_129/*cell*849592  ( .A1(n1915), .A2(n2615), .B1(n2657), .B2(
        n2845), .ZN(n2617) );
  AOI22_X1 \ash_129/*cell*849593  ( .A1(n2842), .A2(n2614), .B1(n2634), .B2(
        n1913), .ZN(n2657) );
  AOI22_X1 \ash_129/*cell*849594  ( .A1(n2840), .A2(n2613), .B1(n2624), .B2(
        n1916), .ZN(n2634) );
  AOI22_X1 \ash_129/*cell*849595  ( .A1(n2709), .A2(\DataP/alu_a_in[18] ), 
        .B1(\DataP/alu_a_in[19] ), .B2(n2710), .ZN(n2624) );
  NOR2_X1 \ash_129/*cell*849597  ( .A1(n2846), .A2(n2612), .ZN(n2673) );
  AOI22_X1 \ash_129/*cell*849599  ( .A1(n2842), .A2(n2610), .B1(n2629), .B2(
        n1913), .ZN(n2653) );
  AOI22_X1 \ash_129/*cell*849600  ( .A1(n2839), .A2(n2609), .B1(n2619), .B2(
        n1916), .ZN(n2629) );
  AOI22_X1 \ash_129/*cell*849601  ( .A1(n2709), .A2(\DataP/alu_a_in[17] ), 
        .B1(\DataP/alu_a_in[18] ), .B2(n2710), .ZN(n2619) );
  NOR2_X1 \ash_129/*cell*849603  ( .A1(n2846), .A2(n2649), .ZN(n2618) );
  NAND2_X1 \ash_129/*cell*849604  ( .A1(n2608), .A2(n1913), .ZN(n2649) );
  AOI22_X1 \ash_129/*cell*849606  ( .A1(n2842), .A2(n2607), .B1(n2625), .B2(
        n1913), .ZN(n2647) );
  AOI22_X1 \ash_129/*cell*849607  ( .A1(n2840), .A2(n2606), .B1(n2613), .B2(
        n1916), .ZN(n2625) );
  AOI22_X1 \ash_129/*cell*849608  ( .A1(n2709), .A2(\DataP/alu_a_in[16] ), 
        .B1(\DataP/alu_a_in[17] ), .B2(n2710), .ZN(n2613) );
  AOI22_X1 \ash_129/*cell*849609  ( .A1(n2842), .A2(n2605), .B1(n2604), .B2(
        n1913), .ZN(n2648) );
  MUX2_X1 \ash_129/*cell*849610  ( .A(n2603), .B(n2602), .S(\lt_x_135/B[4] ), 
        .Z(\DataP/ALU_C/shifter/N34 ) );
  AOI22_X1 \ash_129/*cell*849611  ( .A1(n1915), .A2(n2641), .B1(n2640), .B2(
        n2845), .ZN(n2603) );
  AOI22_X1 \ash_129/*cell*849612  ( .A1(n2842), .A2(n2601), .B1(n2620), .B2(
        n1913), .ZN(n2640) );
  AOI22_X1 \ash_129/*cell*849613  ( .A1(n2840), .A2(n2600), .B1(n2609), .B2(
        n1916), .ZN(n2620) );
  AOI22_X1 \ash_129/*cell*849614  ( .A1(n2709), .A2(n1841), .B1(
        \DataP/alu_a_in[16] ), .B2(n2710), .ZN(n2609) );
  AOI22_X1 \ash_129/*cell*849615  ( .A1(n2842), .A2(n2599), .B1(n2598), .B2(
        n1913), .ZN(n2641) );
  NOR2_X1 \ash_129/*cell*849616  ( .A1(\lt_x_134/B[4] ), .A2(n2702), .ZN(
        \DataP/ALU_C/shifter/N33 ) );
  AOI22_X1 \ash_129/*cell*849618  ( .A1(n2846), .A2(n2636), .B1(n2635), .B2(
        n2127), .ZN(n2688) );
  AOI22_X1 \ash_129/*cell*849619  ( .A1(n2841), .A2(n2597), .B1(n2614), .B2(
        n1913), .ZN(n2635) );
  AOI22_X1 \ash_129/*cell*849620  ( .A1(n2839), .A2(n2596), .B1(n2606), .B2(
        n1916), .ZN(n2614) );
  AOI22_X1 \ash_129/*cell*849621  ( .A1(n2709), .A2(\DataP/alu_a_in[14] ), 
        .B1(\DataP/alu_a_in[15] ), .B2(n2710), .ZN(n2606) );
  AOI22_X1 \ash_129/*cell*849622  ( .A1(n2841), .A2(n2595), .B1(n2594), .B2(
        n1913), .ZN(n2636) );
  NOR2_X1 \ash_129/*cell*849623  ( .A1(\lt_x_135/B[4] ), .A2(n2701), .ZN(
        \DataP/ALU_C/shifter/N32 ) );
  AOI22_X1 \ash_129/*cell*849625  ( .A1(n1915), .A2(n2631), .B1(n2630), .B2(
        n2845), .ZN(n2680) );
  AOI22_X1 \ash_129/*cell*849626  ( .A1(n2841), .A2(n2593), .B1(n2610), .B2(
        n2989), .ZN(n2630) );
  AOI22_X1 \ash_129/*cell*849627  ( .A1(n2839), .A2(n2592), .B1(n2600), .B2(
        n1916), .ZN(n2610) );
  AOI22_X1 \ash_129/*cell*849628  ( .A1(n2709), .A2(\DataP/alu_a_in[13] ), 
        .B1(\DataP/alu_a_in[14] ), .B2(n2710), .ZN(n2600) );
  AOI22_X1 \ash_129/*cell*849629  ( .A1(n2841), .A2(n2591), .B1(n2590), .B2(
        n1913), .ZN(n2631) );
  NOR2_X1 \ash_129/*cell*849630  ( .A1(\lt_x_134/B[4] ), .A2(n2700), .ZN(
        \DataP/ALU_C/shifter/N31 ) );
  AOI22_X1 \ash_129/*cell*849632  ( .A1(n2846), .A2(n2627), .B1(n2626), .B2(
        n2127), .ZN(n2671) );
  AOI22_X1 \ash_129/*cell*849633  ( .A1(n2841), .A2(n2604), .B1(n2607), .B2(
        n1913), .ZN(n2626) );
  AOI22_X1 \ash_129/*cell*849634  ( .A1(n2839), .A2(n2589), .B1(n2596), .B2(
        n1916), .ZN(n2607) );
  AOI22_X1 \ash_129/*cell*849635  ( .A1(n2709), .A2(\DataP/alu_a_in[12] ), 
        .B1(\DataP/alu_a_in[13] ), .B2(n2710), .ZN(n2596) );
  AOI22_X1 \ash_129/*cell*849636  ( .A1(n2839), .A2(n2588), .B1(n2587), .B2(
        n1916), .ZN(n2604) );
  AOI22_X1 \ash_129/*cell*849637  ( .A1(n2841), .A2(n2608), .B1(n2605), .B2(
        n1913), .ZN(n2627) );
  AOI22_X1 \ash_129/*cell*849638  ( .A1(n2713), .A2(n2586), .B1(n2585), .B2(
        n1916), .ZN(n2605) );
  NOR2_X1 \ash_129/*cell*849639  ( .A1(n2713), .A2(n2584), .ZN(n2608) );
  NOR2_X1 \ash_129/*cell*849640  ( .A1(\lt_x_135/B[4] ), .A2(n2699), .ZN(
        \DataP/ALU_C/shifter/N30 ) );
  AOI22_X1 \ash_129/*cell*849642  ( .A1(n2846), .A2(n2622), .B1(n2621), .B2(
        n2064), .ZN(n2664) );
  AOI22_X1 \ash_129/*cell*849643  ( .A1(n2841), .A2(n2598), .B1(n2601), .B2(
        n1913), .ZN(n2621) );
  AOI22_X1 \ash_129/*cell*849644  ( .A1(n2713), .A2(n2583), .B1(n2592), .B2(
        n1916), .ZN(n2601) );
  AOI22_X1 \ash_129/*cell*849645  ( .A1(n2709), .A2(\DataP/alu_a_in[11] ), 
        .B1(\DataP/alu_a_in[12] ), .B2(n2710), .ZN(n2592) );
  AOI22_X1 \ash_129/*cell*849646  ( .A1(n2713), .A2(n2582), .B1(n2581), .B2(
        n1916), .ZN(n2598) );
  AOI22_X1 \ash_129/*cell*849648  ( .A1(n2713), .A2(n2580), .B1(n2579), .B2(
        n1916), .ZN(n2599) );
  NOR2_X1 \ash_129/*cell*849650  ( .A1(\lt_x_135/B[4] ), .A2(n2698), .ZN(
        \DataP/ALU_C/shifter/N29 ) );
  AOI22_X1 \ash_129/*cell*849652  ( .A1(n2846), .A2(n2616), .B1(n2615), .B2(
        n2127), .ZN(n2658) );
  AOI22_X1 \ash_129/*cell*849653  ( .A1(n2842), .A2(n2594), .B1(n2597), .B2(
        n1913), .ZN(n2615) );
  AOI22_X1 \ash_129/*cell*849654  ( .A1(n2713), .A2(n2587), .B1(n2589), .B2(
        n1916), .ZN(n2597) );
  AOI22_X1 \ash_129/*cell*849655  ( .A1(n2709), .A2(\DataP/alu_a_in[10] ), 
        .B1(\DataP/alu_a_in[11] ), .B2(n2710), .ZN(n2589) );
  AOI22_X1 \ash_129/*cell*849656  ( .A1(n2709), .A2(\DataP/alu_a_in[8] ), .B1(
        \DataP/alu_a_in[9] ), .B2(n2711), .ZN(n2587) );
  AOI22_X1 \ash_129/*cell*849657  ( .A1(n2713), .A2(n2585), .B1(n2588), .B2(
        n1916), .ZN(n2594) );
  AOI22_X1 \ash_129/*cell*849658  ( .A1(n2709), .A2(\DataP/alu_a_in[6] ), .B1(
        \DataP/alu_a_in[7] ), .B2(n2711), .ZN(n2588) );
  AOI22_X1 \ash_129/*cell*849659  ( .A1(n2709), .A2(\DataP/alu_a_in[4] ), .B1(
        \DataP/alu_a_in[5] ), .B2(n2711), .ZN(n2585) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[5]  ( .D(n2161), .CK(Clk), .SN(Rst), 
        .Q(n3049), .QN(\DataP/opcode_W[5] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[1]  ( .D(n2559), .CK(Clk), .SN(Rst), .QN(
        \DataP/Rs2[1] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[0]  ( .D(n2558), .CK(Clk), .SN(Rst), .Q(
        n1885), .QN(\DataP/Rs2[0] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[3]  ( .D(n2557), .CK(Clk), .SN(Rst), .QN(
        \DataP/Rs2[3] ) );
  DFFS_X1 \DataP/MEM_WB_s/RD_OUT_reg[1]  ( .D(n529), .CK(Clk), .SN(Rst), .Q(
        n1891), .QN(\DataP/add_D[1] ) );
  DFFS_X1 \DataP/MEM_WB_s/RD_OUT_reg[3]  ( .D(n2570), .CK(Clk), .SN(Rst), .Q(
        n2568), .QN(\DataP/add_D[3] ) );
  DFFS_X2 \DataP/IF_IDs/IR_OUT_reg[28]  ( .D(IRAM_DATA_OUT[28]), .CK(Clk), 
        .SN(n164), .Q(IR_CU_28), .QN(n510) );
  DFFS_X1 \DataP/IF_IDs/IR_OUT_reg[30]  ( .D(IRAM_DATA_OUT[30]), .CK(Clk), 
        .SN(n164), .Q(n2129), .QN(n515) );
  DFF_X2 \DataP/PC_reg/O_reg[29]  ( .D(\DataP/PC_reg/N31 ), .CK(Clk), .Q(
        \DataP/pc_out[29] ) );
  AOI21_X1 \lt_x_134/*cell*849092  ( .B1(\DataP/alu_a_in[4] ), .B2(n2847), .A(
        n2023), .ZN(n2024) );
  NOR2_X1 \lt_x_134/*cell*849116  ( .A1(n1572), .A2(n1863), .ZN(n2028) );
  NAND2_X1 \lt_x_134/*cell*849143  ( .A1(\DataP/alu_b_in[31] ), .A2(n1923), 
        .ZN(n2013) );
  DFF_X2 \DataP/PC_reg/O_reg[30]  ( .D(\DataP/PC_reg/N32 ), .CK(Clk), .Q(
        \DataP/pc_out[30] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[26]  ( .D(n1599), .CK(Clk), .SN(Rst), 
        .Q(n2169), .QN(\DataP/alu_out_M[26] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[31]  ( .D(n297), .CK(Clk), .SN(Rst), .Q(
        n2185), .QN(\DataP/alu_out_M[31] ) );
  DFFR_X1 \DataP/EX_MEM_s/RD_OUT_reg[0]  ( .D(n1956), .CK(Clk), .RN(Rst), .Q(
        \DataP/dest_M[0] ), .QN(n528) );
  DFFR_X1 \DataP/MEM_WB_s/RD_OUT_reg[2]  ( .D(\DataP/dest_M[2] ), .CK(Clk), 
        .RN(Rst), .Q(\DataP/add_D[2] ), .QN(n538) );
  DFF_X1 \DataP/PC_reg/O_reg[31]  ( .D(\DataP/PC_reg/N33 ), .CK(Clk), .Q(
        \DataP/pc_out[31] ) );
  DFFR_X1 \CU_I/cw1_reg[4]  ( .D(\CU_I/cw[4] ), .CK(Clk), .RN(Rst), .QN(n132)
         );
  DFFR_X1 \CU_I/cw1_reg[6]  ( .D(\CU_I/cw[6] ), .CK(Clk), .RN(Rst), .QN(n130)
         );
  DFFR_X1 \CU_I/cw1_reg[3]  ( .D(\CU_I/cw[3] ), .CK(Clk), .RN(Rst), .QN(n131)
         );
  DFFR_X1 \CU_I/cw1_reg[7]  ( .D(\CU_I/cw[7] ), .CK(Clk), .RN(Rst), .QN(n143)
         );
  DFFR_X1 \CU_I/cw1_reg[1]  ( .D(\CU_I/cw[1] ), .CK(Clk), .RN(Rst), .QN(n129)
         );
  DFFR_X1 \CU_I/cw1_reg[0]  ( .D(\CU_I/cw[0] ), .CK(Clk), .RN(Rst), .QN(n136)
         );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[4]  ( .D(\DataP/dest_D[4] ), .CK(Clk), .RN(
        Rst), .QN(n142) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[3]  ( .D(\DataP/dest_D[3] ), .CK(Clk), .RN(
        Rst), .QN(n141) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[2]  ( .D(\DataP/dest_D[2] ), .CK(Clk), .RN(
        Rst), .QN(n140) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[1]  ( .D(\DataP/dest_D[1] ), .CK(Clk), .RN(
        Rst), .QN(n139) );
  DFFR_X1 \DataP/ID_EXs/RD_OUT_reg[0]  ( .D(\DataP/dest_D[0] ), .CK(Clk), .RN(
        Rst), .Q(n1956) );
  DFFR_X1 \DataP/IF_IDs/PR_OUT_reg  ( .D(\DataP/prediction ), .CK(
        \DataP/IF_IDs/net834167 ), .RN(Rst), .QN(n258) );
  DFFR_X1 \DataP/ID_EXs/RS1_OUT_reg[3]  ( .D(\DataP/IR1[24] ), .CK(Clk), .RN(
        Rst), .QN(n523) );
  DFFRS_X1 \DataP/PC_reg/O_reg[13]  ( .D(\DataP/PC_reg/N15 ), .CK(Clk), .RN(
        1'b1), .SN(1'b1), .Q(\DataP/pc_out[13] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[17]  ( .D(n1604), .CK(Clk), .SN(Rst), 
        .Q(n2170), .QN(\DataP/alu_out_M[17] ) );
  DFFS_X1 \DataP/ID_EXs/RS2_OUT_reg[4]  ( .D(n1872), .CK(Clk), .SN(Rst), .QN(
        \DataP/Rs2[4] ) );
  DFFS_X1 \DataP/ID_EXs/RS1_OUT_reg[1]  ( .D(n153), .CK(Clk), .SN(Rst), .Q(
        n2160), .QN(\DataP/Rs1[1] ) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[0]  ( .D(n497), .CK(Clk), .SN(Rst), .Q(
        n151), .QN(\DataP/opcode_E[0] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[19]  ( .D(n319), .CK(Clk), .SN(Rst), .Q(
        n2174), .QN(\DataP/alu_out_M[19] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[15]  ( .D(n330), .CK(Clk), .SN(Rst), .Q(
        n2166), .QN(\DataP/alu_out_M[15] ) );
  DFFS_X1 \DataP/EX_MEM_s/ALU_OUT_reg[30]  ( .D(n2567), .CK(Clk), .SN(Rst), 
        .Q(n2187), .QN(\DataP/alu_out_M[30] ) );
  DFFS_X1 \DataP/ID_EXs/OPCODE_OUT_reg[1]  ( .D(n504), .CK(Clk), .SN(Rst), .Q(
        n520), .QN(n2573) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[4]  ( .D(n147), .CK(Clk), .SN(Rst), 
        .Q(n146), .QN(\DataP/opcode_M[4] ) );
  DFFS_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[0]  ( .D(n151), .CK(Clk), .SN(Rst), 
        .Q(n150), .QN(\DataP/opcode_M[0] ) );
  DFFR_X1 \DataP/ID_EXs/RS1_OUT_reg[0]  ( .D(\DataP/IR1[21] ), .CK(Clk), .RN(
        Rst), .QN(n2154) );
  DFF_X2 \DataP/PC_reg/O_reg[15]  ( .D(\DataP/PC_reg/N17 ), .CK(Clk), .Q(
        \DataP/pc_out[15] ) );
  DFF_X1 \DataP/PC_reg/O_reg[19]  ( .D(\DataP/PC_reg/N21 ), .CK(Clk), .Q(
        \DataP/pc_out[19] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[23]  ( .D(n1549), .CK(Clk), .SN(Rst), 
        .Q(n2168), .QN(\DataP/alu_out_M[23] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[2]  ( .D(n1543), .CK(Clk), .SN(Rst), 
        .Q(n1545), .QN(\DataP/opcode_W[2] ) );
  DFFR_X1 \DataP/EX_MEM_s/OPCODE_OUT_reg[2]  ( .D(n2574), .CK(Clk), .RN(Rst), 
        .Q(n1895), .QN(n1894) );
  DFF_X1 \DataP/PC_reg/O_reg[28]  ( .D(\DataP/PC_reg/N30 ), .CK(Clk), .Q(
        \DataP/pc_out[28] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[28]  ( .D(n1540), .CK(Clk), .SN(Rst), 
        .Q(n2178), .QN(\DataP/alu_out_M[28] ) );
  DFF_X2 \DataP/PC_reg/O_reg[26]  ( .D(\DataP/PC_reg/N28 ), .CK(Clk), .Q(
        \DataP/pc_out[26] ) );
  DFFS_X1 \DataP/MEM_WB_s/OPCODE_OUT_reg[1]  ( .D(n2576), .CK(Clk), .SN(Rst), 
        .Q(n2571), .QN(\DataP/opcode_W[1] ) );
  DFFRS_X2 \DataP/PC_reg/O_reg[22]  ( .D(\DataP/PC_reg/N24 ), .CK(Clk), .RN(
        1'b1), .SN(1'b1), .Q(\DataP/pc_out[22] ) );
  DFFS_X2 \DataP/EX_MEM_s/ALU_OUT_reg[22]  ( .D(n1519), .CK(Clk), .SN(Rst), 
        .Q(n2180), .QN(\DataP/alu_out_M[22] ) );
  BUF_X1 U1451 ( .A(n2564), .Z(n1515) );
  AND2_X2 U1452 ( .A1(\DataP/alu_a_in[0] ), .A2(n1537), .ZN(n3361) );
  AND3_X2 U1453 ( .A1(n3329), .A2(n3046), .A3(n2189), .ZN(n3328) );
  INV_X4 U1454 ( .A(n2712), .ZN(n2710) );
  INV_X1 U1455 ( .A(n3496), .ZN(n1516) );
  BUF_X1 U1456 ( .A(n1886), .Z(n1517) );
  AND3_X2 U1457 ( .A1(n3329), .A2(n3046), .A3(n399), .ZN(n1518) );
  AND3_X1 U1458 ( .A1(n3329), .A2(n3046), .A3(n399), .ZN(n3327) );
  BUF_X1 U1459 ( .A(n311), .Z(n1519) );
  NAND2_X1 U1460 ( .A1(n3458), .A2(n2299), .ZN(n1520) );
  AND2_X1 U1461 ( .A1(n1669), .A2(n1594), .ZN(n1521) );
  AND4_X1 U1462 ( .A1(n1586), .A2(n1521), .A3(n3281), .A4(n3291), .ZN(n1522)
         );
  OR2_X1 U1463 ( .A1(n3910), .A2(n3990), .ZN(n1523) );
  INV_X2 U1464 ( .A(n3689), .ZN(n3510) );
  AND4_X1 U1465 ( .A1(n3095), .A2(n3093), .A3(n3092), .A4(n3094), .ZN(n1524)
         );
  AND2_X1 U1466 ( .A1(n3105), .A2(n3106), .ZN(n1525) );
  AND2_X1 U1467 ( .A1(n3307), .A2(n3308), .ZN(n1526) );
  OR2_X1 U1468 ( .A1(n3194), .A2(n2213), .ZN(n1527) );
  INV_X2 U1469 ( .A(n1561), .ZN(\DataP/alu_a_in[2] ) );
  AND3_X2 U1470 ( .A1(n1868), .A2(n3111), .A3(n1527), .ZN(n1561) );
  BUF_X1 U1471 ( .A(n2403), .Z(n1528) );
  BUF_X2 U1472 ( .A(n3330), .Z(n3005) );
  OAI211_X1 U1473 ( .C1(n1636), .C2(n2185), .A(n3306), .B(n1809), .ZN(
        \DataP/alu_b_in[31] ) );
  AOI211_X1 U1474 ( .C1(n2055), .C2(n1772), .A(n1773), .B(n1774), .ZN(n2119)
         );
  BUF_X1 U1475 ( .A(n2542), .Z(n1529) );
  BUF_X1 U1476 ( .A(n3330), .Z(n3004) );
  AOI21_X1 U1477 ( .B1(n3001), .B2(\DataP/B_s[14] ), .A(n1671), .ZN(n1530) );
  AND2_X1 U1478 ( .A1(n2296), .A2(\DataP/alu_a_in[18] ), .ZN(n1531) );
  INV_X1 U1479 ( .A(n1863), .ZN(\DataP/alu_a_in[11] ) );
  OR2_X4 U1480 ( .A1(n3143), .A2(n3142), .ZN(\DataP/alu_a_in[27] ) );
  INV_X2 U1481 ( .A(n1603), .ZN(\DataP/alu_b_in[6] ) );
  INV_X1 U1482 ( .A(n2571), .ZN(n1532) );
  INV_X2 U1483 ( .A(n2712), .ZN(n2711) );
  BUF_X2 U1484 ( .A(n2004), .Z(n2712) );
  AND2_X1 U1485 ( .A1(n3578), .A2(n3580), .ZN(n1533) );
  NAND3_X1 U1486 ( .A1(n3310), .A2(n3309), .A3(n1526), .ZN(
        \DataP/alu_b_in[13] ) );
  AND2_X1 U1487 ( .A1(n1615), .A2(n149), .ZN(n1616) );
  XOR2_X1 U1488 ( .A(\DataP/Rs2[4] ), .B(n2569), .Z(n1534) );
  AND2_X1 U1489 ( .A1(n147), .A2(n145), .ZN(n1618) );
  AND2_X2 U1490 ( .A1(n151), .A2(n521), .ZN(n1619) );
  NAND4_X1 U1491 ( .A1(n1616), .A2(n1534), .A3(n1618), .A4(n1619), .ZN(n1535)
         );
  NOR2_X1 U1492 ( .A1(n2157), .A2(n1535), .ZN(n1617) );
  INV_X1 U1493 ( .A(n1619), .ZN(n3031) );
  NAND2_X1 U1494 ( .A1(n3381), .A2(n3377), .ZN(n1536) );
  AOI21_X1 U1495 ( .B1(n3205), .B2(n3676), .A(n1536), .ZN(n1886) );
  OAI211_X1 U1496 ( .C1(n1886), .C2(n3212), .A(n3211), .B(n3387), .ZN(n3269)
         );
  NAND4_X1 U1497 ( .A1(n1542), .A2(n3089), .A3(n3091), .A4(n3088), .ZN(n1537)
         );
  NAND2_X1 U1498 ( .A1(n1538), .A2(n1553), .ZN(n1552) );
  OR2_X1 U1499 ( .A1(n1538), .A2(\DataP/alu_a_in[19] ), .ZN(n2378) );
  NAND2_X1 U1500 ( .A1(n1699), .A2(n1700), .ZN(n1538) );
  NAND4_X1 U1501 ( .A1(n2332), .A2(n1584), .A3(n2336), .A4(n1585), .ZN(
        \DataP/alu_b_in[8] ) );
  BUF_X2 U1502 ( .A(n2560), .Z(n1539) );
  BUF_X1 U1503 ( .A(n2560), .Z(n2562) );
  BUF_X1 U1504 ( .A(n300), .Z(n1540) );
  BUF_X1 U1505 ( .A(n3455), .Z(n1541) );
  BUF_X1 U1506 ( .A(n3090), .Z(n1542) );
  BUF_X1 U1507 ( .A(n1894), .Z(n1543) );
  BUF_X1 U1508 ( .A(n2008), .Z(n1544) );
  INV_X1 U1509 ( .A(n1545), .ZN(n1546) );
  INV_X1 U1510 ( .A(n2467), .ZN(n1547) );
  BUF_X1 U1511 ( .A(n3506), .Z(n1548) );
  OAI211_X1 U1512 ( .C1(n2566), .C2(n2175), .A(n3306), .B(n1721), .ZN(
        \DataP/alu_b_in[25] ) );
  AOI21_X1 U1513 ( .B1(n1541), .B2(n3691), .A(n3454), .ZN(n1549) );
  AND4_X2 U1514 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n1550)
         );
  INV_X4 U1515 ( .A(n1550), .ZN(\DataP/alu_b_in[24] ) );
  NAND2_X1 U1516 ( .A1(n3427), .A2(n3510), .ZN(n1551) );
  INV_X2 U1517 ( .A(n1945), .ZN(n1553) );
  AND3_X1 U1518 ( .A1(n1620), .A2(n2314), .A3(n1617), .ZN(n1554) );
  AND4_X1 U1519 ( .A1(n3063), .A2(n3062), .A3(n3027), .A4(n3028), .ZN(n1555)
         );
  AND4_X1 U1520 ( .A1(n3063), .A2(n3062), .A3(n3027), .A4(n3028), .ZN(n3029)
         );
  AND4_X1 U1521 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n1556)
         );
  INV_X2 U1522 ( .A(n1556), .ZN(\DataP/alu_b_in[20] ) );
  AND3_X1 U1523 ( .A1(n1620), .A2(n2314), .A3(n1617), .ZN(n2313) );
  NAND2_X1 U1524 ( .A1(n1551), .A2(n1558), .ZN(n1557) );
  AND2_X1 U1525 ( .A1(n1884), .A2(n2297), .ZN(n1558) );
  AND2_X1 U1526 ( .A1(n2378), .A2(n1552), .ZN(n1559) );
  AND2_X1 U1527 ( .A1(n2378), .A2(n1552), .ZN(n1877) );
  AND2_X2 U1528 ( .A1(n3424), .A2(n3425), .ZN(n2245) );
  NAND2_X1 U1529 ( .A1(n2007), .A2(\DataP/alu_a_in[20] ), .ZN(n1560) );
  OAI21_X1 U1530 ( .B1(n1567), .B2(n121), .A(n3115), .ZN(n1562) );
  OR2_X2 U1531 ( .A1(n1562), .A2(n3116), .ZN(\DataP/alu_a_in[1] ) );
  AND2_X2 U1532 ( .A1(n3420), .A2(n3421), .ZN(n1563) );
  AND4_X1 U1533 ( .A1(n3305), .A2(n2519), .A3(n3303), .A4(n3304), .ZN(n1580)
         );
  OR2_X2 U1534 ( .A1(n3184), .A2(n3183), .ZN(\DataP/alu_a_in[13] ) );
  INV_X2 U1535 ( .A(n2005), .ZN(n3002) );
  AND2_X2 U1536 ( .A1(n2315), .A2(n1554), .ZN(n2005) );
  NAND2_X1 U1537 ( .A1(n1518), .A2(\DataP/B_s[0] ), .ZN(n1564) );
  NAND4_X1 U1538 ( .A1(n1861), .A2(n3030), .A3(n2472), .A4(n2471), .ZN(n1565)
         );
  NAND4_X1 U1539 ( .A1(n1861), .A2(n3030), .A3(n2472), .A4(n2471), .ZN(n3046)
         );
  NAND3_X1 U1540 ( .A1(n3029), .A2(n2472), .A3(n3030), .ZN(n1566) );
  NOR2_X2 U1541 ( .A1(n1596), .A2(n1595), .ZN(n3030) );
  NAND3_X1 U1542 ( .A1(n1568), .A2(n2998), .A3(n2155), .ZN(n1567) );
  INV_X1 U1543 ( .A(n3191), .ZN(n1568) );
  AND3_X2 U1544 ( .A1(n3104), .A2(n1525), .A3(n3107), .ZN(n1569) );
  INV_X2 U1545 ( .A(\DataP/alu_b_in[8] ), .ZN(n3663) );
  NAND2_X2 U1546 ( .A1(n1570), .A2(n1571), .ZN(n1572) );
  AND2_X1 U1547 ( .A1(n3244), .A2(n3245), .ZN(n1570) );
  AND2_X1 U1548 ( .A1(n3246), .A2(n3247), .ZN(n1571) );
  OR2_X2 U1549 ( .A1(n3155), .A2(n3154), .ZN(\DataP/alu_a_in[23] ) );
  AOI211_X1 U1550 ( .C1(\DataP/alu_a_in[28] ), .C2(n1917), .A(n2067), .B(n2048), .ZN(n1573) );
  INV_X1 U1551 ( .A(n1575), .ZN(n3104) );
  AND2_X1 U1552 ( .A1(n3004), .A2(\DataP/alu_out_W[5] ), .ZN(n1575) );
  AOI21_X1 U1553 ( .B1(n2325), .B2(n2130), .A(n1948), .ZN(n1574) );
  CLKBUF_X3 U1554 ( .A(\DataP/alu_b_in[5] ), .Z(\lt_x_134/B[5] ) );
  AOI211_X4 U1555 ( .C1(n2047), .C2(n2107), .A(n2105), .B(n1810), .ZN(n2057)
         );
  NAND2_X1 U1556 ( .A1(n1576), .A2(n3048), .ZN(n2389) );
  AND2_X1 U1557 ( .A1(n3047), .A2(n2391), .ZN(n1576) );
  AND2_X2 U1558 ( .A1(n1900), .A2(n1637), .ZN(n1577) );
  AND2_X2 U1559 ( .A1(n1578), .A2(n1579), .ZN(n3417) );
  AND3_X1 U1560 ( .A1(n3301), .A2(n3300), .A3(n3302), .ZN(n1578) );
  NAND2_X1 U1561 ( .A1(n1839), .A2(\DataP/B_s[15] ), .ZN(n1579) );
  NAND4_X1 U1562 ( .A1(n3095), .A2(n3093), .A3(n3092), .A4(n3094), .ZN(n1581)
         );
  NAND2_X1 U1563 ( .A1(n1584), .A2(n1583), .ZN(n1582) );
  AND2_X1 U1564 ( .A1(n1585), .A2(n2332), .ZN(n1583) );
  NAND2_X1 U1565 ( .A1(n2331), .A2(DRAM_ADDRESS[8]), .ZN(n1584) );
  NAND2_X1 U1566 ( .A1(n1518), .A2(\DataP/B_s[8] ), .ZN(n1585) );
  BUF_X4 U1567 ( .A(n2712), .Z(n2709) );
  NAND2_X2 U1568 ( .A1(n3224), .A2(n3343), .ZN(n3689) );
  NOR2_X2 U1569 ( .A1(ALU_OPCODE_i[3]), .A2(ALU_OPCODE_i[0]), .ZN(n3343) );
  AND3_X2 U1570 ( .A1(n2442), .A2(n1994), .A3(n2010), .ZN(n3421) );
  OR2_X2 U1571 ( .A1(n3164), .A2(n3163), .ZN(\DataP/alu_a_in[20] ) );
  AND3_X2 U1572 ( .A1(n1998), .A2(n3460), .A3(n3457), .ZN(n3494) );
  INV_X1 U1573 ( .A(n2145), .ZN(n1586) );
  NAND2_X1 U1574 ( .A1(n1993), .A2(n3678), .ZN(n1587) );
  OR2_X2 U1575 ( .A1(n3149), .A2(n3148), .ZN(\DataP/alu_a_in[25] ) );
  OR2_X2 U1576 ( .A1(n3003), .A2(n2234), .ZN(n3089) );
  AND2_X1 U1577 ( .A1(n3021), .A2(n3022), .ZN(n1588) );
  NOR2_X1 U1578 ( .A1(n3161), .A2(n3160), .ZN(n1589) );
  AND4_X1 U1579 ( .A1(n3087), .A2(n3085), .A3(n3086), .A4(n3084), .ZN(n1907)
         );
  NAND3_X1 U1580 ( .A1(n3101), .A2(n3100), .A3(n3102), .ZN(n1625) );
  OR2_X1 U1581 ( .A1(n2389), .A2(n1846), .ZN(\DataP/alu_b_in[9] ) );
  XOR2_X1 U1582 ( .A(n3011), .B(n3203), .Z(n1957) );
  BUF_X1 U1583 ( .A(n3532), .Z(n1590) );
  BUF_X1 U1584 ( .A(n1531), .Z(n1591) );
  NOR3_X1 U1585 ( .A1(n1582), .A2(n2389), .A3(n2333), .ZN(n1592) );
  AND2_X2 U1586 ( .A1(n1569), .A2(n1843), .ZN(n1994) );
  NAND2_X2 U1587 ( .A1(n3464), .A2(\DataP/alu_a_in[23] ), .ZN(n3497) );
  BUF_X2 U1588 ( .A(\DataP/alu_b_in[12] ), .Z(n1880) );
  NOR2_X2 U1589 ( .A1(n3639), .A2(n1962), .ZN(n2225) );
  OAI21_X1 U1590 ( .B1(n309), .B2(n3911), .A(n1593), .ZN(\DataP/PC_reg/N25 )
         );
  OR2_X1 U1591 ( .A1(n3910), .A2(n4013), .ZN(n1593) );
  OAI21_X2 U1592 ( .B1(n2434), .B2(n3911), .A(n1523), .ZN(n2346) );
  BUF_X2 U1593 ( .A(n3327), .Z(n1839) );
  NAND3_X1 U1594 ( .A1(n1555), .A2(n2472), .A3(n3030), .ZN(n2315) );
  NOR2_X1 U1595 ( .A1(n3024), .A2(n3025), .ZN(n3028) );
  NAND3_X1 U1596 ( .A1(n1994), .A2(n2442), .A3(n1903), .ZN(n2440) );
  AND3_X1 U1597 ( .A1(n3067), .A2(n3066), .A3(n432), .ZN(n2143) );
  AND4_X2 U1598 ( .A1(n1577), .A2(n2501), .A3(n1569), .A4(n1624), .ZN(n3207)
         );
  NAND2_X1 U1599 ( .A1(n2331), .A2(\DataP/alu_out_M[18] ), .ZN(n1594) );
  NAND2_X1 U1600 ( .A1(n3020), .A2(n3019), .ZN(n1595) );
  AOI21_X1 U1601 ( .B1(n1597), .B2(n3017), .A(n3049), .ZN(n1596) );
  NAND2_X1 U1602 ( .A1(n1953), .A2(\DataP/opcode_W[5] ), .ZN(n3017) );
  AND2_X1 U1603 ( .A1(n3016), .A2(\DataP/opcode_W[3] ), .ZN(n1597) );
  OAI211_X1 U1604 ( .C1(\DataP/opcode_W[4] ), .C2(\DataP/opcode_W[0] ), .A(
        \DataP/opcode_W[2] ), .B(\DataP/opcode_W[1] ), .ZN(n3016) );
  OR2_X4 U1605 ( .A1(n3110), .A2(n3109), .ZN(\DataP/alu_a_in[3] ) );
  OR2_X2 U1606 ( .A1(n3181), .A2(n3180), .ZN(\DataP/alu_a_in[14] ) );
  AND4_X1 U1607 ( .A1(n3262), .A2(n2390), .A3(n3419), .A4(n3263), .ZN(n1598)
         );
  AND4_X1 U1608 ( .A1(n3262), .A2(n3419), .A3(n2390), .A4(n1896), .ZN(n3420)
         );
  AOI21_X1 U1609 ( .B1(n3542), .B2(n3691), .A(n3541), .ZN(n1599) );
  XNOR2_X1 U1610 ( .A(n1959), .B(n1600), .ZN(n3621) );
  AND2_X2 U1611 ( .A1(n3611), .A2(n1757), .ZN(n1600) );
  OR2_X1 U1612 ( .A1(n1997), .A2(n2244), .ZN(n1601) );
  OR2_X1 U1613 ( .A1(n1997), .A2(n2244), .ZN(n3641) );
  BUF_X1 U1614 ( .A(n1983), .Z(n1602) );
  NOR2_X1 U1615 ( .A1(n1911), .A2(n1965), .ZN(n1603) );
  AOI21_X1 U1616 ( .B1(n3621), .B2(n3691), .A(n3620), .ZN(n1604) );
  BUF_X2 U1617 ( .A(\DataP/alu_a_in[0] ), .Z(n1605) );
  NAND2_X1 U1618 ( .A1(n2425), .A2(n2540), .ZN(n1606) );
  OAI21_X1 U1619 ( .B1(n1957), .B2(n1918), .A(n2366), .ZN(n1607) );
  OR2_X2 U1620 ( .A1(n3050), .A2(n1865), .ZN(n2472) );
  AND4_X2 U1621 ( .A1(n1847), .A2(n3028), .A3(n3027), .A4(n3062), .ZN(n1861)
         );
  NOR2_X1 U1622 ( .A1(\DataP/alu_b_in[3] ), .A2(\DataP/alu_b_in[2] ), .ZN(
        n1608) );
  OR2_X1 U1623 ( .A1(n3692), .A2(n3674), .ZN(n1609) );
  INV_X1 U1624 ( .A(n1530), .ZN(n1932) );
  NOR2_X2 U1625 ( .A1(n2555), .A2(n2554), .ZN(n2552) );
  BUF_X1 U1626 ( .A(n1552), .Z(n1610) );
  NAND4_X2 U1627 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(
        \DataP/alu_b_in[21] ) );
  INV_X1 U1628 ( .A(\DataP/alu_b_in[6] ), .ZN(n1611) );
  NOR2_X1 U1629 ( .A1(n1911), .A2(n1965), .ZN(n2362) );
  INV_X1 U1630 ( .A(n1907), .ZN(n1612) );
  NAND2_X1 U1631 ( .A1(n3677), .A2(n3678), .ZN(n3676) );
  NAND2_X1 U1632 ( .A1(n1613), .A2(n3370), .ZN(n3677) );
  NAND2_X1 U1633 ( .A1(n3372), .A2(n3371), .ZN(n1613) );
  NAND2_X1 U1634 ( .A1(n1561), .A2(n2419), .ZN(n3371) );
  NAND2_X1 U1635 ( .A1(n1816), .A2(n3359), .ZN(n3372) );
  NAND2_X1 U1636 ( .A1(n1619), .A2(n1614), .ZN(n3065) );
  AND2_X1 U1637 ( .A1(n1618), .A2(n1616), .ZN(n1614) );
  NOR2_X1 U1638 ( .A1(n2573), .A2(n2468), .ZN(n1615) );
  NAND2_X1 U1639 ( .A1(n3038), .A2(n3039), .ZN(n1620) );
  OAI211_X1 U1640 ( .C1(n3033), .C2(\DataP/opcode_M[4] ), .A(n1622), .B(n1621), 
        .ZN(n3039) );
  AOI21_X1 U1641 ( .B1(n1543), .B2(\DataP/opcode_M[4] ), .A(
        \DataP/opcode_M[5] ), .ZN(n1621) );
  INV_X1 U1642 ( .A(n3032), .ZN(n1622) );
  NAND2_X1 U1643 ( .A1(n1623), .A2(\DataP/opcode_M[3] ), .ZN(n3038) );
  OAI21_X1 U1644 ( .B1(n3036), .B2(n146), .A(n3035), .ZN(n1623) );
  NOR2_X1 U1645 ( .A1(n1626), .A2(n1625), .ZN(n1624) );
  INV_X1 U1646 ( .A(n3103), .ZN(n1626) );
  OAI21_X1 U1647 ( .B1(n150), .B2(\DataP/opcode_M[1] ), .A(n1627), .ZN(n3032)
         );
  NAND2_X1 U1648 ( .A1(\DataP/opcode_M[1] ), .A2(\DataP/opcode_M[3] ), .ZN(
        n1627) );
  INV_X1 U1649 ( .A(n2243), .ZN(n1632) );
  OAI211_X1 U1650 ( .C1(n1544), .C2(n1633), .A(n1629), .B(n1628), .ZN(n2418)
         );
  NAND3_X1 U1651 ( .A1(n2008), .A2(n2430), .A3(n1632), .ZN(n1628) );
  INV_X1 U1652 ( .A(n1630), .ZN(n1629) );
  OAI21_X1 U1653 ( .B1(n2430), .B2(n1633), .A(n1631), .ZN(n1630) );
  NAND2_X2 U1654 ( .A1(n1632), .A2(n2426), .ZN(n1631) );
  NAND2_X2 U1655 ( .A1(n2515), .A2(n2243), .ZN(n1633) );
  NAND2_X1 U1656 ( .A1(n1634), .A2(n1980), .ZN(\DataP/PC_reg/N31 ) );
  NAND2_X1 U1657 ( .A1(n2418), .A2(n1982), .ZN(n1634) );
  NAND4_X1 U1658 ( .A1(n3095), .A2(n3093), .A3(n3092), .A4(n3094), .ZN(
        \DataP/alu_b_in[3] ) );
  BUF_X1 U1659 ( .A(n3327), .Z(n1635) );
  INV_X1 U1660 ( .A(n2331), .ZN(n1636) );
  AND3_X1 U1661 ( .A1(n3087), .A2(n3090), .A3(n3089), .ZN(n1637) );
  OAI21_X1 U1662 ( .B1(n2380), .B2(n2577), .A(n2379), .ZN(n1638) );
  BUF_X1 U1663 ( .A(n3565), .Z(n1639) );
  INV_X1 U1664 ( .A(n2130), .ZN(\sra_131/SH[4] ) );
  AND4_X1 U1665 ( .A1(n3673), .A2(n3681), .A3(n3380), .A4(n3316), .ZN(n1856)
         );
  OR2_X1 U1666 ( .A1(n3003), .A2(n2233), .ZN(n3085) );
  BUF_X2 U1667 ( .A(n1887), .Z(n1837) );
  BUF_X1 U1668 ( .A(n3612), .Z(n1959) );
  OR2_X1 U1669 ( .A1(n3512), .A2(n2539), .ZN(n2226) );
  INV_X1 U1670 ( .A(n2450), .ZN(n1976) );
  INV_X2 U1671 ( .A(n2845), .ZN(n2846) );
  INV_X1 U1672 ( .A(n2048), .ZN(n1640) );
  OAI22_X1 U1673 ( .A1(\DataP/alu_b_in[31] ), .A2(n1923), .B1(
        \DataP/alu_a_in[30] ), .B2(n2053), .ZN(n1641) );
  AOI211_X1 U1674 ( .C1(n2055), .C2(n1640), .A(n2054), .B(n1641), .ZN(n2056)
         );
  INV_X1 U1675 ( .A(\lt_x_135/B[4] ), .ZN(n1642) );
  OAI21_X1 U1676 ( .B1(n3671), .B2(n1642), .A(n3694), .ZN(n1643) );
  AOI22_X1 U1677 ( .A1(\DataP/alu_a_in[4] ), .A2(n1643), .B1(\lt_x_134/B[4] ), 
        .B2(n3697), .ZN(n3672) );
  OAI21_X1 U1678 ( .B1(n2065), .B2(n2984), .A(n2980), .ZN(n1644) );
  INV_X1 U1679 ( .A(\lt_x_134/B[4] ), .ZN(n1645) );
  INV_X1 U1680 ( .A(\lt_x_135/B[4] ), .ZN(n1646) );
  OAI221_X1 U1681 ( .B1(\lt_x_135/B[4] ), .B2(n2837), .C1(n1646), .C2(n2836), 
        .A(n3006), .ZN(n1647) );
  NAND2_X1 U1682 ( .A1(n1645), .A2(n3007), .ZN(n1648) );
  OAI21_X1 U1683 ( .B1(n2708), .B2(n1648), .A(n1647), .ZN(n1649) );
  AOI21_X1 U1684 ( .B1(n3659), .B2(n3656), .A(n3217), .ZN(n1650) );
  NAND2_X1 U1685 ( .A1(n3232), .A2(n3266), .ZN(n1651) );
  AOI21_X1 U1686 ( .B1(n1650), .B2(n1651), .A(n3674), .ZN(n1652) );
  OAI21_X1 U1687 ( .B1(n1650), .B2(n1651), .A(n1652), .ZN(n1653) );
  OAI211_X1 U1688 ( .C1(n3700), .C2(n3282), .A(n3228), .B(n1653), .ZN(n1654)
         );
  AOI211_X1 U1689 ( .C1(n3675), .C2(n1644), .A(n1649), .B(n1654), .ZN(n341) );
  NAND4_X1 U1690 ( .A1(n2467), .A2(n1550), .A3(n2503), .A4(n2133), .ZN(n1655)
         );
  OAI211_X1 U1691 ( .C1(n2467), .C2(n2133), .A(n2367), .B(n1655), .ZN(n1656)
         );
  NAND2_X1 U1692 ( .A1(n1547), .A2(n2321), .ZN(n1657) );
  OAI21_X1 U1693 ( .B1(n2368), .B2(n1656), .A(n1657), .ZN(n3470) );
  OAI21_X1 U1694 ( .B1(n2847), .B2(n2983), .A(n2977), .ZN(n1658) );
  OAI22_X1 U1695 ( .A1(n3663), .A2(n3664), .B1(n1921), .B2(n3662), .ZN(n1659)
         );
  INV_X1 U1696 ( .A(\lt_x_134/B[4] ), .ZN(n1660) );
  OAI221_X1 U1697 ( .B1(\lt_x_134/B[4] ), .B2(n2833), .C1(n1660), .C2(n2832), 
        .A(n3703), .ZN(n1661) );
  NOR2_X1 U1698 ( .A1(\lt_x_135/B[4] ), .A2(n2707), .ZN(n1662) );
  XNOR2_X1 U1699 ( .A(\DataP/alu_a_in[8] ), .B(n3658), .ZN(n1663) );
  AOI21_X1 U1700 ( .B1(n3657), .B2(n3656), .A(n3659), .ZN(n1664) );
  AOI211_X1 U1701 ( .C1(n3659), .C2(n1663), .A(n1664), .B(n3674), .ZN(n1665)
         );
  AOI21_X1 U1702 ( .B1(n3706), .B2(n1662), .A(n1665), .ZN(n1666) );
  NAND2_X1 U1703 ( .A1(n1661), .A2(n1666), .ZN(n1667) );
  AOI211_X1 U1704 ( .C1(n3675), .C2(n1658), .A(n1659), .B(n1667), .ZN(n345) );
  NAND3_X1 U1705 ( .A1(n3488), .A2(n3509), .A3(n1917), .ZN(n1668) );
  XOR2_X1 U1706 ( .A(\DataP/alu_b_in[29] ), .B(n1668), .Z(n2371) );
  NAND2_X1 U1707 ( .A1(n2565), .A2(\DataP/IMM_s[18] ), .ZN(n1669) );
  NAND2_X1 U1708 ( .A1(n2564), .A2(\DataP/ir_E[14] ), .ZN(n1670) );
  NAND3_X1 U1709 ( .A1(n1670), .A2(n3312), .A3(n3311), .ZN(n1671) );
  AOI21_X1 U1710 ( .B1(n3001), .B2(\DataP/B_s[14] ), .A(n1671), .ZN(n3418) );
  XOR2_X1 U1711 ( .A(n3665), .B(n1851), .Z(n1672) );
  AOI22_X1 U1712 ( .A1(n1915), .A2(n2823), .B1(n2064), .B2(n2822), .ZN(n1673)
         );
  INV_X1 U1713 ( .A(\lt_x_135/B[4] ), .ZN(n1674) );
  OAI221_X1 U1714 ( .B1(\lt_x_135/B[4] ), .B2(n1673), .C1(n1674), .C2(n2824), 
        .A(n3703), .ZN(n1675) );
  INV_X1 U1715 ( .A(n2968), .ZN(n1676) );
  INV_X1 U1716 ( .A(n2065), .ZN(n1677) );
  OAI221_X1 U1717 ( .B1(n2065), .B2(n1676), .C1(n1677), .C2(n2967), .A(n3675), 
        .ZN(n1678) );
  OAI211_X1 U1718 ( .C1(n1672), .C2(n3674), .A(n1675), .B(n1678), .ZN(n1679)
         );
  AOI21_X1 U1719 ( .B1(n3667), .B2(n3694), .A(n2363), .ZN(n1680) );
  AOI21_X1 U1720 ( .B1(n3697), .B2(\DataP/alu_a_in[6] ), .A(n1680), .ZN(n1681)
         );
  NAND3_X1 U1721 ( .A1(n3007), .A2(n2693), .A3(n1674), .ZN(n1682) );
  OAI211_X1 U1722 ( .C1(n3700), .C2(n3668), .A(n1681), .B(n1682), .ZN(n1683)
         );
  NOR2_X1 U1723 ( .A1(n1679), .A2(n1683), .ZN(n353) );
  AOI22_X1 U1724 ( .A1(n3005), .A2(\DataP/alu_out_W[26] ), .B1(n3001), .B2(
        \DataP/B_s[26] ), .ZN(n1684) );
  OAI211_X1 U1725 ( .C1(n1636), .C2(n2169), .A(n3306), .B(n1684), .ZN(
        \DataP/alu_b_in[26] ) );
  AOI22_X1 U1726 ( .A1(\DataP/alu_a_in[5] ), .A2(n3379), .B1(\lt_x_134/B[5] ), 
        .B2(n3697), .ZN(n1685) );
  INV_X1 U1727 ( .A(\lt_x_134/B[4] ), .ZN(n1686) );
  NAND3_X1 U1728 ( .A1(n3007), .A2(n2692), .A3(n1686), .ZN(n1687) );
  OAI211_X1 U1729 ( .C1(n3380), .C2(n3700), .A(n1685), .B(n1687), .ZN(n1688)
         );
  NAND2_X1 U1730 ( .A1(n1899), .A2(n3382), .ZN(n1689) );
  XNOR2_X1 U1731 ( .A(n1689), .B(n3383), .ZN(n1690) );
  AOI22_X1 U1732 ( .A1(n2064), .A2(n2817), .B1(n1915), .B2(n2818), .ZN(n1691)
         );
  OAI221_X1 U1733 ( .B1(\lt_x_134/B[4] ), .B2(n1691), .C1(n1686), .C2(n2819), 
        .A(n3006), .ZN(n1692) );
  OAI21_X1 U1734 ( .B1(n2065), .B2(n2963), .A(n2962), .ZN(n1693) );
  NAND2_X1 U1735 ( .A1(n1693), .A2(n3675), .ZN(n1694) );
  OAI211_X1 U1736 ( .C1(n3674), .C2(n1690), .A(n1692), .B(n1694), .ZN(n1695)
         );
  NOR2_X1 U1737 ( .A1(n1688), .A2(n1695), .ZN(n354) );
  INV_X1 U1738 ( .A(n3392), .ZN(n1696) );
  NAND3_X1 U1739 ( .A1(n3510), .A2(n1841), .A3(n1696), .ZN(n3416) );
  AOI22_X1 U1740 ( .A1(n2846), .A2(n2635), .B1(n2127), .B2(n2687), .ZN(n1697)
         );
  INV_X1 U1741 ( .A(\lt_x_135/B[4] ), .ZN(n1698) );
  OAI221_X1 U1742 ( .B1(\lt_x_135/B[4] ), .B2(n1697), .C1(n1698), .C2(n2694), 
        .A(n3706), .ZN(n3451) );
  AND3_X2 U1743 ( .A1(n2245), .A2(n2306), .A3(n1522), .ZN(n2136) );
  AOI21_X1 U1744 ( .B1(n2301), .B2(n2300), .A(n2183), .ZN(n1699) );
  OAI211_X1 U1745 ( .C1(n1946), .C2(\DataP/alu_b_in[18] ), .A(n3426), .B(n2496), .ZN(n1700) );
  NAND2_X1 U1746 ( .A1(n1932), .A2(n2478), .ZN(n1701) );
  NAND2_X1 U1747 ( .A1(n3510), .A2(n2377), .ZN(n1702) );
  NAND2_X1 U1748 ( .A1(n3400), .A2(n2372), .ZN(n1703) );
  OAI211_X1 U1749 ( .C1(n1702), .C2(n3400), .A(n1703), .B(n1701), .ZN(n3401)
         );
  AOI22_X1 U1750 ( .A1(n3005), .A2(\DataP/alu_out_W[30] ), .B1(\DataP/B_s[30] ), .B2(n1859), .ZN(n1704) );
  OAI211_X1 U1751 ( .C1(n2566), .C2(n2187), .A(n3306), .B(n1704), .ZN(
        \DataP/alu_b_in[30] ) );
  NOR2_X1 U1752 ( .A1(\lt_x_134/B[4] ), .A2(n2705), .ZN(n1705) );
  XNOR2_X1 U1753 ( .A(\DataP/alu_a_in[4] ), .B(n3670), .ZN(n1706) );
  XNOR2_X1 U1754 ( .A(n1706), .B(n1961), .ZN(n1707) );
  OAI21_X1 U1755 ( .B1(n2847), .B2(n2956), .A(n2955), .ZN(n1708) );
  NAND2_X1 U1756 ( .A1(n1708), .A2(n3675), .ZN(n1709) );
  OAI21_X1 U1757 ( .B1(n3674), .B2(n1707), .A(n1709), .ZN(n1710) );
  OAI221_X1 U1758 ( .B1(\lt_x_134/B[4] ), .B2(n2814), .C1(n1645), .C2(n2813), 
        .A(n3703), .ZN(n1711) );
  OAI211_X1 U1759 ( .C1(n3673), .C2(n3700), .A(n3672), .B(n1711), .ZN(n1712)
         );
  AOI211_X1 U1760 ( .C1(n3007), .C2(n1705), .A(n1710), .B(n1712), .ZN(n355) );
  AOI21_X1 U1761 ( .B1(n2478), .B2(n2407), .A(\DataP/alu_a_in[29] ), .ZN(n2279) );
  XNOR2_X1 U1762 ( .A(\DataP/alu_a_in[8] ), .B(n3663), .ZN(n1713) );
  AOI211_X1 U1763 ( .C1(n3335), .C2(n3317), .A(n3402), .B(n1713), .ZN(n1714)
         );
  AND3_X1 U1764 ( .A1(n2452), .A2(n1714), .A3(n3668), .ZN(n1853) );
  OAI21_X1 U1765 ( .B1(n2573), .B2(n151), .A(\DataP/opcode_E[4] ), .ZN(n1715)
         );
  AND2_X1 U1766 ( .A1(\DataP/opcode_E[3] ), .A2(n2573), .ZN(n1716) );
  OAI33_X1 U1767 ( .A1(n1715), .A2(n2575), .A3(n1716), .B1(\DataP/opcode_E[4] ), .B2(\DataP/opcode_E[0] ), .B3(n149), .ZN(n1717) );
  AOI21_X1 U1768 ( .B1(n3060), .B2(\DataP/opcode_E[4] ), .A(n145), .ZN(n1718)
         );
  OAI21_X1 U1769 ( .B1(n521), .B2(n520), .A(\DataP/opcode_E[3] ), .ZN(n1719)
         );
  NOR2_X1 U1770 ( .A1(n1718), .A2(n1719), .ZN(n1720) );
  AOI21_X1 U1771 ( .B1(n145), .B2(n1717), .A(n1720), .ZN(n3073) );
  AOI22_X1 U1772 ( .A1(n3001), .A2(\DataP/B_s[25] ), .B1(n3005), .B2(
        \DataP/alu_out_W[25] ), .ZN(n1721) );
  NAND4_X1 U1773 ( .A1(n1882), .A2(n3458), .A3(n2526), .A4(n2540), .ZN(n2424)
         );
  AOI22_X1 U1774 ( .A1(n2843), .A2(n2826), .B1(n2844), .B2(n2825), .ZN(n1722)
         );
  AOI22_X1 U1775 ( .A1(n1915), .A2(n2827), .B1(n2845), .B2(n1722), .ZN(n2829)
         );
  NOR2_X1 U1776 ( .A1(n3510), .A2(n2279), .ZN(n1723) );
  NAND2_X1 U1777 ( .A1(n2281), .A2(n2279), .ZN(n1724) );
  OAI211_X1 U1778 ( .C1(n2371), .C2(n1723), .A(n2280), .B(n1724), .ZN(n2513)
         );
  NOR2_X1 U1779 ( .A1(n2177), .A2(n2566), .ZN(n1725) );
  AOI21_X1 U1780 ( .B1(n1515), .B2(\DataP/ir_E[12] ), .A(n1725), .ZN(n1726) );
  NAND3_X1 U1781 ( .A1(n1726), .A2(n3261), .A3(n2387), .ZN(
        \DataP/alu_b_in[12] ) );
  NOR2_X1 U1782 ( .A1(n3249), .A2(n1879), .ZN(n1727) );
  XNOR2_X1 U1783 ( .A(n1727), .B(n1572), .ZN(n3251) );
  OAI221_X1 U1784 ( .B1(n2122), .B2(n2120), .C1(n2122), .C2(n2121), .A(n2119), 
        .ZN(n1728) );
  MUX2_X1 U1785 ( .A(n1983), .B(n1728), .S(ALU_OPCODE_i[2]), .Z(n3346) );
  NOR2_X1 U1786 ( .A1(n2713), .A2(n2578), .ZN(n1729) );
  AOI22_X1 U1787 ( .A1(n2599), .A2(n1930), .B1(n2842), .B2(n1729), .ZN(n2622)
         );
  AOI22_X1 U1788 ( .A1(n3423), .A2(n1520), .B1(n2002), .B2(n1840), .ZN(n1730)
         );
  OAI21_X1 U1789 ( .B1(n1591), .B2(n1730), .A(n1960), .ZN(n3428) );
  OAI21_X1 U1790 ( .B1(\DataP/alu_a_in[25] ), .B2(n1547), .A(n3697), .ZN(n1731) );
  NAND3_X1 U1791 ( .A1(\DataP/alu_a_in[25] ), .A2(n1547), .A3(n3693), .ZN(
        n1732) );
  OAI211_X1 U1792 ( .C1(n3547), .C2(n3700), .A(n1731), .B(n1732), .ZN(n3548)
         );
  AOI22_X1 U1793 ( .A1(n2508), .A2(n2003), .B1(n3689), .B2(n3663), .ZN(n1733)
         );
  NAND3_X1 U1794 ( .A1(n2509), .A2(n2507), .A3(n1733), .ZN(n3658) );
  OAI21_X1 U1795 ( .B1(n2065), .B2(n2949), .A(n2948), .ZN(n1734) );
  AOI22_X1 U1796 ( .A1(n1916), .A2(n2805), .B1(n2840), .B2(n2806), .ZN(n1735)
         );
  AOI22_X1 U1797 ( .A1(n2842), .A2(n2825), .B1(n1930), .B2(n1735), .ZN(n1736)
         );
  AOI22_X1 U1798 ( .A1(n2330), .A2(n1736), .B1(n2846), .B2(n2807), .ZN(n1737)
         );
  INV_X1 U1799 ( .A(\lt_x_135/B[4] ), .ZN(n1738) );
  OAI221_X1 U1800 ( .B1(\lt_x_135/B[4] ), .B2(n1737), .C1(n1738), .C2(n2808), 
        .A(n3006), .ZN(n1739) );
  INV_X1 U1801 ( .A(n2690), .ZN(n1740) );
  AOI22_X1 U1802 ( .A1(\DataP/alu_a_in[3] ), .A2(n3680), .B1(n1963), .B2(n3697), .ZN(n1741) );
  OAI211_X1 U1803 ( .C1(n3678), .C2(n1993), .A(n2001), .B(n3691), .ZN(n1742)
         );
  OAI211_X1 U1804 ( .C1(n3700), .C2(n3681), .A(n1741), .B(n1742), .ZN(n1743)
         );
  NOR2_X1 U1805 ( .A1(n1740), .A2(\lt_x_134/B[4] ), .ZN(n1744) );
  AOI21_X1 U1806 ( .B1(n1744), .B2(n3706), .A(n1743), .ZN(n1745) );
  NAND2_X1 U1807 ( .A1(n1745), .A2(n1739), .ZN(n1746) );
  AOI21_X1 U1808 ( .B1(n3675), .B2(n1734), .A(n1746), .ZN(n356) );
  OAI21_X1 U1809 ( .B1(n1589), .B2(\DataP/alu_b_in[21] ), .A(
        \DataP/alu_b_in[20] ), .ZN(n1747) );
  OAI22_X1 U1810 ( .A1(\DataP/alu_a_in[20] ), .A2(n1747), .B1(
        \DataP/alu_a_in[21] ), .B2(n1952), .ZN(n2107) );
  INV_X1 U1811 ( .A(n1838), .ZN(n1748) );
  NAND2_X1 U1812 ( .A1(n2493), .A2(n3510), .ZN(n1749) );
  AOI21_X1 U1813 ( .B1(n2538), .B2(n1749), .A(n1748), .ZN(n2491) );
  NAND2_X1 U1814 ( .A1(n1947), .A2(n1881), .ZN(n1750) );
  NAND2_X1 U1815 ( .A1(n1932), .A2(n1750), .ZN(n2377) );
  INV_X1 U1816 ( .A(n1605), .ZN(n1751) );
  NAND2_X1 U1817 ( .A1(n2985), .A2(n1751), .ZN(n3335) );
  AND4_X1 U1818 ( .A1(n2476), .A2(n3058), .A3(n2477), .A4(n2163), .ZN(n1752)
         );
  NAND4_X1 U1819 ( .A1(n3062), .A2(n3064), .A3(n1752), .A4(n1883), .ZN(n3069)
         );
  AOI22_X1 U1820 ( .A1(n3005), .A2(\DataP/alu_out_W[29] ), .B1(n1859), .B2(
        \DataP/B_s[29] ), .ZN(n1753) );
  NAND2_X1 U1821 ( .A1(n2331), .A2(\DataP/alu_out_M[29] ), .ZN(n1754) );
  NAND3_X1 U1822 ( .A1(n1754), .A2(n1753), .A3(n3306), .ZN(
        \DataP/alu_b_in[29] ) );
  NAND3_X1 U1823 ( .A1(n3510), .A2(\DataP/alu_a_in[11] ), .A3(n3251), .ZN(
        n3272) );
  INV_X1 U1824 ( .A(n3202), .ZN(n1755) );
  NAND2_X1 U1825 ( .A1(\DataP/alu_a_in[3] ), .A2(n1755), .ZN(n3375) );
  OAI21_X1 U1826 ( .B1(\DataP/alu_b_in[22] ), .B2(n3510), .A(
        \DataP/alu_a_in[22] ), .ZN(n1756) );
  AOI21_X1 U1827 ( .B1(n3446), .B2(n3510), .A(n1756), .ZN(n2312) );
  NAND2_X1 U1828 ( .A1(n1986), .A2(n1878), .ZN(n1757) );
  OAI22_X1 U1829 ( .A1(n2989), .A2(n3694), .B1(n1561), .B2(n3373), .ZN(n1758)
         );
  NOR2_X1 U1830 ( .A1(\lt_x_135/B[4] ), .A2(n2704), .ZN(n1759) );
  NAND2_X1 U1831 ( .A1(n3370), .A2(n3371), .ZN(n1760) );
  XNOR2_X1 U1832 ( .A(n1760), .B(n3372), .ZN(n1761) );
  AOI22_X1 U1833 ( .A1(n1759), .A2(n3706), .B1(n1761), .B2(n3691), .ZN(n1762)
         );
  INV_X1 U1834 ( .A(n2937), .ZN(n1763) );
  INV_X1 U1835 ( .A(n2065), .ZN(n1764) );
  AOI22_X1 U1836 ( .A1(n2841), .A2(n2964), .B1(n2935), .B2(n2989), .ZN(n1765)
         );
  AOI22_X1 U1837 ( .A1(n2846), .A2(n2936), .B1(n2845), .B2(n1765), .ZN(n1766)
         );
  OAI221_X1 U1838 ( .B1(n2065), .B2(n1763), .C1(n1764), .C2(n1766), .A(n3675), 
        .ZN(n1767) );
  AOI22_X1 U1839 ( .A1(n2846), .A2(n2799), .B1(n2845), .B2(n2798), .ZN(n1768)
         );
  OAI221_X1 U1840 ( .B1(\lt_x_134/B[4] ), .B2(n1768), .C1(n1660), .C2(n2800), 
        .A(n3703), .ZN(n1769) );
  NAND3_X1 U1841 ( .A1(n1762), .A2(n1767), .A3(n1769), .ZN(n1770) );
  AOI211_X1 U1842 ( .C1(n3374), .C2(n1939), .A(n1758), .B(n1770), .ZN(n357) );
  XNOR2_X1 U1843 ( .A(n1946), .B(\DataP/alu_b_in[18] ), .ZN(n2300) );
  AOI22_X1 U1844 ( .A1(n2997), .A2(\DataP/alu_out_M[17] ), .B1(
        \DataP/alu_out_W[17] ), .B2(n2992), .ZN(n1771) );
  OAI21_X1 U1845 ( .B1(n57), .B2(n2999), .A(n1771), .ZN(n3172) );
  INV_X1 U1846 ( .A(n2109), .ZN(n1772) );
  AOI221_X1 U1847 ( .B1(n2123), .B2(n2117), .C1(n2116), .C2(n2117), .A(n2124), 
        .ZN(n1773) );
  OAI22_X1 U1848 ( .A1(\DataP/alu_a_in[31] ), .A2(n1935), .B1(
        \DataP/alu_a_in[30] ), .B2(n2118), .ZN(n1774) );
  INV_X1 U1849 ( .A(n3490), .ZN(n1775) );
  NAND2_X1 U1850 ( .A1(n3510), .A2(n1775), .ZN(n1776) );
  XNOR2_X1 U1851 ( .A(n1917), .B(n1776), .ZN(n3523) );
  OAI221_X1 U1852 ( .B1(n3510), .B2(n2358), .C1(n2383), .C2(n3233), .A(n3236), 
        .ZN(n3268) );
  AOI21_X1 U1853 ( .B1(n2383), .B2(n2382), .A(\DataP/alu_a_in[21] ), .ZN(n2379) );
  AOI21_X1 U1854 ( .B1(n3465), .B2(n2131), .A(n2421), .ZN(n1777) );
  NAND2_X1 U1855 ( .A1(n2422), .A2(n1777), .ZN(n3533) );
  AOI211_X1 U1856 ( .C1(n3353), .C2(n3352), .A(n2132), .B(ALU_OPCODE_i[0]), 
        .ZN(n1778) );
  AOI211_X1 U1857 ( .C1(n3353), .C2(\DataP/ALU_C/comp/N24 ), .A(
        ALU_OPCODE_i[1]), .B(n2150), .ZN(n1779) );
  OR2_X1 U1858 ( .A1(n1778), .A2(n1779), .ZN(n3354) );
  OAI221_X1 U1859 ( .B1(n1520), .B2(n3456), .C1(n1520), .C2(n2002), .A(n3423), 
        .ZN(n1987) );
  AND4_X1 U1860 ( .A1(n2477), .A2(n2476), .A3(n3058), .A4(n2163), .ZN(n1780)
         );
  AND3_X1 U1861 ( .A1(n3062), .A2(Rst), .A3(n1780), .ZN(n2475) );
  INV_X1 U1862 ( .A(n1899), .ZN(n1781) );
  AOI21_X1 U1863 ( .B1(n3382), .B2(n3383), .A(n1781), .ZN(n3665) );
  NOR2_X1 U1864 ( .A1(\DataP/alu_b_in[19] ), .A2(n1938), .ZN(n2496) );
  NAND2_X1 U1865 ( .A1(\DataP/alu_a_in[26] ), .A2(n1936), .ZN(n1782) );
  OAI21_X1 U1866 ( .B1(n1912), .B2(\DataP/alu_b_in[27] ), .A(n1782), .ZN(n2060) );
  AOI21_X1 U1867 ( .B1(n2478), .B2(n2512), .A(\DataP/alu_a_in[16] ), .ZN(n1979) );
  NOR2_X1 U1868 ( .A1(n3554), .A2(n2556), .ZN(n2131) );
  AOI22_X1 U1869 ( .A1(n3001), .A2(\DataP/B_s[23] ), .B1(n2565), .B2(
        \DataP/IMM_s[23] ), .ZN(n1783) );
  NAND2_X1 U1870 ( .A1(n3005), .A2(\DataP/alu_out_W[23] ), .ZN(n1784) );
  OAI211_X1 U1871 ( .C1(n1636), .C2(n2168), .A(n1783), .B(n1784), .ZN(
        \DataP/alu_b_in[23] ) );
  AOI22_X1 U1872 ( .A1(n2846), .A2(n2648), .B1(n2127), .B2(n2647), .ZN(n1785)
         );
  INV_X1 U1873 ( .A(\lt_x_135/B[4] ), .ZN(n1786) );
  OAI221_X1 U1874 ( .B1(\lt_x_135/B[4] ), .B2(n1785), .C1(n1786), .C2(n2618), 
        .A(n3007), .ZN(n3617) );
  AOI22_X1 U1875 ( .A1(n2842), .A2(n2652), .B1(n1913), .B2(n2677), .ZN(n1787)
         );
  AOI22_X1 U1876 ( .A1(n2127), .A2(n1787), .B1(n2653), .B2(n1915), .ZN(n1788)
         );
  OAI221_X1 U1877 ( .B1(\lt_x_134/B[4] ), .B2(n1788), .C1(n1686), .C2(n2654), 
        .A(n3007), .ZN(n3540) );
  OAI211_X1 U1878 ( .C1(n2321), .C2(n2365), .A(n2364), .B(n1944), .ZN(n3580)
         );
  INV_X1 U1879 ( .A(n1960), .ZN(n1789) );
  NOR2_X1 U1880 ( .A1(n1591), .A2(n1789), .ZN(n2572) );
  NAND3_X1 U1881 ( .A1(\DataP/alu_a_in[14] ), .A2(n1932), .A3(n3693), .ZN(
        n1790) );
  OAI21_X1 U1882 ( .B1(\DataP/alu_a_in[14] ), .B2(n1932), .A(n3697), .ZN(n1791) );
  OAI211_X1 U1883 ( .C1(n3633), .C2(n3700), .A(n1790), .B(n1791), .ZN(n3634)
         );
  NAND2_X1 U1884 ( .A1(n3657), .A2(n3266), .ZN(n1792) );
  INV_X1 U1885 ( .A(n3659), .ZN(n1793) );
  NAND2_X1 U1886 ( .A1(n3232), .A2(n1792), .ZN(n1794) );
  OAI21_X1 U1887 ( .B1(n1793), .B2(n3267), .A(n1794), .ZN(n3248) );
  AOI22_X1 U1888 ( .A1(n2127), .A2(n2978), .B1(n1915), .B2(n2979), .ZN(n1795)
         );
  NAND2_X1 U1889 ( .A1(n2065), .A2(n1795), .ZN(n2980) );
  AOI22_X1 U1890 ( .A1(n2064), .A2(n2975), .B1(n1915), .B2(n2976), .ZN(n1796)
         );
  NAND2_X1 U1891 ( .A1(n2065), .A2(n1796), .ZN(n2977) );
  AOI22_X1 U1892 ( .A1(n1914), .A2(\DataP/alu_a_in[2] ), .B1(n1931), .B2(
        \DataP/alu_a_in[1] ), .ZN(n1797) );
  AOI22_X1 U1893 ( .A1(\sra_131/SH[1] ), .A2(n2805), .B1(n1916), .B2(n1797), 
        .ZN(n2772) );
  AOI21_X1 U1894 ( .B1(n3050), .B2(n3049), .A(n1865), .ZN(n1798) );
  INV_X1 U1895 ( .A(n1798), .ZN(n3064) );
  INV_X1 U1896 ( .A(n3983), .ZN(n1799) );
  AOI221_X1 U1897 ( .B1(n3984), .B2(n3983), .C1(n3709), .C2(n1799), .A(n3982), 
        .ZN(\DataP/wrong_br ) );
  NOR2_X1 U1898 ( .A1(\lt_x_134/B[4] ), .A2(n2706), .ZN(n1800) );
  OAI21_X1 U1899 ( .B1(n3665), .B2(n3386), .A(n3385), .ZN(n1801) );
  XOR2_X1 U1900 ( .A(\DataP/alu_a_in[7] ), .B(n3213), .Z(n1802) );
  XNOR2_X1 U1901 ( .A(n1801), .B(n1802), .ZN(n1803) );
  NAND2_X1 U1902 ( .A1(\DataP/ALU_C/shifter/N89 ), .A2(n3675), .ZN(n1804) );
  OAI21_X1 U1903 ( .B1(n3674), .B2(n1803), .A(n1804), .ZN(n1805) );
  INV_X1 U1904 ( .A(\lt_x_134/B[4] ), .ZN(n1806) );
  OAI221_X1 U1905 ( .B1(\lt_x_134/B[4] ), .B2(n2829), .C1(n1806), .C2(n2828), 
        .A(n3006), .ZN(n1807) );
  OAI211_X1 U1906 ( .C1(n3700), .C2(n3390), .A(n3389), .B(n1807), .ZN(n1808)
         );
  AOI211_X1 U1907 ( .C1(n3007), .C2(n1800), .A(n1805), .B(n1808), .ZN(n350) );
  AOI22_X1 U1908 ( .A1(n3005), .A2(\DataP/alu_out_W[31] ), .B1(\DataP/B_s[31] ), .B2(n1859), .ZN(n1809) );
  AOI221_X1 U1909 ( .B1(n3709), .B2(n3983), .C1(n3984), .C2(n1799), .A(n3982), 
        .ZN(\DataP/right_br ) );
  AOI221_X1 U1910 ( .B1(n2061), .B2(n2103), .C1(n2102), .C2(n2103), .A(n2046), 
        .ZN(n1810) );
  INV_X1 U1911 ( .A(\DataP/alu_a_in[28] ), .ZN(n1811) );
  NAND2_X1 U1912 ( .A1(n3523), .A2(n1811), .ZN(n2515) );
  NAND2_X1 U1913 ( .A1(n2006), .A2(\DataP/alu_out_W[10] ), .ZN(n2388) );
  OR2_X1 U1914 ( .A1(\sra_131/SH[4] ), .A2(n3510), .ZN(n2461) );
  INV_X1 U1915 ( .A(n3470), .ZN(n1812) );
  NAND2_X1 U1916 ( .A1(n1929), .A2(n1812), .ZN(n3543) );
  INV_X1 U1917 ( .A(n3493), .ZN(n1813) );
  NAND2_X1 U1918 ( .A1(\DataP/alu_a_in[30] ), .A2(n1813), .ZN(n3683) );
  OR2_X1 U1919 ( .A1(n3401), .A2(\DataP/alu_a_in[14] ), .ZN(n3410) );
  AOI21_X1 U1920 ( .B1(n2543), .B2(n2547), .A(\DataP/alu_a_in[12] ), .ZN(n2542) );
  NAND2_X1 U1921 ( .A1(n3203), .A2(n3011), .ZN(n1814) );
  NAND2_X1 U1922 ( .A1(n1814), .A2(n3510), .ZN(n1815) );
  XNOR2_X1 U1923 ( .A(n1815), .B(n2330), .ZN(n3202) );
  NAND2_X1 U1924 ( .A1(n3358), .A2(n3361), .ZN(n1816) );
  NAND3_X1 U1925 ( .A1(n3007), .A2(n2602), .A3(n1806), .ZN(n3339) );
  OAI221_X1 U1926 ( .B1(n2981), .B2(n2924), .C1(n2981), .C2(n2065), .A(n3675), 
        .ZN(n3538) );
  AOI21_X1 U1927 ( .B1(n3466), .B2(n3467), .A(n3465), .ZN(n1817) );
  INV_X1 U1928 ( .A(n1817), .ZN(n2423) );
  AOI22_X1 U1929 ( .A1(n2127), .A2(n2670), .B1(n2846), .B2(n2626), .ZN(n1818)
         );
  MUX2_X1 U1930 ( .A(n1818), .B(n2692), .S(\lt_x_135/B[4] ), .Z(
        \DataP/ALU_C/shifter/N39 ) );
  AOI22_X1 U1931 ( .A1(n2064), .A2(n2653), .B1(n2846), .B2(n2611), .ZN(n1819)
         );
  MUX2_X1 U1932 ( .A(n1819), .B(n2673), .S(\lt_x_134/B[4] ), .Z(
        \DataP/ALU_C/shifter/N36 ) );
  INV_X1 U1933 ( .A(n3658), .ZN(n1820) );
  NAND2_X1 U1934 ( .A1(\DataP/alu_a_in[8] ), .A2(n1820), .ZN(n3657) );
  AOI22_X1 U1935 ( .A1(n2841), .A2(n2965), .B1(n2989), .B2(n2964), .ZN(n1821)
         );
  AOI22_X1 U1936 ( .A1(n1915), .A2(n2966), .B1(n2845), .B2(n1821), .ZN(n2967)
         );
  AOI22_X1 U1937 ( .A1(n2987), .A2(\DataP/alu_a_in[2] ), .B1(n2710), .B2(
        \DataP/alu_a_in[1] ), .ZN(n1822) );
  AOI22_X1 U1938 ( .A1(\sra_131/SH[1] ), .A2(n2942), .B1(n2988), .B2(n1822), 
        .ZN(n2905) );
  NOR3_X1 U1939 ( .A1(n3806), .A2(IR_CU[4]), .A3(IR_CU[5]), .ZN(n1823) );
  AOI21_X1 U1940 ( .B1(n3797), .B2(n606), .A(n1823), .ZN(n1824) );
  OAI221_X1 U1941 ( .B1(n3837), .B2(n3828), .C1(n3837), .C2(n3817), .A(n1824), 
        .ZN(n3807) );
  AOI22_X1 U1942 ( .A1(n2842), .A2(n2656), .B1(n1913), .B2(n2685), .ZN(n1825)
         );
  AOI22_X1 U1943 ( .A1(n2127), .A2(n1825), .B1(n2657), .B2(n1915), .ZN(n1826)
         );
  OAI221_X1 U1944 ( .B1(\lt_x_134/B[4] ), .B2(n1826), .C1(n1806), .C2(n2658), 
        .A(n3007), .ZN(n3480) );
  AND3_X1 U1945 ( .A1(n2475), .A2(n3070), .A3(n3064), .ZN(n3710) );
  NAND2_X1 U1946 ( .A1(n3765), .A2(n3766), .ZN(n1827) );
  NOR3_X1 U1947 ( .A1(n3770), .A2(n3771), .A3(n3772), .ZN(n1828) );
  NAND4_X1 U1948 ( .A1(n3773), .A2(n3774), .A3(n3769), .A4(n1828), .ZN(n1829)
         );
  NOR4_X1 U1949 ( .A1(n3767), .A2(n3768), .A3(n1827), .A4(n1829), .ZN(n1830)
         );
  INV_X1 U1950 ( .A(n3757), .ZN(n1831) );
  NAND4_X1 U1951 ( .A1(n3758), .A2(n3759), .A3(n3760), .A4(n1831), .ZN(n1832)
         );
  NOR2_X1 U1952 ( .A1(n3755), .A2(n3756), .ZN(n1833) );
  NAND3_X1 U1953 ( .A1(n3754), .A2(n3753), .A3(n1833), .ZN(n1834) );
  NOR4_X1 U1954 ( .A1(n3761), .A2(n3762), .A3(n1832), .A4(n1834), .ZN(n1835)
         );
  NAND4_X1 U1955 ( .A1(n3763), .A2(n3764), .A3(n1830), .A4(n1835), .ZN(n1836)
         );
  NAND2_X1 U1956 ( .A1(n3775), .A2(n1836), .ZN(\DataP/NPC_add/N0 ) );
  CLKBUF_X3 U1957 ( .A(n1907), .Z(n2988) );
  NAND4_X1 U1958 ( .A1(n2388), .A2(n3231), .A3(n3230), .A4(n2335), .ZN(n1879)
         );
  NOR2_X1 U1959 ( .A1(n3172), .A2(n3171), .ZN(n1838) );
  OR2_X2 U1960 ( .A1(n3131), .A2(n3130), .ZN(\DataP/alu_a_in[31] ) );
  AND2_X1 U1961 ( .A1(n3456), .A2(n3423), .ZN(n1840) );
  BUF_X2 U1962 ( .A(n3193), .Z(n2999) );
  INV_X1 U1963 ( .A(n1864), .ZN(n1841) );
  INV_X1 U1964 ( .A(\DataP/alu_a_in[15] ), .ZN(n1842) );
  INV_X1 U1965 ( .A(n1864), .ZN(\DataP/alu_a_in[15] ) );
  NOR2_X1 U1966 ( .A1(n3178), .A2(n3177), .ZN(n1864) );
  AND4_X1 U1967 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n1843)
         );
  BUF_X4 U1968 ( .A(\sra_131/SH[4] ), .Z(\lt_x_134/B[4] ) );
  NAND2_X1 U1969 ( .A1(n2469), .A2(n2470), .ZN(n1844) );
  NAND2_X1 U1970 ( .A1(n2469), .A2(n2470), .ZN(n1845) );
  NAND2_X1 U1971 ( .A1(n2469), .A2(n2470), .ZN(n2998) );
  OR2_X4 U1972 ( .A1(n3119), .A2(n3118), .ZN(\DataP/alu_a_in[4] ) );
  AND2_X1 U1973 ( .A1(n1518), .A2(\DataP/B_s[9] ), .ZN(n1846) );
  NAND4_X1 U1974 ( .A1(n1588), .A2(n2186), .A3(n3023), .A4(n2140), .ZN(n1847)
         );
  BUF_X1 U1975 ( .A(n3328), .Z(n1848) );
  BUF_X1 U1976 ( .A(n3328), .Z(n2565) );
  BUF_X1 U1977 ( .A(n3328), .Z(n1905) );
  AOI21_X2 U1978 ( .B1(n3412), .B2(n3411), .A(n2541), .ZN(n2540) );
  NAND3_X1 U1979 ( .A1(n1967), .A2(n3494), .A3(n3497), .ZN(n1849) );
  NAND3_X1 U1980 ( .A1(n3501), .A2(n3499), .A3(n3500), .ZN(n1850) );
  BUF_X1 U1981 ( .A(n3666), .Z(n1851) );
  INV_X1 U1982 ( .A(n1862), .ZN(n1852) );
  AND4_X2 U1983 ( .A1(n1853), .A2(n1854), .A3(n1855), .A4(n1856), .ZN(n2369)
         );
  AND3_X1 U1984 ( .A1(n3484), .A2(n3701), .A3(n3633), .ZN(n1854) );
  AND4_X1 U1985 ( .A1(n3615), .A2(n3624), .A3(n3651), .A4(n3390), .ZN(n1855)
         );
  AND2_X1 U1986 ( .A1(n3067), .A2(n3066), .ZN(n1857) );
  INV_X1 U1987 ( .A(n3001), .ZN(n1858) );
  INV_X1 U1988 ( .A(n1858), .ZN(n1859) );
  INV_X1 U1989 ( .A(n3396), .ZN(n1860) );
  AND3_X1 U1990 ( .A1(n2442), .A2(n1994), .A3(n2010), .ZN(n1889) );
  INV_X1 U1991 ( .A(n1565), .ZN(n3330) );
  BUF_X1 U1992 ( .A(n536), .Z(n1862) );
  NOR2_X2 U1993 ( .A1(n3190), .A2(n3189), .ZN(n1863) );
  AND3_X1 U1994 ( .A1(n3016), .A2(n3017), .A3(\DataP/opcode_W[3] ), .ZN(n1865)
         );
  AND2_X1 U1995 ( .A1(n2322), .A2(n2320), .ZN(n1866) );
  XOR2_X1 U1996 ( .A(n2570), .B(\DataP/add_D[3] ), .Z(n2186) );
  BUF_X1 U1997 ( .A(n1548), .Z(n1867) );
  OR2_X1 U1998 ( .A1(n1567), .A2(n117), .ZN(n1868) );
  INV_X1 U1999 ( .A(\DataP/dest_M[0] ), .ZN(n1869) );
  XNOR2_X1 U2000 ( .A(n2576), .B(n1894), .ZN(n3036) );
  XNOR2_X1 U2001 ( .A(n1870), .B(n1933), .ZN(n3446) );
  NOR2_X1 U2002 ( .A1(n3444), .A2(n3445), .ZN(n1870) );
  BUF_X1 U2003 ( .A(n538), .Z(n1871) );
  INV_X2 U2004 ( .A(n2126), .ZN(n2839) );
  INV_X2 U2005 ( .A(n1963), .ZN(n2845) );
  INV_X4 U2006 ( .A(n2845), .ZN(n1915) );
  INV_X1 U2007 ( .A(n1581), .ZN(n2064) );
  NOR2_X4 U2008 ( .A1(n3013), .A2(n4022), .ZN(n164) );
  INV_X1 U2009 ( .A(\DataP/add_S2[4] ), .ZN(n1872) );
  OR2_X2 U2012 ( .A1(n3167), .A2(n3166), .ZN(\DataP/alu_a_in[19] ) );
  AOI211_X2 U2013 ( .C1(n2108), .C2(n2107), .A(n2106), .B(n2105), .ZN(n2120)
         );
  NAND3_X1 U2014 ( .A1(n2449), .A2(n2448), .A3(n3270), .ZN(n1875) );
  OAI221_X1 U2015 ( .B1(n2122), .B2(n2121), .C1(n2122), .C2(n2120), .A(n2119), 
        .ZN(n1876) );
  INV_X2 U2016 ( .A(n1844), .ZN(n2995) );
  INV_X1 U2017 ( .A(n1893), .ZN(n1878) );
  NAND4_X1 U2018 ( .A1(n2388), .A2(n3231), .A3(n3230), .A4(n2335), .ZN(
        \DataP/alu_b_in[10] ) );
  BUF_X1 U2019 ( .A(n1581), .Z(n1963) );
  OR2_X1 U2020 ( .A1(\DataP/alu_b_in[13] ), .A2(\DataP/alu_b_in[12] ), .ZN(
        n1881) );
  NAND2_X1 U2021 ( .A1(n1875), .A2(n2225), .ZN(n1882) );
  BUF_X1 U2022 ( .A(n1847), .Z(n1883) );
  AND2_X1 U2023 ( .A1(n2576), .A2(n1543), .ZN(n3033) );
  INV_X1 U2024 ( .A(\DataP/alu_a_in[18] ), .ZN(n1884) );
  XNOR2_X1 U2025 ( .A(\DataP/add_D[0] ), .B(n1885), .ZN(n3025) );
  NAND3_X1 U2026 ( .A1(n2994), .A2(n2998), .A3(n2155), .ZN(n1887) );
  NAND3_X1 U2027 ( .A1(n1568), .A2(n2998), .A3(n2155), .ZN(n3193) );
  BUF_X1 U2028 ( .A(n3384), .Z(n1888) );
  MUX2_X2 U2029 ( .A(n3690), .B(n3701), .S(n3689), .Z(n3692) );
  NAND2_X1 U2030 ( .A1(n3545), .A2(n2552), .ZN(n1890) );
  INV_X1 U2031 ( .A(n1891), .ZN(n1892) );
  OR2_X2 U2032 ( .A1(n3076), .A2(n3075), .ZN(\DataP/alu_a_in[9] ) );
  AND2_X1 U2033 ( .A1(n1978), .A2(n1979), .ZN(n1893) );
  NOR3_X1 U2034 ( .A1(n1582), .A2(n2389), .A3(n2333), .ZN(n1896) );
  NOR3_X1 U2035 ( .A1(n1582), .A2(n2389), .A3(n2333), .ZN(n1897) );
  NOR3_X1 U2036 ( .A1(n1582), .A2(n2389), .A3(n2333), .ZN(n3263) );
  OR2_X2 U2037 ( .A1(n3079), .A2(n3078), .ZN(\DataP/alu_a_in[7] ) );
  NOR2_X1 U2038 ( .A1(n1572), .A2(\DataP/alu_b_in[10] ), .ZN(n1898) );
  BUF_X1 U2039 ( .A(n3381), .Z(n1899) );
  AND4_X1 U2040 ( .A1(n1564), .A2(n2498), .A3(n3086), .A4(n3085), .ZN(n1900)
         );
  AND2_X1 U2041 ( .A1(n1879), .A2(n2083), .ZN(n1901) );
  AND2_X1 U2042 ( .A1(n1572), .A2(n1863), .ZN(n1902) );
  NOR2_X1 U2043 ( .A1(n1901), .A2(n1902), .ZN(n2088) );
  NOR2_X1 U2044 ( .A1(n1966), .A2(n1910), .ZN(n1903) );
  AOI21_X1 U2045 ( .B1(n3039), .B2(n3038), .A(n2157), .ZN(n1904) );
  NOR2_X1 U2046 ( .A1(n1966), .A2(n1910), .ZN(n2010) );
  NAND2_X1 U2047 ( .A1(n3503), .A2(n3502), .ZN(n1906) );
  AOI21_X1 U2048 ( .B1(n1890), .B2(n2224), .A(n2427), .ZN(n1908) );
  OR2_X1 U2049 ( .A1(n3685), .A2(n3684), .ZN(n1909) );
  OR2_X1 U2050 ( .A1(n3685), .A2(n3684), .ZN(n3708) );
  NAND4_X2 U2051 ( .A1(n3098), .A2(n3099), .A3(n3096), .A4(n3097), .ZN(n1910)
         );
  CLKBUF_X3 U2052 ( .A(n3327), .Z(n3001) );
  AND4_X2 U2053 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n2130)
         );
  AND2_X1 U2054 ( .A1(n1635), .A2(\DataP/B_s[6] ), .ZN(n1911) );
  OR2_X2 U2055 ( .A1(\DataP/alu_b_in[17] ), .A2(n3510), .ZN(n2538) );
  INV_X2 U2056 ( .A(n1580), .ZN(\DataP/alu_b_in[17] ) );
  OR2_X2 U2057 ( .A1(n3170), .A2(n3169), .ZN(\DataP/alu_a_in[18] ) );
  NOR2_X2 U2058 ( .A1(n1562), .A2(n3116), .ZN(n1996) );
  NAND4_X1 U2059 ( .A1(n3098), .A2(n3099), .A3(n3096), .A4(n3097), .ZN(
        \DataP/alu_b_in[2] ) );
  INV_X1 U2060 ( .A(\DataP/alu_a_in[27] ), .ZN(n1912) );
  OR2_X1 U2061 ( .A1(n3137), .A2(n3136), .ZN(\DataP/alu_a_in[29] ) );
  OR2_X1 U2062 ( .A1(n3161), .A2(n3160), .ZN(\DataP/alu_a_in[21] ) );
  OR2_X1 U2063 ( .A1(n2302), .A2(n2145), .ZN(\DataP/alu_b_in[18] ) );
  OR2_X1 U2064 ( .A1(n3134), .A2(n3133), .ZN(\DataP/alu_a_in[30] ) );
  OR2_X1 U2065 ( .A1(n3128), .A2(n3127), .ZN(\DataP/alu_a_in[8] ) );
  INV_X1 U2066 ( .A(n2843), .ZN(n1930) );
  BUF_X2 U2067 ( .A(n2990), .Z(n2842) );
  INV_X2 U2068 ( .A(n2714), .ZN(n1913) );
  INV_X2 U2069 ( .A(n2838), .ZN(n1914) );
  BUF_X4 U2070 ( .A(n1907), .Z(n1916) );
  INV_X1 U2071 ( .A(\DataP/alu_b_in[28] ), .ZN(n1917) );
  INV_X1 U2072 ( .A(n3510), .ZN(n1918) );
  INV_X1 U2073 ( .A(n3911), .ZN(n1919) );
  INV_X1 U2074 ( .A(\DataP/alu_a_in[5] ), .ZN(n1920) );
  INV_X1 U2075 ( .A(\DataP/alu_a_in[8] ), .ZN(n1921) );
  INV_X1 U2076 ( .A(\DataP/alu_a_in[9] ), .ZN(n1922) );
  INV_X1 U2077 ( .A(\DataP/alu_a_in[31] ), .ZN(n1923) );
  INV_X1 U2078 ( .A(\DataP/alu_a_in[30] ), .ZN(n1924) );
  INV_X1 U2079 ( .A(\DataP/alu_a_in[29] ), .ZN(n1925) );
  INV_X1 U2080 ( .A(\DataP/alu_a_in[7] ), .ZN(n1926) );
  INV_X1 U2081 ( .A(\DataP/alu_a_in[13] ), .ZN(n1927) );
  INV_X1 U2082 ( .A(\DataP/alu_b_in[18] ), .ZN(n1928) );
  INV_X1 U2083 ( .A(\DataP/alu_a_in[25] ), .ZN(n1929) );
  BUF_X2 U2084 ( .A(n2990), .Z(n2841) );
  BUF_X2 U2085 ( .A(n2838), .Z(n1931) );
  INV_X1 U2086 ( .A(\DataP/alu_b_in[22] ), .ZN(n1933) );
  INV_X1 U2087 ( .A(\DataP/alu_b_in[29] ), .ZN(n1934) );
  INV_X1 U2088 ( .A(\DataP/alu_b_in[31] ), .ZN(n1935) );
  INV_X1 U2089 ( .A(\DataP/alu_b_in[26] ), .ZN(n1936) );
  INV_X1 U2090 ( .A(\DataP/alu_b_in[23] ), .ZN(n1937) );
  INV_X1 U2091 ( .A(n3510), .ZN(n1938) );
  INV_X1 U2092 ( .A(n3700), .ZN(n1939) );
  AOI21_X1 U2093 ( .B1(n3522), .B2(n1919), .A(n1981), .ZN(n1980) );
  NOR2_X1 U2094 ( .A1(n3910), .A2(n4019), .ZN(n1981) );
  AND4_X1 U2095 ( .A1(n2395), .A2(n2393), .A3(n2396), .A4(n2392), .ZN(n301) );
  AND4_X1 U2096 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n2137)
         );
  INV_X2 U2097 ( .A(n3010), .ZN(n1940) );
  OAI21_X1 U2098 ( .B1(n3248), .B2(n1976), .A(n1985), .ZN(n3252) );
  OR2_X1 U2099 ( .A1(n3515), .A2(n3514), .ZN(n2243) );
  NOR2_X1 U2100 ( .A1(n3234), .A2(n1976), .ZN(n3235) );
  AND2_X1 U2101 ( .A1(n3416), .A2(n3415), .ZN(n3456) );
  XNOR2_X1 U2102 ( .A(n3213), .B(\DataP/alu_a_in[7] ), .ZN(n3387) );
  AND2_X1 U2103 ( .A1(n3393), .A2(n3416), .ZN(n3413) );
  AND2_X1 U2104 ( .A1(n2282), .A2(n2283), .ZN(n1958) );
  AND2_X1 U2105 ( .A1(\DataP/alu_a_in[10] ), .A2(n2357), .ZN(n2356) );
  INV_X1 U2106 ( .A(\DataP/alu_a_in[12] ), .ZN(n1941) );
  INV_X1 U2107 ( .A(\DataP/alu_a_in[3] ), .ZN(n1942) );
  OR2_X1 U2108 ( .A1(n3196), .A2(n3195), .ZN(\DataP/alu_a_in[10] ) );
  INV_X1 U2109 ( .A(\DataP/alu_a_in[23] ), .ZN(n1943) );
  OR2_X1 U2110 ( .A1(n3158), .A2(n3157), .ZN(\DataP/alu_a_in[22] ) );
  OR2_X1 U2111 ( .A1(n3175), .A2(n3174), .ZN(\DataP/alu_a_in[16] ) );
  INV_X1 U2112 ( .A(\DataP/alu_a_in[20] ), .ZN(n1944) );
  OR2_X1 U2113 ( .A1(n3152), .A2(n3151), .ZN(\DataP/alu_a_in[24] ) );
  OR2_X1 U2114 ( .A1(n3146), .A2(n3145), .ZN(\DataP/alu_a_in[26] ) );
  INV_X1 U2115 ( .A(\DataP/alu_a_in[19] ), .ZN(n1945) );
  OR2_X1 U2116 ( .A1(n3140), .A2(n3139), .ZN(\DataP/alu_a_in[28] ) );
  INV_X2 U2117 ( .A(n1448), .ZN(n4022) );
  INV_X1 U2118 ( .A(\DataP/alu_b_in[19] ), .ZN(n1946) );
  AND2_X1 U2119 ( .A1(n3473), .A2(n1550), .ZN(n2241) );
  INV_X1 U2120 ( .A(n2985), .ZN(n2987) );
  INV_X1 U2121 ( .A(n1916), .ZN(\sra_131/SH[1] ) );
  BUF_X1 U2122 ( .A(n2990), .Z(n2714) );
  INV_X1 U2123 ( .A(n1932), .ZN(n1947) );
  BUF_X1 U2124 ( .A(n2990), .Z(n2843) );
  INV_X2 U2125 ( .A(n2847), .ZN(\lt_x_135/B[4] ) );
  INV_X1 U2126 ( .A(\DataP/alu_b_in[5] ), .ZN(n1948) );
  INV_X1 U2127 ( .A(\DataP/alu_b_in[21] ), .ZN(n3442) );
  INV_X1 U2128 ( .A(\DataP/alu_b_in[15] ), .ZN(n1949) );
  INV_X1 U2129 ( .A(\DataP/alu_b_in[7] ), .ZN(n1950) );
  INV_X1 U2130 ( .A(\DataP/alu_b_in[16] ), .ZN(n1951) );
  INV_X2 U2131 ( .A(n2004), .ZN(n2985) );
  INV_X1 U2132 ( .A(\DataP/alu_b_in[21] ), .ZN(n1952) );
  NAND2_X1 U2133 ( .A1(n2006), .A2(\DataP/alu_out_W[6] ), .ZN(n2152) );
  INV_X1 U2134 ( .A(n3071), .ZN(n2469) );
  NOR2_X1 U2135 ( .A1(n3674), .A2(n3911), .ZN(n1982) );
  OAI21_X1 U2136 ( .B1(n3948), .B2(n3947), .A(Rst), .ZN(n3949) );
  INV_X1 U2137 ( .A(n3065), .ZN(n2471) );
  NAND2_X2 U2138 ( .A1(n3229), .A2(Rst), .ZN(n3910) );
  OR2_X2 U2139 ( .A1(n3008), .A2(n3943), .ZN(n3946) );
  INV_X1 U2140 ( .A(n3856), .ZN(n3837) );
  AND2_X2 U2141 ( .A1(\WB_MUX_SEL_i[1] ), .A2(n294), .ZN(n3943) );
  CLKBUF_X1 U2142 ( .A(\DataP/add_D[2] ), .Z(n1955) );
  NOR2_X1 U2143 ( .A1(IR_CU_27), .A2(IR_CU_26), .ZN(n3856) );
  AOI21_X1 U2144 ( .B1(n2413), .B2(n3691), .A(n2226), .ZN(n2567) );
  AND3_X1 U2145 ( .A1(n3692), .A2(n3705), .A3(n3691), .ZN(n2153) );
  NOR2_X2 U2146 ( .A1(n3345), .A2(n3903), .ZN(n3703) );
  BUF_X2 U2147 ( .A(n3706), .Z(n3007) );
  NAND2_X2 U2148 ( .A1(n3223), .A2(n3226), .ZN(n3700) );
  NAND3_X1 U2149 ( .A1(n1606), .A2(n3494), .A3(n3497), .ZN(n3501) );
  OAI21_X1 U2150 ( .B1(\DataP/opcode_W[2] ), .B2(\DataP/opcode_W[1] ), .A(
        \DataP/opcode_W[4] ), .ZN(n1953) );
  AND2_X2 U2151 ( .A1(n1563), .A2(n2136), .ZN(n2503) );
  BUF_X1 U2152 ( .A(n3377), .Z(n1954) );
  NAND3_X1 U2153 ( .A1(n2449), .A2(n2448), .A3(n3270), .ZN(n2290) );
  OAI21_X1 U2154 ( .B1(n1957), .B2(n1918), .A(n2366), .ZN(n2419) );
  INV_X1 U2155 ( .A(n1607), .ZN(n2420) );
  NAND3_X1 U2156 ( .A1(n3408), .A2(n2284), .A3(n1958), .ZN(n3647) );
  NAND2_X1 U2157 ( .A1(n3233), .A2(n3510), .ZN(n1977) );
  NAND2_X1 U2158 ( .A1(n1977), .A2(n2356), .ZN(n2450) );
  BUF_X1 U2159 ( .A(n1557), .Z(n1960) );
  BUF_X1 U2160 ( .A(n3669), .Z(n1961) );
  NAND2_X1 U2161 ( .A1(n3411), .A2(n3409), .ZN(n1962) );
  NOR2_X1 U2162 ( .A1(\DataP/alu_b_in[13] ), .A2(\DataP/alu_b_in[12] ), .ZN(
        n3419) );
  NAND2_X1 U2163 ( .A1(n1964), .A2(n3510), .ZN(n2339) );
  XNOR2_X1 U2164 ( .A(n2009), .B(\DataP/alu_b_in[0] ), .ZN(n1964) );
  NAND4_X1 U2165 ( .A1(n3090), .A2(n3089), .A3(n3091), .A4(n3088), .ZN(
        \DataP/alu_b_in[0] ) );
  NAND4_X1 U2166 ( .A1(n1564), .A2(n2498), .A3(n3086), .A4(n3085), .ZN(n2506)
         );
  AND3_X2 U2167 ( .A1(n1524), .A2(n1900), .A3(n2362), .ZN(n2442) );
  NAND3_X1 U2168 ( .A1(n2500), .A2(n2499), .A3(n2152), .ZN(n1965) );
  NAND2_X1 U2169 ( .A1(n1637), .A2(n3214), .ZN(n1966) );
  NAND2_X1 U2170 ( .A1(n2002), .A2(n3494), .ZN(n3467) );
  NAND2_X1 U2171 ( .A1(n2425), .A2(n2540), .ZN(n1967) );
  XNOR2_X1 U2172 ( .A(n3202), .B(\DataP/alu_a_in[3] ), .ZN(n3678) );
  INV_X1 U2173 ( .A(n1968), .ZN(n300) );
  OAI211_X1 U2174 ( .C1(n1975), .C2(n2008), .A(n1972), .B(n1969), .ZN(n1968)
         );
  INV_X1 U2175 ( .A(n1970), .ZN(n1969) );
  OAI21_X1 U2176 ( .B1(n1975), .B2(n2550), .A(n1971), .ZN(n1970) );
  INV_X1 U2177 ( .A(n3531), .ZN(n1971) );
  NAND2_X1 U2178 ( .A1(n2008), .A2(n1973), .ZN(n1972) );
  AND2_X1 U2179 ( .A1(n2550), .A2(n1974), .ZN(n1973) );
  NOR2_X1 U2180 ( .A1(n3524), .A2(n3674), .ZN(n1974) );
  NAND2_X1 U2181 ( .A1(n3524), .A2(n3691), .ZN(n1975) );
  NAND2_X1 U2182 ( .A1(n1906), .A2(n2552), .ZN(n2008) );
  NAND2_X1 U2183 ( .A1(n1978), .A2(n1979), .ZN(n3458) );
  NAND2_X1 U2184 ( .A1(n3422), .A2(n2512), .ZN(n1978) );
  AOI21_X1 U2185 ( .B1(n2418), .B2(n3691), .A(n3522), .ZN(n299) );
  OAI221_X1 U2186 ( .B1(n2059), .B2(n2058), .C1(n2059), .C2(n2057), .A(n2056), 
        .ZN(n1983) );
  AOI21_X1 U2187 ( .B1(n3354), .B2(n2438), .A(n2437), .ZN(n1984) );
  AND2_X1 U2188 ( .A1(n3488), .A2(n3509), .ZN(n3490) );
  BUF_X1 U2189 ( .A(n3268), .Z(n1985) );
  NAND2_X1 U2190 ( .A1(n2002), .A2(n3456), .ZN(n1986) );
  AOI21_X1 U2191 ( .B1(n2131), .B2(n3465), .A(n2421), .ZN(n1988) );
  NAND2_X1 U2192 ( .A1(n2424), .A2(n2523), .ZN(n1989) );
  INV_X1 U2193 ( .A(n2535), .ZN(n1990) );
  BUF_X1 U2194 ( .A(n1909), .Z(n1991) );
  XNOR2_X1 U2195 ( .A(n2293), .B(n2292), .ZN(n1992) );
  BUF_X1 U2196 ( .A(n3677), .Z(n1993) );
  AND2_X1 U2197 ( .A1(n1569), .A2(n2130), .ZN(n1995) );
  AND2_X1 U2198 ( .A1(n3088), .A2(n3084), .ZN(n2498) );
  AND3_X1 U2199 ( .A1(n2449), .A2(n3270), .A3(n2448), .ZN(n1997) );
  AND3_X2 U2200 ( .A1(n3329), .A2(n1565), .A3(n2189), .ZN(n2564) );
  OAI211_X1 U2201 ( .C1(n3441), .C2(n1531), .A(n1559), .B(n1960), .ZN(n1998)
         );
  INV_X1 U2202 ( .A(\DataP/dest_M[2] ), .ZN(n1999) );
  OAI211_X1 U2203 ( .C1(n2492), .C2(n2494), .A(n2489), .B(n2491), .ZN(n2000)
         );
  BUF_X1 U2204 ( .A(n1587), .Z(n2001) );
  NAND2_X1 U2205 ( .A1(n1882), .A2(n2540), .ZN(n2002) );
  NAND2_X1 U2206 ( .A1(n1577), .A2(n1608), .ZN(n2003) );
  NAND2_X1 U2207 ( .A1(n1577), .A2(n1608), .ZN(n3216) );
  NAND4_X1 U2208 ( .A1(n1542), .A2(n1564), .A3(n3089), .A4(n3088), .ZN(n2004)
         );
  INV_X1 U2209 ( .A(n1565), .ZN(n2006) );
  OAI21_X1 U2210 ( .B1(n2365), .B2(n2321), .A(n2364), .ZN(n2007) );
  NAND2_X2 U2211 ( .A1(n1845), .A2(n2143), .ZN(n2561) );
  INV_X1 U2212 ( .A(n2843), .ZN(n2844) );
  NAND4_X1 U2213 ( .A1(n3087), .A2(n3085), .A3(n3086), .A4(n3084), .ZN(n2009)
         );
  OAI21_X1 U2214 ( .B1(n2380), .B2(n2577), .A(n2379), .ZN(n2011) );
  OAI21_X1 U2215 ( .B1(n2577), .B2(n2380), .A(n2379), .ZN(n3577) );
  OAI211_X1 U2216 ( .C1(n3212), .C2(n1517), .A(n3211), .B(n3387), .ZN(n2012)
         );
  OR2_X2 U2217 ( .A1(n3113), .A2(n3114), .ZN(\DataP/alu_a_in[0] ) );
  OAI21_X1 U2218 ( .B1(\DataP/alu_b_in[30] ), .B2(n1924), .A(n2013), .ZN(n2048) );
  AOI211_X1 U2219 ( .C1(\DataP/alu_a_in[28] ), .C2(n1917), .A(n2067), .B(n2048), .ZN(n2050) );
  AOI211_X1 U2220 ( .C1(\DataP/alu_a_in[24] ), .C2(n1550), .A(n2113), .B(n2060), .ZN(n2014) );
  NAND2_X1 U2221 ( .A1(n1573), .A2(n2014), .ZN(n2059) );
  NOR2_X1 U2222 ( .A1(\DataP/alu_b_in[9] ), .A2(n1922), .ZN(n2029) );
  NAND2_X1 U2223 ( .A1(\DataP/alu_a_in[13] ), .A2(n3396), .ZN(n2015) );
  OAI211_X1 U2224 ( .C1(n1880), .C2(n1941), .A(n2035), .B(n2015), .ZN(n2031)
         );
  NOR2_X1 U2225 ( .A1(\DataP/alu_b_in[8] ), .A2(n1921), .ZN(n2017) );
  AOI21_X1 U2226 ( .B1(n2358), .B2(\DataP/alu_a_in[10] ), .A(n2028), .ZN(n2016) );
  OR4_X1 U2227 ( .A1(n2029), .A2(n2031), .A3(n2017), .A4(n2063), .ZN(n2038) );
  OAI21_X1 U2228 ( .B1(\lt_x_134/B[5] ), .B2(n1920), .A(\lt_x_134/B[4] ), .ZN(
        n2018) );
  OAI22_X1 U2229 ( .A1(\DataP/alu_a_in[4] ), .A2(n2018), .B1(
        \DataP/alu_a_in[5] ), .B2(n1948), .ZN(n2026) );
  AOI21_X1 U2230 ( .B1(\DataP/alu_a_in[6] ), .B2(n1611), .A(n2072), .ZN(n2025)
         );
  OAI21_X1 U2231 ( .B1(n1612), .B2(n1996), .A(n1537), .ZN(n2019) );
  OAI22_X1 U2232 ( .A1(n1605), .A2(n2019), .B1(\DataP/alu_a_in[1] ), .B2(n2126), .ZN(n2020) );
  OAI221_X1 U2233 ( .B1(n1963), .B2(n1942), .C1(n1910), .C2(n1561), .A(n2020), 
        .ZN(n2021) );
  OAI221_X1 U2234 ( .B1(\DataP/alu_a_in[3] ), .B2(n2064), .C1(
        \DataP/alu_a_in[2] ), .C2(n2076), .A(n2021), .ZN(n2022) );
  OAI21_X1 U2235 ( .B1(\lt_x_134/B[5] ), .B2(n1920), .A(n2022), .ZN(n2023) );
  AOI221_X1 U2236 ( .B1(n2026), .B2(n2025), .C1(n2024), .C2(n2025), .A(n2080), 
        .ZN(n2037) );
  OAI21_X1 U2237 ( .B1(n1860), .B2(n1927), .A(n1880), .ZN(n2027) );
  AOI22_X1 U2238 ( .A1(n2083), .A2(n1879), .B1(n1572), .B2(n1863), .ZN(n2033)
         );
  NOR2_X1 U2239 ( .A1(\DataP/alu_a_in[8] ), .A2(n2029), .ZN(n2030) );
  AOI22_X1 U2240 ( .A1(n2030), .A2(\DataP/alu_b_in[8] ), .B1(
        \DataP/alu_b_in[9] ), .B2(n1922), .ZN(n2032) );
  AOI221_X1 U2241 ( .B1(n2063), .B2(n2033), .C1(n2032), .C2(n2033), .A(n2031), 
        .ZN(n2034) );
  AOI211_X1 U2242 ( .C1(n2035), .C2(n2092), .A(n2090), .B(n2034), .ZN(n2036)
         );
  OAI21_X1 U2243 ( .B1(n2037), .B2(n2038), .A(n2036), .ZN(n2042) );
  NOR2_X1 U2244 ( .A1(\DataP/alu_b_in[23] ), .A2(n1943), .ZN(n2039) );
  AOI21_X1 U2245 ( .B1(\DataP/alu_a_in[22] ), .B2(n1933), .A(n2039), .ZN(n2047) );
  NAND2_X1 U2246 ( .A1(\DataP/alu_a_in[21] ), .A2(n1952), .ZN(n2040) );
  OAI211_X1 U2247 ( .C1(\DataP/alu_b_in[20] ), .C2(n1944), .A(n2047), .B(n2040), .ZN(n2046) );
  NOR2_X1 U2248 ( .A1(\DataP/alu_b_in[19] ), .A2(n1945), .ZN(n2043) );
  AOI211_X1 U2249 ( .C1(\DataP/alu_a_in[16] ), .C2(n1951), .A(n2046), .B(n2061), .ZN(n2041) );
  NAND3_X1 U2250 ( .A1(n2042), .A2(n2125), .A3(n2041), .ZN(n2058) );
  NOR2_X1 U2251 ( .A1(\DataP/alu_a_in[18] ), .A2(n2043), .ZN(n2044) );
  NOR2_X1 U2252 ( .A1(\DataP/alu_a_in[16] ), .A2(n2100), .ZN(n2045) );
  OAI22_X1 U2253 ( .A1(\DataP/alu_a_in[28] ), .A2(n2110), .B1(
        \DataP/alu_a_in[29] ), .B2(n1934), .ZN(n2055) );
  AOI22_X1 U2254 ( .A1(\DataP/alu_b_in[26] ), .A2(n2112), .B1(
        \DataP/alu_b_in[27] ), .B2(n1912), .ZN(n2052) );
  NOR2_X1 U2255 ( .A1(\DataP/alu_a_in[24] ), .A2(n2113), .ZN(n2049) );
  AOI22_X1 U2256 ( .A1(\DataP/alu_b_in[24] ), .A2(n2049), .B1(
        \DataP/alu_b_in[25] ), .B2(n1929), .ZN(n2051) );
  AOI221_X1 U2257 ( .B1(n2060), .B2(n2052), .C1(n2051), .C2(n2052), .A(n2062), 
        .ZN(n2054) );
  OAI21_X1 U2258 ( .B1(\DataP/alu_a_in[31] ), .B2(n1935), .A(
        \DataP/alu_b_in[30] ), .ZN(n2053) );
  OAI221_X1 U2259 ( .B1(n2059), .B2(n2058), .C1(n2059), .C2(n2057), .A(n2056), 
        .ZN(\DataP/ALU_C/comp/N24 ) );
  INV_X1 U2260 ( .A(\lt_x_134/B[4] ), .ZN(n2065) );
  AOI22_X1 U2261 ( .A1(\DataP/alu_a_in[15] ), .A2(n1949), .B1(
        \DataP/alu_a_in[14] ), .B2(n1947), .ZN(n2035) );
  INV_X1 U2262 ( .A(n2016), .ZN(n2063) );
  INV_X1 U2263 ( .A(n2097), .ZN(n2061) );
  INV_X1 U2264 ( .A(n2050), .ZN(n2062) );
  NOR2_X1 U2265 ( .A1(\DataP/alu_b_in[29] ), .A2(n1925), .ZN(n2067) );
  NAND2_X1 U2266 ( .A1(\DataP/alu_a_in[31] ), .A2(n1935), .ZN(n2066) );
  OAI21_X1 U2267 ( .B1(\DataP/alu_b_in[30] ), .B2(n1924), .A(n2066), .ZN(n2109) );
  AOI211_X1 U2268 ( .C1(\DataP/alu_a_in[28] ), .C2(n1917), .A(n2067), .B(n2109), .ZN(n2115) );
  NOR2_X1 U2269 ( .A1(\DataP/alu_b_in[25] ), .A2(n1929), .ZN(n2113) );
  NOR2_X1 U2270 ( .A1(n1912), .A2(\DataP/alu_b_in[27] ), .ZN(n2111) );
  AOI21_X1 U2271 ( .B1(n1936), .B2(\DataP/alu_a_in[26] ), .A(n2111), .ZN(n2068) );
  AOI211_X1 U2272 ( .C1(\DataP/alu_a_in[24] ), .C2(n1550), .A(n2113), .B(n2123), .ZN(n2069) );
  NAND2_X1 U2273 ( .A1(n2115), .A2(n2069), .ZN(n2122) );
  NOR2_X1 U2274 ( .A1(\DataP/alu_b_in[9] ), .A2(n1922), .ZN(n2084) );
  NOR2_X1 U2275 ( .A1(\DataP/alu_b_in[15] ), .A2(n1864), .ZN(n2070) );
  AOI21_X1 U2276 ( .B1(\DataP/alu_a_in[14] ), .B2(n1947), .A(n2070), .ZN(n2093) );
  OAI211_X1 U2277 ( .C1(n1880), .C2(n1941), .A(n2093), .B(n2015), .ZN(n2086)
         );
  OR4_X1 U2278 ( .A1(n2084), .A2(n2086), .A3(n2017), .A4(n2063), .ZN(n2096) );
  OAI21_X1 U2279 ( .B1(\lt_x_134/B[5] ), .B2(n1920), .A(\lt_x_134/B[4] ), .ZN(
        n2071) );
  OAI22_X1 U2280 ( .A1(\DataP/alu_a_in[4] ), .A2(n2071), .B1(
        \DataP/alu_a_in[5] ), .B2(n1948), .ZN(n2082) );
  NOR2_X1 U2281 ( .A1(\DataP/alu_b_in[7] ), .A2(n1926), .ZN(n2072) );
  OAI21_X1 U2282 ( .B1(n1963), .B2(n1942), .A(n1910), .ZN(n2076) );
  OAI21_X1 U2283 ( .B1(n1612), .B2(n1996), .A(n2004), .ZN(n2073) );
  OAI22_X1 U2284 ( .A1(n1605), .A2(n2073), .B1(\DataP/alu_a_in[1] ), .B2(n2126), .ZN(n2074) );
  OAI221_X1 U2285 ( .B1(n1963), .B2(n1942), .C1(n1910), .C2(n1561), .A(n2074), 
        .ZN(n2075) );
  OAI221_X1 U2286 ( .B1(\DataP/alu_a_in[3] ), .B2(n2127), .C1(
        \DataP/alu_a_in[2] ), .C2(n2076), .A(n2075), .ZN(n2077) );
  OAI21_X1 U2287 ( .B1(\lt_x_134/B[5] ), .B2(n1920), .A(n2077), .ZN(n2078) );
  AOI21_X1 U2288 ( .B1(\DataP/alu_a_in[4] ), .B2(n2847), .A(n2078), .ZN(n2081)
         );
  OAI21_X1 U2289 ( .B1(\DataP/alu_b_in[7] ), .B2(n1926), .A(
        \DataP/alu_b_in[6] ), .ZN(n2079) );
  OAI22_X1 U2290 ( .A1(\DataP/alu_a_in[6] ), .A2(n2079), .B1(
        \DataP/alu_a_in[7] ), .B2(n1950), .ZN(n2080) );
  AOI221_X1 U2291 ( .B1(n2082), .B2(n2025), .C1(n2081), .C2(n2025), .A(n2080), 
        .ZN(n2095) );
  OAI22_X1 U2292 ( .A1(\DataP/alu_a_in[12] ), .A2(n2027), .B1(
        \DataP/alu_a_in[13] ), .B2(n3396), .ZN(n2092) );
  NOR2_X1 U2293 ( .A1(\DataP/alu_a_in[10] ), .A2(n2028), .ZN(n2083) );
  NOR2_X1 U2294 ( .A1(\DataP/alu_a_in[8] ), .A2(n2084), .ZN(n2085) );
  AOI22_X1 U2295 ( .A1(\DataP/alu_b_in[8] ), .A2(n2085), .B1(
        \DataP/alu_b_in[9] ), .B2(n1922), .ZN(n2087) );
  AOI221_X1 U2296 ( .B1(n2063), .B2(n2088), .C1(n2087), .C2(n2088), .A(n2086), 
        .ZN(n2091) );
  OAI21_X1 U2297 ( .B1(\DataP/alu_b_in[15] ), .B2(n1842), .A(n1932), .ZN(n2089) );
  OAI22_X1 U2298 ( .A1(\DataP/alu_a_in[14] ), .A2(n2089), .B1(n1841), .B2(
        n1949), .ZN(n2090) );
  AOI211_X1 U2299 ( .C1(n2093), .C2(n2092), .A(n2090), .B(n2091), .ZN(n2094)
         );
  OAI21_X1 U2300 ( .B1(n2096), .B2(n2095), .A(n2094), .ZN(n2099) );
  NOR2_X1 U2301 ( .A1(\DataP/alu_b_in[17] ), .A2(n1838), .ZN(n2100) );
  AOI21_X1 U2302 ( .B1(\DataP/alu_a_in[22] ), .B2(n1933), .A(n2039), .ZN(n2108) );
  OAI211_X1 U2303 ( .C1(\DataP/alu_b_in[20] ), .C2(n1944), .A(n2108), .B(n2040), .ZN(n2101) );
  AOI21_X1 U2304 ( .B1(n1928), .B2(\DataP/alu_a_in[18] ), .A(n2043), .ZN(n2097) );
  AOI211_X1 U2305 ( .C1(\DataP/alu_a_in[16] ), .C2(n1951), .A(n2101), .B(n2061), .ZN(n2098) );
  NAND3_X1 U2306 ( .A1(n2099), .A2(n2125), .A3(n2098), .ZN(n2121) );
  AOI22_X1 U2307 ( .A1(\DataP/alu_b_in[18] ), .A2(n2044), .B1(
        \DataP/alu_b_in[19] ), .B2(n1945), .ZN(n2103) );
  AOI22_X1 U2308 ( .A1(\DataP/alu_b_in[16] ), .A2(n2045), .B1(
        \DataP/alu_b_in[17] ), .B2(n1838), .ZN(n2102) );
  AOI221_X1 U2309 ( .B1(n2061), .B2(n2103), .C1(n2102), .C2(n2103), .A(n2101), 
        .ZN(n2106) );
  OAI21_X1 U2310 ( .B1(\DataP/alu_b_in[23] ), .B2(n1943), .A(
        \DataP/alu_b_in[22] ), .ZN(n2104) );
  OAI22_X1 U2311 ( .A1(\DataP/alu_a_in[22] ), .A2(n2104), .B1(
        \DataP/alu_a_in[23] ), .B2(n1937), .ZN(n2105) );
  OAI21_X1 U2312 ( .B1(\DataP/alu_b_in[29] ), .B2(n1925), .A(
        \DataP/alu_b_in[28] ), .ZN(n2110) );
  NOR2_X1 U2313 ( .A1(\DataP/alu_a_in[26] ), .A2(n2111), .ZN(n2112) );
  AOI22_X1 U2314 ( .A1(\DataP/alu_b_in[26] ), .A2(n2112), .B1(
        \DataP/alu_b_in[27] ), .B2(n1912), .ZN(n2117) );
  NOR2_X1 U2315 ( .A1(\DataP/alu_a_in[24] ), .A2(n2113), .ZN(n2114) );
  AOI22_X1 U2316 ( .A1(\DataP/alu_b_in[24] ), .A2(n2114), .B1(
        \DataP/alu_b_in[25] ), .B2(n1929), .ZN(n2116) );
  OAI21_X1 U2317 ( .B1(\DataP/alu_b_in[31] ), .B2(n1923), .A(
        \DataP/alu_b_in[30] ), .ZN(n2118) );
  INV_X1 U2318 ( .A(n1612), .ZN(n2126) );
  INV_X1 U2319 ( .A(\DataP/alu_b_in[3] ), .ZN(n2127) );
  INV_X1 U2320 ( .A(n2068), .ZN(n2123) );
  INV_X1 U2321 ( .A(n2100), .ZN(n2125) );
  INV_X1 U2322 ( .A(n2115), .ZN(n2124) );
  NAND2_X1 U2323 ( .A1(n1566), .A2(n2313), .ZN(n3329) );
  AND2_X1 U2324 ( .A1(n3021), .A2(n3022), .ZN(n2480) );
  NAND4_X1 U2325 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(
        \DataP/alu_b_in[5] ) );
  OR2_X1 U2326 ( .A1(n2231), .A2(n3003), .ZN(n3093) );
  OR2_X1 U2327 ( .A1(n3003), .A2(n2227), .ZN(n3105) );
  INV_X1 U2328 ( .A(n1844), .ZN(n2996) );
  OR2_X1 U2329 ( .A1(n3070), .A2(n3012), .ZN(n3071) );
  AND3_X1 U2330 ( .A1(n3655), .A2(n3654), .A3(n3653), .ZN(n333) );
  INV_X1 U2331 ( .A(\sra_131/SH[4] ), .ZN(n2847) );
  OR2_X1 U2332 ( .A1(n3172), .A2(n3171), .ZN(\DataP/alu_a_in[17] ) );
  OR2_X1 U2333 ( .A1(n3953), .A2(\CU_I/cw[7] ), .ZN(n3947) );
  NOR3_X1 U2334 ( .A1(n3795), .A2(n3955), .A3(n3837), .ZN(n3953) );
  BUF_X1 U2335 ( .A(n1910), .Z(n2990) );
  INV_X1 U2336 ( .A(n3425), .ZN(\DataP/alu_b_in[16] ) );
  INV_X1 U2337 ( .A(n2005), .ZN(n3003) );
  OR2_X1 U2338 ( .A1(n3026), .A2(n1892), .ZN(n3062) );
  INV_X1 U2339 ( .A(n3987), .ZN(n492) );
  INV_X1 U2340 ( .A(n3988), .ZN(n491) );
  NOR2_X1 U2341 ( .A1(n3853), .A2(n3852), .ZN(\CU_I/cw[7] ) );
  INV_X1 U2342 ( .A(n3951), .ZN(n3853) );
  INV_X1 U2343 ( .A(n3956), .ZN(n3948) );
  INV_X1 U2344 ( .A(n3695), .ZN(n3675) );
  INV_X1 U2345 ( .A(n3674), .ZN(n3691) );
  AND3_X1 U2346 ( .A1(n3201), .A2(n3689), .A3(n3200), .ZN(n3674) );
  OR2_X1 U2347 ( .A1(n3002), .A2(n2229), .ZN(n3101) );
  INV_X1 U2348 ( .A(n3985), .ZN(n494) );
  INV_X1 U2349 ( .A(n3989), .ZN(n490) );
  INV_X1 U2350 ( .A(n3986), .ZN(n493) );
  NOR2_X1 U2351 ( .A1(n487), .A2(n3949), .ZN(\DataP/add_S2[2] ) );
  NOR2_X1 U2352 ( .A1(n486), .A2(n3949), .ZN(\DataP/add_S2[1] ) );
  INV_X1 U2353 ( .A(n2923), .ZN(n2981) );
  BUF_X1 U2354 ( .A(n3703), .Z(n3006) );
  AND4_X1 U2355 ( .A1(n3037), .A2(n1869), .A3(n1999), .A4(n529), .ZN(n2157) );
  NOR2_X1 U2356 ( .A1(n489), .A2(n3949), .ZN(\DataP/add_S2[4] ) );
  NOR2_X1 U2357 ( .A1(n485), .A2(n3949), .ZN(\DataP/add_S2[0] ) );
  NOR2_X1 U2358 ( .A1(n488), .A2(n3949), .ZN(\DataP/add_S2[3] ) );
  NAND2_X1 U2359 ( .A1(n516), .A2(n510), .ZN(n3795) );
  NOR2_X1 U2360 ( .A1(n504), .A2(n497), .ZN(n3966) );
  AND3_X2 U2361 ( .A1(n2453), .A2(n3272), .A3(n2451), .ZN(n3270) );
  OR2_X1 U2362 ( .A1(n2232), .A2(n3003), .ZN(n3097) );
  NOR2_X1 U2363 ( .A1(n3795), .A2(n2141), .ZN(n144) );
  AND2_X1 U2364 ( .A1(BR_EN_i), .A2(n3901), .ZN(n3711) );
  NAND2_X1 U2365 ( .A1(n514), .A2(n515), .ZN(n3955) );
  NAND3_X1 U2366 ( .A1(n3966), .A2(n144), .A3(n2129), .ZN(n3956) );
  NAND2_X2 U2367 ( .A1(n3711), .A2(Rst), .ZN(n3911) );
  NOR2_X1 U2368 ( .A1(n3221), .A2(n3903), .ZN(n3706) );
  OR2_X2 U2369 ( .A1(n3474), .A2(\DataP/alu_a_in[26] ), .ZN(n3504) );
  AND3_X2 U2370 ( .A1(n3468), .A2(n1933), .A3(n1937), .ZN(n2133) );
  AND4_X2 U2371 ( .A1(n3081), .A2(n3083), .A3(n3080), .A4(n3082), .ZN(n3214)
         );
  AND2_X1 U2372 ( .A1(n3198), .A2(ALU_OPCODE_i[1]), .ZN(n3224) );
  BUF_X1 U2373 ( .A(n4021), .Z(n3009) );
  NOR2_X1 U2374 ( .A1(n1448), .A2(n3013), .ZN(n4021) );
  INV_X1 U2375 ( .A(Rst), .ZN(n3014) );
  INV_X1 U2376 ( .A(Rst), .ZN(n3013) );
  INV_X1 U2377 ( .A(\DataP/npc_mux_sel ), .ZN(n3010) );
  BUF_X1 U2378 ( .A(n3944), .Z(n3008) );
  NOR2_X1 U2379 ( .A1(\WB_MUX_SEL_i[1] ), .A2(n294), .ZN(n3944) );
  INV_X1 U2380 ( .A(n3965), .ZN(n3981) );
  NOR2_X1 U2381 ( .A1(n3711), .A2(\DataP/wrong_br ), .ZN(n1448) );
  AND2_X2 U2382 ( .A1(n2503), .A2(n2133), .ZN(n3488) );
  AND4_X2 U2383 ( .A1(n3315), .A2(n2520), .A3(n3313), .A4(n3314), .ZN(n3425)
         );
  AND4_X2 U2384 ( .A1(n3305), .A2(n2519), .A3(n3303), .A4(n3304), .ZN(n3424)
         );
  AND2_X2 U2385 ( .A1(n3420), .A2(n3421), .ZN(n3437) );
  OR2_X2 U2386 ( .A1(n3187), .A2(n3186), .ZN(\DataP/alu_a_in[12] ) );
  OR2_X2 U2387 ( .A1(n3122), .A2(n3121), .ZN(\DataP/alu_a_in[5] ) );
  INV_X2 U2388 ( .A(n3694), .ZN(n3697) );
  INV_X2 U2389 ( .A(n1857), .ZN(n2991) );
  BUF_X2 U2390 ( .A(n3194), .Z(n2563) );
  OR2_X2 U2391 ( .A1(n3125), .A2(n3124), .ZN(\DataP/alu_a_in[6] ) );
  INV_X2 U2392 ( .A(n1857), .ZN(n2992) );
  BUF_X2 U2393 ( .A(n1887), .Z(n3000) );
  NOR4_X1 U2394 ( .A1(n443), .A2(ALU_OPCODE_i[3]), .A3(ALU_OPCODE_i[2]), .A4(
        ALU_OPCODE_i[1]), .ZN(n3901) );
  NAND2_X1 U2395 ( .A1(n3226), .A2(ALU_OPCODE_i[0]), .ZN(n3709) );
  AOI211_X1 U2396 ( .C1(n3675), .C2(\DataP/ALU_C/shifter/N83 ), .A(n3369), .B(
        n3368), .ZN(n358) );
  AND2_X1 U2397 ( .A1(\DataP/ALU_C/shifter/N51 ), .A2(n3006), .ZN(n3368) );
  OAI211_X1 U2398 ( .C1(n3674), .C2(n3367), .A(n3366), .B(n3365), .ZN(n3369)
         );
  AOI21_X1 U2399 ( .B1(n1939), .B2(n3364), .A(n3363), .ZN(n3365) );
  NAND2_X1 U2400 ( .A1(\DataP/ALU_C/shifter/N19 ), .A2(n3007), .ZN(n3366) );
  INV_X1 U2401 ( .A(n2618), .ZN(n2703) );
  NAND2_X1 U2402 ( .A1(n3359), .A2(n3358), .ZN(n3360) );
  INV_X1 U2403 ( .A(\DataP/add_S2[1] ), .ZN(n2559) );
  AOI21_X1 U2404 ( .B1(n2990), .B2(n3693), .A(n3697), .ZN(n3373) );
  INV_X1 U2405 ( .A(n2673), .ZN(n2704) );
  OAI22_X1 U2406 ( .A1(n355), .A2(n3911), .B1(n3994), .B2(n3910), .ZN(
        \DataP/PC_reg/N6 ) );
  INV_X1 U2407 ( .A(n2691), .ZN(n2705) );
  OAI22_X1 U2408 ( .A1(n356), .A2(n3911), .B1(n3993), .B2(n3910), .ZN(
        \DataP/PC_reg/N5 ) );
  AOI21_X1 U2409 ( .B1(n2330), .B2(n3694), .A(n3679), .ZN(n3680) );
  INV_X1 U2410 ( .A(\DataP/add_S2[3] ), .ZN(n2557) );
  INV_X1 U2411 ( .A(\DataP/add_S2[0] ), .ZN(n2558) );
  OAI22_X1 U2412 ( .A1(n353), .A2(n3911), .B1(n3996), .B2(n3910), .ZN(
        \DataP/PC_reg/N8 ) );
  NAND2_X1 U2413 ( .A1(\DataP/alu_b_in[6] ), .A2(n3660), .ZN(n2363) );
  AOI22_X1 U2414 ( .A1(n3388), .A2(\DataP/alu_b_in[7] ), .B1(n3697), .B2(
        \DataP/alu_a_in[7] ), .ZN(n3389) );
  OAI21_X1 U2415 ( .B1(n1926), .B2(n3671), .A(n3694), .ZN(n3388) );
  INV_X1 U2416 ( .A(n2694), .ZN(n2706) );
  INV_X1 U2417 ( .A(n1888), .ZN(n3386) );
  OAI21_X1 U2418 ( .B1(n3670), .B2(n3378), .A(n1954), .ZN(n3383) );
  INV_X1 U2419 ( .A(n3376), .ZN(n3378) );
  NAND2_X1 U2420 ( .A1(n2001), .A2(n3375), .ZN(n3670) );
  OAI22_X1 U2421 ( .A1(n345), .A2(n3911), .B1(n3998), .B2(n3910), .ZN(
        \DataP/PC_reg/N10 ) );
  AOI21_X1 U2422 ( .B1(n3663), .B2(n1939), .A(n3697), .ZN(n3662) );
  NOR2_X1 U2423 ( .A1(n1939), .A2(n3697), .ZN(n3661) );
  INV_X1 U2424 ( .A(n2695), .ZN(n2707) );
  AOI22_X1 U2425 ( .A1(n3227), .A2(\DataP/alu_b_in[9] ), .B1(n3697), .B2(
        \DataP/alu_a_in[9] ), .ZN(n3228) );
  OAI21_X1 U2426 ( .B1(n1922), .B2(n3671), .A(n3694), .ZN(n3227) );
  INV_X1 U2427 ( .A(n2696), .ZN(n2708) );
  INV_X1 U2428 ( .A(n3657), .ZN(n3217) );
  NOR2_X1 U2429 ( .A1(n3911), .A2(n443), .ZN(n2347) );
  INV_X1 U2430 ( .A(n3243), .ZN(n340) );
  OAI211_X1 U2431 ( .C1(n3674), .C2(n3242), .A(n3241), .B(n3240), .ZN(n3243)
         );
  AOI22_X1 U2432 ( .A1(n3006), .A2(\DataP/ALU_C/shifter/N60 ), .B1(
        \DataP/ALU_C/shifter/N92 ), .B2(n3675), .ZN(n3240) );
  AOI21_X1 U2433 ( .B1(\DataP/ALU_C/shifter/N28 ), .B2(n3007), .A(n3239), .ZN(
        n3241) );
  OAI21_X1 U2434 ( .B1(n3700), .B2(n3283), .A(n3238), .ZN(n3239) );
  AOI22_X1 U2435 ( .A1(n3237), .A2(n1879), .B1(n3697), .B2(
        \DataP/alu_a_in[10] ), .ZN(n3238) );
  OAI21_X1 U2436 ( .B1(n3236), .B2(n3671), .A(n3694), .ZN(n3237) );
  INV_X1 U2437 ( .A(n2654), .ZN(n2697) );
  XNOR2_X1 U2438 ( .A(n3248), .B(n3235), .ZN(n3242) );
  INV_X1 U2439 ( .A(n1985), .ZN(n3234) );
  NAND2_X1 U2440 ( .A1(n2343), .A2(n2342), .ZN(n296) );
  INV_X1 U2441 ( .A(\DataP/ALU_C/comp/N24 ), .ZN(n3352) );
  NAND2_X1 U2442 ( .A1(n2345), .A2(n2344), .ZN(n2343) );
  NOR3_X1 U2443 ( .A1(n2431), .A2(n2349), .A3(n443), .ZN(n2344) );
  NAND4_X1 U2444 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3357)
         );
  OAI21_X1 U2445 ( .B1(n3336), .B2(n3697), .A(n3335), .ZN(n3337) );
  AOI21_X1 U2446 ( .B1(n3674), .B2(n3700), .A(n3361), .ZN(n3336) );
  NAND2_X1 U2447 ( .A1(n3361), .A2(n3693), .ZN(n3338) );
  NAND2_X1 U2448 ( .A1(\DataP/ALU_C/shifter/N50 ), .A2(n3006), .ZN(n3340) );
  OAI21_X1 U2449 ( .B1(n3350), .B2(n3356), .A(n3349), .ZN(n3351) );
  INV_X1 U2450 ( .A(n3355), .ZN(n3349) );
  INV_X1 U2451 ( .A(n1876), .ZN(n3350) );
  AND2_X1 U2452 ( .A1(n3353), .A2(n3223), .ZN(n3341) );
  NAND2_X1 U2453 ( .A1(n2516), .A2(n2369), .ZN(n3353) );
  INV_X1 U2454 ( .A(n3374), .ZN(n3316) );
  XNOR2_X1 U2455 ( .A(\DataP/alu_a_in[2] ), .B(n2844), .ZN(n3374) );
  XNOR2_X1 U2456 ( .A(\DataP/alu_a_in[4] ), .B(\lt_x_134/B[4] ), .ZN(n3673) );
  XNOR2_X1 U2457 ( .A(\DataP/alu_a_in[7] ), .B(\DataP/alu_b_in[7] ), .ZN(n3390) );
  XNOR2_X1 U2458 ( .A(\DataP/alu_a_in[6] ), .B(\DataP/alu_b_in[6] ), .ZN(n3668) );
  INV_X1 U2459 ( .A(n3361), .ZN(n3317) );
  AND2_X1 U2460 ( .A1(n2517), .A2(n3904), .ZN(n2516) );
  NOR3_X1 U2461 ( .A1(n3299), .A2(n3364), .A3(n3298), .ZN(n3904) );
  NAND4_X1 U2462 ( .A1(n3518), .A2(n3527), .A3(n3477), .A4(n3536), .ZN(n3298)
         );
  INV_X1 U2463 ( .A(n3547), .ZN(n3299) );
  NOR2_X1 U2464 ( .A1(n3905), .A2(n2518), .ZN(n2517) );
  NAND4_X1 U2465 ( .A1(n3586), .A2(n3908), .A3(n3909), .A4(n3570), .ZN(n2518)
         );
  AND4_X1 U2466 ( .A1(n3605), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n2222)
         );
  XNOR2_X1 U2467 ( .A(\DataP/alu_a_in[9] ), .B(\DataP/alu_b_in[9] ), .ZN(n3282) );
  XNOR2_X1 U2468 ( .A(\DataP/alu_a_in[10] ), .B(n1879), .ZN(n3283) );
  OAI21_X1 U2469 ( .B1(n3346), .B2(n3345), .A(n3344), .ZN(n3347) );
  OAI22_X1 U2470 ( .A1(n317), .A2(n3911), .B1(n3910), .B2(n4010), .ZN(
        \DataP/PC_reg/N22 ) );
  INV_X1 U2471 ( .A(\DataP/npc[20] ), .ZN(n4010) );
  AOI21_X1 U2472 ( .B1(n3601), .B2(n3691), .A(n3600), .ZN(n317) );
  NAND2_X1 U2473 ( .A1(\DataP/ALU_C/shifter/N38 ), .A2(n3007), .ZN(n3597) );
  AOI21_X1 U2474 ( .B1(\DataP/ALU_C/shifter/N70 ), .B2(n3703), .A(n3596), .ZN(
        n3598) );
  OAI211_X1 U2475 ( .C1(n3907), .C2(n3700), .A(n3595), .B(n3594), .ZN(n3596)
         );
  NAND2_X1 U2476 ( .A1(\DataP/alu_a_in[20] ), .A2(n3697), .ZN(n3594) );
  OAI211_X1 U2477 ( .C1(\DataP/alu_a_in[20] ), .C2(n3697), .A(
        \DataP/alu_b_in[20] ), .B(n3660), .ZN(n3595) );
  XNOR2_X1 U2478 ( .A(\DataP/alu_a_in[20] ), .B(\DataP/alu_b_in[20] ), .ZN(
        n3907) );
  NAND2_X1 U2479 ( .A1(\DataP/ALU_C/shifter/N102 ), .A2(n3675), .ZN(n3599) );
  OAI22_X1 U2480 ( .A1(n326), .A2(n3911), .B1(n3910), .B2(n4006), .ZN(
        \DataP/PC_reg/N18 ) );
  INV_X1 U2481 ( .A(\DataP/npc[16] ), .ZN(n4006) );
  AOI21_X1 U2482 ( .B1(n3630), .B2(n3691), .A(n3629), .ZN(n326) );
  NAND2_X1 U2483 ( .A1(\DataP/ALU_C/shifter/N34 ), .A2(n3007), .ZN(n3626) );
  NAND2_X1 U2484 ( .A1(\DataP/ALU_C/shifter/N98 ), .A2(n3675), .ZN(n3627) );
  INV_X1 U2485 ( .A(n2894), .ZN(\DataP/ALU_C/shifter/N98 ) );
  AOI21_X1 U2486 ( .B1(\DataP/ALU_C/shifter/N66 ), .B2(n3703), .A(n3625), .ZN(
        n3628) );
  OAI211_X1 U2487 ( .C1(n3624), .C2(n3700), .A(n3623), .B(n3622), .ZN(n3625)
         );
  OAI21_X1 U2488 ( .B1(\DataP/alu_a_in[16] ), .B2(\DataP/alu_b_in[16] ), .A(
        n3697), .ZN(n3622) );
  XNOR2_X1 U2489 ( .A(\DataP/alu_a_in[16] ), .B(\DataP/alu_b_in[16] ), .ZN(
        n3624) );
  INV_X1 U2490 ( .A(n3280), .ZN(n337) );
  OAI211_X1 U2491 ( .C1(n3279), .C2(n3674), .A(n3278), .B(n3277), .ZN(n3280)
         );
  AOI22_X1 U2492 ( .A1(\DataP/ALU_C/shifter/N30 ), .A2(n3007), .B1(n3675), 
        .B2(\DataP/ALU_C/shifter/N94 ), .ZN(n3277) );
  INV_X1 U2493 ( .A(n2664), .ZN(n2699) );
  AOI21_X1 U2494 ( .B1(\DataP/ALU_C/shifter/N62 ), .B2(n3006), .A(n3276), .ZN(
        n3278) );
  OAI211_X1 U2495 ( .C1(n3284), .C2(n3700), .A(n3275), .B(n3274), .ZN(n3276)
         );
  OAI21_X1 U2496 ( .B1(\DataP/alu_a_in[12] ), .B2(n1880), .A(n3697), .ZN(n3275) );
  XNOR2_X1 U2497 ( .A(\DataP/alu_a_in[12] ), .B(n1880), .ZN(n3284) );
  NAND2_X1 U2498 ( .A1(n3642), .A2(n3640), .ZN(n3273) );
  NAND2_X1 U2499 ( .A1(\DataP/ALU_C/shifter/N29 ), .A2(n3007), .ZN(n3257) );
  INV_X1 U2500 ( .A(n2658), .ZN(n2698) );
  AOI21_X1 U2501 ( .B1(n3318), .B2(n1939), .A(n3256), .ZN(n3258) );
  OAI22_X1 U2502 ( .A1(n3255), .A2(n3254), .B1(n1863), .B2(n3694), .ZN(n3256)
         );
  AOI21_X1 U2503 ( .B1(\DataP/alu_a_in[11] ), .B2(n3693), .A(n3697), .ZN(n3255) );
  AOI22_X1 U2504 ( .A1(n3006), .A2(\DataP/ALU_C/shifter/N61 ), .B1(
        \DataP/ALU_C/shifter/N93 ), .B2(n3675), .ZN(n3259) );
  NAND2_X1 U2505 ( .A1(n3253), .A2(n3691), .ZN(n3260) );
  XNOR2_X1 U2506 ( .A(n3252), .B(n3270), .ZN(n3253) );
  NAND2_X1 U2507 ( .A1(n2012), .A2(n3265), .ZN(n3659) );
  OAI22_X1 U2508 ( .A1(n333), .A2(n3911), .B1(n3910), .B2(n4003), .ZN(
        \DataP/PC_reg/N15 ) );
  INV_X1 U2509 ( .A(\DataP/npc[13] ), .ZN(n4003) );
  AOI22_X1 U2510 ( .A1(n3006), .A2(\DataP/ALU_C/shifter/N63 ), .B1(
        \DataP/ALU_C/shifter/N95 ), .B2(n3675), .ZN(n3653) );
  AOI21_X1 U2511 ( .B1(\DataP/ALU_C/shifter/N31 ), .B2(n3007), .A(n3652), .ZN(
        n3654) );
  OAI211_X1 U2512 ( .C1(n3651), .C2(n3700), .A(n3650), .B(n3649), .ZN(n3652)
         );
  INV_X1 U2513 ( .A(n2671), .ZN(n2700) );
  OAI211_X1 U2514 ( .C1(n3648), .C2(n3647), .A(n3646), .B(n3691), .ZN(n3655)
         );
  OAI211_X1 U2515 ( .C1(n3645), .C2(n3644), .A(n3643), .B(n3642), .ZN(n3646)
         );
  NAND2_X1 U2516 ( .A1(n1601), .A2(n3640), .ZN(n3643) );
  NOR2_X1 U2517 ( .A1(n1997), .A2(n3639), .ZN(n3648) );
  OAI22_X1 U2518 ( .A1(n301), .A2(n3911), .B1(n3910), .B2(n4017), .ZN(
        \DataP/PC_reg/N29 ) );
  INV_X1 U2519 ( .A(\DataP/npc[27] ), .ZN(n4017) );
  NOR2_X1 U2520 ( .A1(n2397), .A2(n3481), .ZN(n2396) );
  OAI211_X1 U2521 ( .C1(n3695), .C2(n2926), .A(n3480), .B(n3479), .ZN(n3481)
         );
  AOI21_X1 U2522 ( .B1(\DataP/ALU_C/shifter/N77 ), .B2(n3006), .A(n3478), .ZN(
        n3479) );
  OAI21_X1 U2523 ( .B1(n3700), .B2(n3477), .A(n3476), .ZN(n3478) );
  AOI22_X1 U2524 ( .A1(n3475), .A2(\DataP/alu_b_in[27] ), .B1(n3697), .B2(
        \DataP/alu_a_in[27] ), .ZN(n3476) );
  OAI21_X1 U2525 ( .B1(n1912), .B2(n3671), .A(n3694), .ZN(n3475) );
  XNOR2_X1 U2526 ( .A(\DataP/alu_a_in[27] ), .B(\DataP/alu_b_in[27] ), .ZN(
        n3477) );
  NAND2_X1 U2527 ( .A1(n2400), .A2(n2398), .ZN(n2397) );
  NAND2_X1 U2528 ( .A1(n1867), .A2(n2399), .ZN(n2398) );
  NOR2_X1 U2529 ( .A1(n3504), .A2(n3674), .ZN(n2399) );
  NAND2_X1 U2530 ( .A1(n2401), .A2(n2553), .ZN(n2400) );
  OR2_X1 U2531 ( .A1(n2422), .A2(n2394), .ZN(n2393) );
  NOR2_X1 U2532 ( .A1(n1867), .A2(n2402), .ZN(n2401) );
  NAND2_X1 U2533 ( .A1(n3504), .A2(n3691), .ZN(n2402) );
  OAI22_X1 U2534 ( .A1(n313), .A2(n3911), .B1(n3910), .B2(n4011), .ZN(
        \DataP/PC_reg/N23 ) );
  INV_X1 U2535 ( .A(\DataP/npc[21] ), .ZN(n4011) );
  AOI21_X1 U2536 ( .B1(n3591), .B2(n3691), .A(n3590), .ZN(n313) );
  OAI21_X1 U2537 ( .B1(n3695), .B2(n3589), .A(n3588), .ZN(n3590) );
  AOI21_X1 U2538 ( .B1(n3007), .B2(\DataP/ALU_C/shifter/N39 ), .A(n3587), .ZN(
        n3588) );
  OAI211_X1 U2539 ( .C1(n3700), .C2(n3586), .A(n3585), .B(n3584), .ZN(n3587)
         );
  AOI22_X1 U2540 ( .A1(n3583), .A2(\DataP/alu_b_in[21] ), .B1(n3697), .B2(
        \DataP/alu_a_in[21] ), .ZN(n3584) );
  OAI21_X1 U2541 ( .B1(n1589), .B2(n3671), .A(n3694), .ZN(n3583) );
  NAND2_X1 U2542 ( .A1(\DataP/ALU_C/shifter/N71 ), .A2(n3006), .ZN(n3585) );
  XNOR2_X1 U2543 ( .A(\DataP/alu_a_in[21] ), .B(\DataP/alu_b_in[21] ), .ZN(
        n3586) );
  INV_X1 U2544 ( .A(\DataP/ALU_C/shifter/N103 ), .ZN(n3589) );
  AOI21_X1 U2545 ( .B1(n1989), .B2(n3580), .A(n3579), .ZN(n3581) );
  INV_X1 U2546 ( .A(n1560), .ZN(n3579) );
  OAI22_X1 U2547 ( .A1(n304), .A2(n3911), .B1(n3910), .B2(n4015), .ZN(
        \DataP/PC_reg/N27 ) );
  INV_X1 U2548 ( .A(\DataP/npc[25] ), .ZN(n4015) );
  AOI21_X1 U2549 ( .B1(n3553), .B2(n3691), .A(n3552), .ZN(n304) );
  AOI21_X1 U2550 ( .B1(\DataP/ALU_C/shifter/N75 ), .B2(n3703), .A(n3548), .ZN(
        n3549) );
  XNOR2_X1 U2551 ( .A(\DataP/alu_a_in[25] ), .B(\DataP/alu_b_in[25] ), .ZN(
        n3547) );
  NAND2_X1 U2552 ( .A1(\DataP/ALU_C/shifter/N43 ), .A2(n3007), .ZN(n3550) );
  NAND2_X1 U2553 ( .A1(\DataP/ALU_C/shifter/N107 ), .A2(n3675), .ZN(n3551) );
  INV_X1 U2554 ( .A(n2922), .ZN(n2984) );
  NOR2_X1 U2555 ( .A1(n2556), .A2(n3544), .ZN(n3546) );
  OAI22_X1 U2556 ( .A1(n311), .A2(n3911), .B1(n3910), .B2(n4012), .ZN(
        \DataP/PC_reg/N24 ) );
  INV_X1 U2557 ( .A(\DataP/npc[22] ), .ZN(n4012) );
  AOI21_X1 U2558 ( .B1(n3575), .B2(n3691), .A(n3574), .ZN(n311) );
  OAI21_X1 U2559 ( .B1(n3695), .B2(n3573), .A(n3572), .ZN(n3574) );
  AOI21_X1 U2560 ( .B1(n3007), .B2(\DataP/ALU_C/shifter/N40 ), .A(n3571), .ZN(
        n3572) );
  OAI211_X1 U2561 ( .C1(n3700), .C2(n3570), .A(n3569), .B(n3568), .ZN(n3571)
         );
  AOI22_X1 U2562 ( .A1(n3567), .A2(\DataP/alu_b_in[22] ), .B1(n3697), .B2(
        \DataP/alu_a_in[22] ), .ZN(n3568) );
  OAI21_X1 U2563 ( .B1(n3566), .B2(n3671), .A(n3694), .ZN(n3567) );
  NAND2_X1 U2564 ( .A1(\DataP/ALU_C/shifter/N72 ), .A2(n3006), .ZN(n3569) );
  XNOR2_X1 U2565 ( .A(\DataP/alu_a_in[22] ), .B(\DataP/alu_b_in[22] ), .ZN(
        n3570) );
  INV_X1 U2566 ( .A(\DataP/ALU_C/shifter/N104 ), .ZN(n3573) );
  XNOR2_X1 U2567 ( .A(n1639), .B(n3564), .ZN(n3575) );
  OAI22_X1 U2568 ( .A1(n308), .A2(n3911), .B1(n3910), .B2(n4014), .ZN(
        \DataP/PC_reg/N26 ) );
  INV_X1 U2569 ( .A(\DataP/npc[24] ), .ZN(n4014) );
  AOI21_X1 U2570 ( .B1(n3563), .B2(n3691), .A(n3562), .ZN(n308) );
  NAND2_X1 U2571 ( .A1(\DataP/ALU_C/shifter/N42 ), .A2(n3007), .ZN(n3559) );
  AOI21_X1 U2572 ( .B1(\DataP/ALU_C/shifter/N74 ), .B2(n3703), .A(n3558), .ZN(
        n3560) );
  OAI211_X1 U2573 ( .C1(n3909), .C2(n3700), .A(n3557), .B(n3556), .ZN(n3558)
         );
  NAND2_X1 U2574 ( .A1(\DataP/alu_a_in[24] ), .A2(n3697), .ZN(n3556) );
  OAI211_X1 U2575 ( .C1(\DataP/alu_a_in[24] ), .C2(n3697), .A(
        \DataP/alu_b_in[24] ), .B(n3660), .ZN(n3557) );
  XNOR2_X1 U2576 ( .A(\DataP/alu_a_in[24] ), .B(\DataP/alu_b_in[24] ), .ZN(
        n3909) );
  NAND2_X1 U2577 ( .A1(\DataP/ALU_C/shifter/N106 ), .A2(n3675), .ZN(n3561) );
  INV_X1 U2578 ( .A(n2919), .ZN(n2983) );
  XNOR2_X1 U2579 ( .A(n2423), .B(n2158), .ZN(n3563) );
  OAI22_X1 U2580 ( .A1(n323), .A2(n3911), .B1(n3910), .B2(n4007), .ZN(
        \DataP/PC_reg/N19 ) );
  INV_X1 U2581 ( .A(\DataP/npc[17] ), .ZN(n4007) );
  AOI21_X1 U2582 ( .B1(n3621), .B2(n3691), .A(n3620), .ZN(n323) );
  AOI21_X1 U2583 ( .B1(\DataP/ALU_C/shifter/N67 ), .B2(n3703), .A(n3616), .ZN(
        n3618) );
  OAI211_X1 U2584 ( .C1(n3615), .C2(n3700), .A(n3614), .B(n3613), .ZN(n3616)
         );
  OAI211_X1 U2585 ( .C1(\DataP/alu_a_in[17] ), .C2(n3697), .A(
        \DataP/alu_b_in[17] ), .B(n3660), .ZN(n3613) );
  NAND2_X1 U2586 ( .A1(\DataP/alu_a_in[17] ), .A2(n3697), .ZN(n3614) );
  XNOR2_X1 U2587 ( .A(\DataP/alu_a_in[17] ), .B(\DataP/alu_b_in[17] ), .ZN(
        n3615) );
  NAND2_X1 U2588 ( .A1(\DataP/ALU_C/shifter/N99 ), .A2(n3675), .ZN(n3619) );
  OAI22_X1 U2589 ( .A1(n303), .A2(n3911), .B1(n3910), .B2(n4016), .ZN(
        \DataP/PC_reg/N28 ) );
  INV_X1 U2590 ( .A(\DataP/npc[26] ), .ZN(n4016) );
  AOI21_X1 U2591 ( .B1(n3542), .B2(n3691), .A(n3541), .ZN(n303) );
  AOI21_X1 U2592 ( .B1(\DataP/ALU_C/shifter/N76 ), .B2(n3703), .A(n3537), .ZN(
        n3539) );
  OAI211_X1 U2593 ( .C1(n3536), .C2(n3700), .A(n3535), .B(n3534), .ZN(n3537)
         );
  NAND2_X1 U2594 ( .A1(\DataP/alu_a_in[26] ), .A2(n3697), .ZN(n3534) );
  OAI211_X1 U2595 ( .C1(\DataP/alu_a_in[26] ), .C2(n3697), .A(
        \DataP/alu_b_in[26] ), .B(n3660), .ZN(n3535) );
  XNOR2_X1 U2596 ( .A(\DataP/alu_a_in[26] ), .B(\DataP/alu_b_in[26] ), .ZN(
        n3536) );
  XNOR2_X1 U2597 ( .A(n1590), .B(n3533), .ZN(n3542) );
  INV_X1 U2598 ( .A(n3472), .ZN(n2421) );
  OAI21_X1 U2599 ( .B1(n3544), .B2(n3555), .A(n3543), .ZN(n3472) );
  INV_X1 U2600 ( .A(n3502), .ZN(n3555) );
  INV_X1 U2601 ( .A(n3497), .ZN(n3465) );
  INV_X1 U2602 ( .A(\DataP/npc[28] ), .ZN(n4018) );
  OAI211_X1 U2603 ( .C1(n3695), .C2(n2928), .A(n3530), .B(n3529), .ZN(n3531)
         );
  AOI21_X1 U2604 ( .B1(\DataP/ALU_C/shifter/N78 ), .B2(n3703), .A(n3528), .ZN(
        n3529) );
  OAI21_X1 U2605 ( .B1(n3700), .B2(n3527), .A(n3526), .ZN(n3528) );
  AOI22_X1 U2606 ( .A1(n3525), .A2(\DataP/alu_b_in[28] ), .B1(n3697), .B2(
        \DataP/alu_a_in[28] ), .ZN(n3526) );
  OAI21_X1 U2607 ( .B1(n1811), .B2(n3671), .A(n3694), .ZN(n3525) );
  XNOR2_X1 U2608 ( .A(\DataP/alu_a_in[28] ), .B(\DataP/alu_b_in[28] ), .ZN(
        n3527) );
  NAND2_X1 U2609 ( .A1(\DataP/ALU_C/shifter/N46 ), .A2(n3007), .ZN(n3530) );
  XNOR2_X1 U2610 ( .A(n3523), .B(n1811), .ZN(n3524) );
  INV_X1 U2611 ( .A(\DataP/npc[23] ), .ZN(n4013) );
  AOI21_X1 U2612 ( .B1(n3455), .B2(n3691), .A(n3454), .ZN(n309) );
  OAI211_X1 U2613 ( .C1(n3453), .C2(n3695), .A(n3452), .B(n3451), .ZN(n3454)
         );
  AOI21_X1 U2614 ( .B1(\DataP/ALU_C/shifter/N73 ), .B2(n3703), .A(n3450), .ZN(
        n3452) );
  OAI211_X1 U2615 ( .C1(n3908), .C2(n3700), .A(n3449), .B(n3448), .ZN(n3450)
         );
  NAND2_X1 U2616 ( .A1(\DataP/alu_a_in[23] ), .A2(n3697), .ZN(n3448) );
  OAI211_X1 U2617 ( .C1(\DataP/alu_a_in[23] ), .C2(n3697), .A(
        \DataP/alu_b_in[23] ), .B(n3660), .ZN(n3449) );
  XNOR2_X1 U2618 ( .A(\DataP/alu_a_in[23] ), .B(\DataP/alu_b_in[23] ), .ZN(
        n3908) );
  INV_X1 U2619 ( .A(\DataP/ALU_C/shifter/N105 ), .ZN(n3453) );
  INV_X1 U2620 ( .A(n2917), .ZN(n2982) );
  AND2_X1 U2621 ( .A1(n2527), .A2(n2524), .ZN(n2523) );
  NAND2_X1 U2622 ( .A1(n2526), .A2(n2525), .ZN(n2524) );
  NOR2_X1 U2623 ( .A1(n3456), .A2(n1893), .ZN(n2525) );
  AND2_X1 U2624 ( .A1(n1998), .A2(n1610), .ZN(n2527) );
  AND3_X1 U2625 ( .A1(n1559), .A2(n1557), .A3(n1959), .ZN(n2526) );
  INV_X1 U2626 ( .A(\DataP/npc[31] ), .ZN(n4023) );
  OAI22_X1 U2627 ( .A1(n319), .A2(n3911), .B1(n3910), .B2(n4009), .ZN(
        \DataP/PC_reg/N21 ) );
  INV_X1 U2628 ( .A(\DataP/npc[19] ), .ZN(n4009) );
  AOI21_X1 U2629 ( .B1(n3436), .B2(n3691), .A(n3435), .ZN(n319) );
  NAND2_X1 U2630 ( .A1(\DataP/ALU_C/shifter/N37 ), .A2(n3007), .ZN(n3432) );
  AOI21_X1 U2631 ( .B1(\DataP/ALU_C/shifter/N69 ), .B2(n3006), .A(n3431), .ZN(
        n3433) );
  OAI211_X1 U2632 ( .C1(n3906), .C2(n3700), .A(n3430), .B(n3429), .ZN(n3431)
         );
  NAND2_X1 U2633 ( .A1(n1553), .A2(n3697), .ZN(n3429) );
  OAI211_X1 U2634 ( .C1(n1553), .C2(n3697), .A(\DataP/alu_b_in[19] ), .B(n3660), .ZN(n3430) );
  XNOR2_X1 U2635 ( .A(n1553), .B(\DataP/alu_b_in[19] ), .ZN(n3906) );
  NAND2_X1 U2636 ( .A1(\DataP/ALU_C/shifter/N101 ), .A2(n3675), .ZN(n3434) );
  AOI21_X1 U2637 ( .B1(n2226), .B2(n1919), .A(n2223), .ZN(n2411) );
  INV_X1 U2638 ( .A(\DataP/npc[30] ), .ZN(n4020) );
  NOR2_X1 U2639 ( .A1(n3674), .A2(n3911), .ZN(n2412) );
  OAI22_X1 U2640 ( .A1(n322), .A2(n3911), .B1(n3910), .B2(n4008), .ZN(
        \DataP/PC_reg/N20 ) );
  INV_X1 U2641 ( .A(\DataP/npc[18] ), .ZN(n4008) );
  INV_X1 U2642 ( .A(n3610), .ZN(n322) );
  OAI211_X1 U2643 ( .C1(n3609), .C2(n3674), .A(n3608), .B(n3607), .ZN(n3610)
         );
  NAND2_X1 U2644 ( .A1(\DataP/ALU_C/shifter/N100 ), .A2(n3675), .ZN(n3607) );
  AOI21_X1 U2645 ( .B1(n3007), .B2(\DataP/ALU_C/shifter/N36 ), .A(n3606), .ZN(
        n3608) );
  OAI211_X1 U2646 ( .C1(n3700), .C2(n3605), .A(n3604), .B(n3603), .ZN(n3606)
         );
  AOI22_X1 U2647 ( .A1(n3602), .A2(\DataP/alu_b_in[18] ), .B1(n3697), .B2(
        \DataP/alu_a_in[18] ), .ZN(n3603) );
  OAI21_X1 U2648 ( .B1(n1884), .B2(n3671), .A(n3694), .ZN(n3602) );
  NAND2_X1 U2649 ( .A1(\DataP/ALU_C/shifter/N68 ), .A2(n3006), .ZN(n3604) );
  XNOR2_X1 U2650 ( .A(\DataP/alu_a_in[18] ), .B(\DataP/alu_b_in[18] ), .ZN(
        n3605) );
  INV_X1 U2651 ( .A(n3441), .ZN(n3423) );
  OAI22_X1 U2652 ( .A1(n332), .A2(n3911), .B1(n3910), .B2(n4004), .ZN(
        \DataP/PC_reg/N16 ) );
  INV_X1 U2653 ( .A(\DataP/npc[14] ), .ZN(n4004) );
  INV_X1 U2654 ( .A(n3638), .ZN(n332) );
  OAI211_X1 U2655 ( .C1(n3637), .C2(n3674), .A(n3636), .B(n3635), .ZN(n3638)
         );
  AOI22_X1 U2656 ( .A1(\DataP/ALU_C/shifter/N32 ), .A2(n3706), .B1(n3675), 
        .B2(\DataP/ALU_C/shifter/N96 ), .ZN(n3635) );
  INV_X1 U2657 ( .A(n2680), .ZN(n2701) );
  AOI21_X1 U2658 ( .B1(\DataP/ALU_C/shifter/N64 ), .B2(n3006), .A(n3634), .ZN(
        n3636) );
  XNOR2_X1 U2659 ( .A(\DataP/alu_a_in[14] ), .B(n1932), .ZN(n3633) );
  XNOR2_X1 U2660 ( .A(n3632), .B(n3631), .ZN(n3637) );
  OAI21_X1 U2661 ( .B1(n2939), .B2(n3695), .A(n3486), .ZN(n3512) );
  AOI21_X1 U2662 ( .B1(\DataP/ALU_C/shifter/N80 ), .B2(n3006), .A(n3485), .ZN(
        n3486) );
  OAI211_X1 U2663 ( .C1(n3484), .C2(n3700), .A(n3483), .B(n3482), .ZN(n3485)
         );
  NAND2_X1 U2664 ( .A1(\DataP/alu_a_in[30] ), .A2(n3697), .ZN(n3482) );
  OAI211_X1 U2665 ( .C1(\DataP/alu_a_in[30] ), .C2(n3697), .A(
        \DataP/alu_b_in[30] ), .B(n3660), .ZN(n3483) );
  XNOR2_X1 U2666 ( .A(\DataP/alu_a_in[30] ), .B(\DataP/alu_b_in[30] ), .ZN(
        n3484) );
  NAND2_X1 U2667 ( .A1(n3705), .A2(n3683), .ZN(n3511) );
  OAI22_X1 U2668 ( .A1(n330), .A2(n3911), .B1(n3910), .B2(n4005), .ZN(
        \DataP/PC_reg/N17 ) );
  INV_X1 U2669 ( .A(\DataP/npc[15] ), .ZN(n4005) );
  AOI21_X1 U2670 ( .B1(n2385), .B2(n3691), .A(n2384), .ZN(n330) );
  NAND2_X1 U2671 ( .A1(n3406), .A2(n3407), .ZN(n2384) );
  AOI21_X1 U2672 ( .B1(\DataP/ALU_C/shifter/N65 ), .B2(n3006), .A(n3405), .ZN(
        n3407) );
  OAI211_X1 U2673 ( .C1(n1842), .C2(n3694), .A(n3404), .B(n3403), .ZN(n3405)
         );
  NAND2_X1 U2674 ( .A1(n3694), .A2(n3671), .ZN(n3660) );
  NAND2_X1 U2675 ( .A1(n3402), .A2(n1939), .ZN(n3404) );
  AOI22_X1 U2676 ( .A1(\DataP/ALU_C/shifter/N33 ), .A2(n3706), .B1(n3675), 
        .B2(\DataP/ALU_C/shifter/N97 ), .ZN(n3406) );
  INV_X1 U2677 ( .A(n2688), .ZN(n2702) );
  XNOR2_X1 U2678 ( .A(n2386), .B(n3413), .ZN(n2385) );
  OAI21_X1 U2679 ( .B1(n3632), .B2(n3414), .A(n3410), .ZN(n2386) );
  AOI21_X1 U2680 ( .B1(n3399), .B2(n3409), .A(n3644), .ZN(n3632) );
  INV_X1 U2681 ( .A(n3408), .ZN(n3644) );
  OAI21_X1 U2682 ( .B1(n3641), .B2(n3394), .A(n3640), .ZN(n3399) );
  OAI21_X1 U2683 ( .B1(n3264), .B2(n2481), .A(n1529), .ZN(n3640) );
  INV_X1 U2684 ( .A(n3642), .ZN(n3394) );
  NAND2_X1 U2685 ( .A1(n2288), .A2(n2294), .ZN(n3642) );
  NAND2_X1 U2686 ( .A1(n3264), .A2(n3510), .ZN(n2288) );
  INV_X1 U2687 ( .A(\DataP/npc[29] ), .ZN(n4019) );
  INV_X1 U2688 ( .A(n3711), .ZN(n3229) );
  OAI211_X1 U2689 ( .C1(n3695), .C2(n2930), .A(n3521), .B(n3520), .ZN(n3522)
         );
  AOI21_X1 U2690 ( .B1(\DataP/ALU_C/shifter/N79 ), .B2(n3703), .A(n3519), .ZN(
        n3520) );
  OAI21_X1 U2691 ( .B1(n3700), .B2(n3518), .A(n3517), .ZN(n3519) );
  AOI22_X1 U2692 ( .A1(n3516), .A2(\DataP/alu_b_in[29] ), .B1(n3697), .B2(
        \DataP/alu_a_in[29] ), .ZN(n3517) );
  OAI21_X1 U2693 ( .B1(n1925), .B2(n3671), .A(n3694), .ZN(n3516) );
  XNOR2_X1 U2694 ( .A(\DataP/alu_a_in[29] ), .B(\DataP/alu_b_in[29] ), .ZN(
        n3518) );
  NAND2_X1 U2695 ( .A1(\DataP/ALU_C/shifter/N47 ), .A2(n3007), .ZN(n3521) );
  INV_X1 U2696 ( .A(n2514), .ZN(n3514) );
  INV_X1 U2697 ( .A(n3513), .ZN(n3515) );
  OAI21_X1 U2698 ( .B1(n2371), .B2(n2321), .A(n2280), .ZN(n3513) );
  INV_X1 U2699 ( .A(n2515), .ZN(n2426) );
  AND2_X1 U2700 ( .A1(n2550), .A2(n2147), .ZN(n2430) );
  AOI21_X1 U2701 ( .B1(n2417), .B2(n2416), .A(n2414), .ZN(n3707) );
  NAND2_X1 U2702 ( .A1(n2415), .A2(n3704), .ZN(n2414) );
  AOI21_X1 U2703 ( .B1(\DataP/ALU_C/shifter/N81 ), .B2(n3006), .A(n3702), .ZN(
        n3704) );
  OAI21_X1 U2704 ( .B1(n3701), .B2(n3700), .A(n3699), .ZN(n3702) );
  AOI22_X1 U2705 ( .A1(\DataP/alu_a_in[31] ), .A2(n3698), .B1(n3697), .B2(
        \DataP/alu_b_in[31] ), .ZN(n3699) );
  NAND2_X1 U2706 ( .A1(n3226), .A2(n3343), .ZN(n3694) );
  INV_X1 U2707 ( .A(n3903), .ZN(n3222) );
  NAND2_X1 U2708 ( .A1(\DataP/alu_b_in[31] ), .A2(n3693), .ZN(n3696) );
  INV_X1 U2709 ( .A(n3671), .ZN(n3693) );
  OR2_X1 U2710 ( .A1(n3225), .A2(n3345), .ZN(n3671) );
  INV_X1 U2711 ( .A(n3224), .ZN(n3225) );
  NOR2_X1 U2712 ( .A1(n3015), .A2(ALU_OPCODE_i[1]), .ZN(n3226) );
  NAND2_X1 U2713 ( .A1(ALU_OPCODE_i[2]), .A2(n443), .ZN(n3015) );
  NAND2_X1 U2714 ( .A1(\DataP/ALU_C/shifter/N49 ), .A2(n3007), .ZN(n2415) );
  INV_X1 U2715 ( .A(n3343), .ZN(n3221) );
  NOR2_X1 U2716 ( .A1(n3692), .A2(n3674), .ZN(n2416) );
  INV_X1 U2717 ( .A(n3705), .ZN(n2417) );
  XNOR2_X1 U2718 ( .A(ALU_OPCODE_i[2]), .B(n3902), .ZN(n3199) );
  NAND2_X1 U2719 ( .A1(n3197), .A2(n3348), .ZN(n3201) );
  NOR2_X1 U2720 ( .A1(ALU_OPCODE_i[2]), .A2(ALU_OPCODE_i[1]), .ZN(n3348) );
  OAI21_X1 U2721 ( .B1(n443), .B2(ALU_OPCODE_i[3]), .A(n3345), .ZN(n3197) );
  NAND2_X1 U2722 ( .A1(n3493), .A2(n1924), .ZN(n3705) );
  INV_X1 U2723 ( .A(n3687), .ZN(n3701) );
  XNOR2_X1 U2724 ( .A(n3688), .B(n3687), .ZN(n3690) );
  XNOR2_X1 U2725 ( .A(\DataP/alu_a_in[31] ), .B(n1935), .ZN(n3687) );
  NOR2_X1 U2726 ( .A1(n2562), .A2(n2191), .ZN(n3130) );
  OAI21_X1 U2727 ( .B1(n1837), .B2(n1), .A(n3129), .ZN(n3131) );
  OR2_X1 U2728 ( .A1(n3686), .A2(\DataP/alu_b_in[30] ), .ZN(n3688) );
  INV_X1 U2729 ( .A(n3683), .ZN(n3684) );
  NOR2_X1 U2730 ( .A1(n2563), .A2(n2192), .ZN(n3133) );
  OAI21_X1 U2731 ( .B1(n2999), .B2(n5), .A(n3132), .ZN(n3134) );
  XNOR2_X1 U2732 ( .A(n3686), .B(\DataP/alu_b_in[30] ), .ZN(n3491) );
  NAND2_X1 U2733 ( .A1(n3490), .A2(n3489), .ZN(n3686) );
  NOR2_X1 U2734 ( .A1(\DataP/alu_b_in[29] ), .A2(\DataP/alu_b_in[28] ), .ZN(
        n3489) );
  INV_X1 U2735 ( .A(\DataP/alu_b_in[30] ), .ZN(n3492) );
  AND2_X1 U2736 ( .A1(n2429), .A2(n2513), .ZN(n2427) );
  NAND2_X1 U2737 ( .A1(n2515), .A2(n2514), .ZN(n2429) );
  NAND2_X1 U2738 ( .A1(n2278), .A2(n2279), .ZN(n2514) );
  NAND2_X1 U2739 ( .A1(n2371), .A2(n2407), .ZN(n2278) );
  AND2_X1 U2740 ( .A1(n2513), .A2(n2147), .ZN(n2428) );
  NOR2_X1 U2741 ( .A1(n2563), .A2(n2206), .ZN(n3139) );
  OAI21_X1 U2742 ( .B1(n2999), .B2(n13), .A(n3138), .ZN(n3140) );
  AOI22_X1 U2743 ( .A1(n2995), .A2(\DataP/alu_out_M[28] ), .B1(n2991), .B2(
        \DataP/alu_out_W[28] ), .ZN(n3138) );
  NOR2_X1 U2744 ( .A1(n1925), .A2(n2281), .ZN(n2280) );
  NOR2_X1 U2745 ( .A1(n2561), .A2(n2199), .ZN(n3136) );
  OAI21_X1 U2746 ( .B1(n2999), .B2(n9), .A(n3135), .ZN(n3137) );
  AOI22_X1 U2747 ( .A1(n2996), .A2(\DataP/alu_out_M[29] ), .B1(n2992), .B2(
        \DataP/alu_out_W[29] ), .ZN(n3135) );
  NAND4_X1 U2748 ( .A1(n3306), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(
        \DataP/alu_b_in[28] ) );
  NAND2_X1 U2749 ( .A1(n3005), .A2(\DataP/alu_out_W[28] ), .ZN(n3292) );
  OR2_X1 U2750 ( .A1(n1636), .A2(n2178), .ZN(n3293) );
  NAND2_X1 U2751 ( .A1(n3001), .A2(\DataP/B_s[28] ), .ZN(n3294) );
  NOR2_X1 U2752 ( .A1(n3487), .A2(\DataP/alu_b_in[27] ), .ZN(n3509) );
  NAND2_X1 U2753 ( .A1(n3507), .A2(\DataP/alu_a_in[27] ), .ZN(n3508) );
  NAND2_X1 U2754 ( .A1(n2474), .A2(n2473), .ZN(n3507) );
  INV_X1 U2755 ( .A(n1548), .ZN(n2554) );
  NOR2_X1 U2756 ( .A1(n2563), .A2(n2193), .ZN(n3142) );
  OAI21_X1 U2757 ( .B1(n1837), .B2(n17), .A(n3141), .ZN(n3143) );
  AOI22_X1 U2758 ( .A1(n2996), .A2(\DataP/alu_out_M[27] ), .B1(n2991), .B2(
        \DataP/alu_out_W[27] ), .ZN(n3141) );
  INV_X1 U2759 ( .A(n3487), .ZN(n2497) );
  NAND2_X1 U2760 ( .A1(n2241), .A2(n1936), .ZN(n3487) );
  NAND4_X1 U2761 ( .A1(n3306), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(
        \DataP/alu_b_in[27] ) );
  NAND2_X1 U2762 ( .A1(n3005), .A2(\DataP/alu_out_W[27] ), .ZN(n3295) );
  OR2_X1 U2763 ( .A1(n2566), .A2(n2165), .ZN(n3296) );
  NAND2_X1 U2764 ( .A1(n1859), .A2(\DataP/B_s[27] ), .ZN(n3297) );
  OR2_X1 U2765 ( .A1(n3532), .A2(n2556), .ZN(n2555) );
  NOR2_X1 U2766 ( .A1(n2563), .A2(n2207), .ZN(n3148) );
  OAI21_X1 U2767 ( .B1(n2999), .B2(n25), .A(n3147), .ZN(n3149) );
  AOI22_X1 U2768 ( .A1(n2996), .A2(\DataP/alu_out_M[25] ), .B1(n2991), .B2(
        \DataP/alu_out_W[25] ), .ZN(n3147) );
  NOR2_X1 U2769 ( .A1(n2563), .A2(n2200), .ZN(n3145) );
  OAI21_X1 U2770 ( .B1(n3000), .B2(n21), .A(n3144), .ZN(n3146) );
  AOI22_X1 U2771 ( .A1(n2995), .A2(\DataP/alu_out_M[26] ), .B1(n2991), .B2(
        \DataP/alu_out_W[26] ), .ZN(n3144) );
  NAND2_X1 U2772 ( .A1(\DataP/alu_b_in[26] ), .A2(n1938), .ZN(n2502) );
  INV_X1 U2773 ( .A(\DataP/alu_b_in[25] ), .ZN(n3473) );
  NAND2_X1 U2774 ( .A1(n2565), .A2(\DataP/IMM_s[31] ), .ZN(n3306) );
  NAND2_X1 U2775 ( .A1(n3471), .A2(\DataP/alu_a_in[24] ), .ZN(n3502) );
  AND2_X1 U2776 ( .A1(n3497), .A2(n3496), .ZN(n2353) );
  NAND2_X1 U2777 ( .A1(n3496), .A2(n3463), .ZN(n3564) );
  NAND2_X1 U2778 ( .A1(n3447), .A2(n3566), .ZN(n3463) );
  INV_X1 U2779 ( .A(\DataP/alu_a_in[22] ), .ZN(n3566) );
  AND2_X1 U2780 ( .A1(n3459), .A2(n1533), .ZN(n2352) );
  AND2_X1 U2781 ( .A1(n3578), .A2(n3580), .ZN(n3593) );
  AOI21_X1 U2782 ( .B1(n3495), .B2(n3497), .A(n3554), .ZN(n3500) );
  NOR2_X1 U2783 ( .A1(n3471), .A2(\DataP/alu_a_in[24] ), .ZN(n3554) );
  NOR2_X1 U2784 ( .A1(n1539), .A2(n2217), .ZN(n3151) );
  OAI21_X1 U2785 ( .B1(n3000), .B2(n29), .A(n3150), .ZN(n3152) );
  AOI22_X1 U2786 ( .A1(n2995), .A2(\DataP/alu_out_M[24] ), .B1(n2991), .B2(
        \DataP/alu_out_W[24] ), .ZN(n3150) );
  XNOR2_X1 U2787 ( .A(n3488), .B(\DataP/alu_b_in[24] ), .ZN(n3469) );
  NAND2_X1 U2788 ( .A1(n3005), .A2(\DataP/alu_out_W[24] ), .ZN(n3319) );
  OR2_X1 U2789 ( .A1(n1636), .A2(n2179), .ZN(n3320) );
  NAND2_X1 U2790 ( .A1(n1905), .A2(\DataP/IMM_s[24] ), .ZN(n3321) );
  NAND2_X1 U2791 ( .A1(n3001), .A2(\DataP/B_s[24] ), .ZN(n3322) );
  XNOR2_X1 U2792 ( .A(n3464), .B(\DataP/alu_a_in[23] ), .ZN(n3495) );
  NOR2_X1 U2793 ( .A1(n1539), .A2(n2194), .ZN(n3154) );
  OAI21_X1 U2794 ( .B1(n1837), .B2(n33), .A(n3153), .ZN(n3155) );
  AOI22_X1 U2795 ( .A1(n2995), .A2(\DataP/alu_out_M[23] ), .B1(n2992), .B2(
        \DataP/alu_out_W[23] ), .ZN(n3153) );
  XNOR2_X1 U2796 ( .A(n3439), .B(n1937), .ZN(n3440) );
  INV_X1 U2797 ( .A(n3444), .ZN(n3468) );
  INV_X1 U2798 ( .A(n2382), .ZN(n2380) );
  NAND2_X1 U2799 ( .A1(n1560), .A2(n3576), .ZN(n3443) );
  AND2_X1 U2800 ( .A1(n2382), .A2(\DataP/alu_a_in[21] ), .ZN(n2370) );
  NOR2_X1 U2801 ( .A1(n2563), .A2(n2201), .ZN(n3160) );
  OAI21_X1 U2802 ( .B1(n2999), .B2(n41), .A(n3159), .ZN(n3161) );
  AOI22_X1 U2803 ( .A1(n2995), .A2(\DataP/alu_out_M[21] ), .B1(n2991), .B2(
        \DataP/alu_out_W[21] ), .ZN(n3159) );
  NAND2_X1 U2804 ( .A1(n2007), .A2(\DataP/alu_a_in[20] ), .ZN(n3578) );
  NOR2_X1 U2805 ( .A1(n2561), .A2(n2208), .ZN(n3163) );
  OAI21_X1 U2806 ( .B1(n2999), .B2(n45), .A(n3162), .ZN(n3164) );
  AOI22_X1 U2807 ( .A1(n2995), .A2(\DataP/alu_out_M[20] ), .B1(n2991), .B2(
        \DataP/alu_out_W[20] ), .ZN(n3162) );
  AND3_X1 U2808 ( .A1(n3496), .A2(n1610), .A3(n3456), .ZN(n3457) );
  NOR2_X1 U2809 ( .A1(n2561), .A2(n2218), .ZN(n3157) );
  OAI21_X1 U2810 ( .B1(n2999), .B2(n37), .A(n3156), .ZN(n3158) );
  AOI22_X1 U2811 ( .A1(n2995), .A2(\DataP/alu_out_M[22] ), .B1(n2991), .B2(
        \DataP/alu_out_W[22] ), .ZN(n3156) );
  NAND4_X1 U2812 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(
        \DataP/alu_b_in[22] ) );
  NAND2_X1 U2813 ( .A1(n3005), .A2(\DataP/alu_out_W[22] ), .ZN(n3323) );
  OR2_X1 U2814 ( .A1(n3002), .A2(n2180), .ZN(n3324) );
  NAND2_X1 U2815 ( .A1(n1848), .A2(\DataP/IMM_s[22] ), .ZN(n3325) );
  NAND2_X1 U2816 ( .A1(n3001), .A2(\DataP/B_s[22] ), .ZN(n3326) );
  NAND2_X1 U2817 ( .A1(n3442), .A2(n1556), .ZN(n3444) );
  NAND2_X1 U2818 ( .A1(n3005), .A2(\DataP/alu_out_W[20] ), .ZN(n3285) );
  OR2_X1 U2819 ( .A1(n1636), .A2(n2173), .ZN(n3286) );
  NAND2_X1 U2820 ( .A1(n1905), .A2(\DataP/IMM_s[20] ), .ZN(n3287) );
  NAND2_X1 U2821 ( .A1(n3001), .A2(\DataP/B_s[20] ), .ZN(n3288) );
  NAND2_X1 U2822 ( .A1(n3005), .A2(\DataP/alu_out_W[21] ), .ZN(n3331) );
  OR2_X1 U2823 ( .A1(n3002), .A2(n2172), .ZN(n3332) );
  NAND2_X1 U2824 ( .A1(n1848), .A2(\DataP/IMM_s[21] ), .ZN(n3333) );
  NAND2_X1 U2825 ( .A1(n3001), .A2(\DataP/B_s[21] ), .ZN(n3334) );
  OAI211_X1 U2826 ( .C1(n3441), .C2(n1531), .A(n1877), .B(n1557), .ZN(n3462)
         );
  NOR2_X1 U2827 ( .A1(n2561), .A2(n2202), .ZN(n3166) );
  OAI21_X1 U2828 ( .B1(n3000), .B2(n49), .A(n3165), .ZN(n3167) );
  AOI22_X1 U2829 ( .A1(n2996), .A2(\DataP/alu_out_M[19] ), .B1(n2991), .B2(
        \DataP/alu_out_W[19] ), .ZN(n3165) );
  NAND2_X1 U2830 ( .A1(n2306), .A2(n3291), .ZN(\DataP/alu_b_in[19] ) );
  NAND2_X1 U2831 ( .A1(n3001), .A2(\DataP/B_s[19] ), .ZN(n3291) );
  NAND2_X1 U2832 ( .A1(n3289), .A2(n3290), .ZN(n2307) );
  OR2_X1 U2833 ( .A1(n3002), .A2(n2174), .ZN(n3289) );
  NOR2_X1 U2834 ( .A1(n1539), .A2(n2209), .ZN(n3169) );
  OAI21_X1 U2835 ( .B1(n2999), .B2(n53), .A(n3168), .ZN(n3170) );
  AOI22_X1 U2836 ( .A1(n2996), .A2(\DataP/alu_out_M[18] ), .B1(n2991), .B2(
        \DataP/alu_out_W[18] ), .ZN(n3168) );
  NAND2_X1 U2837 ( .A1(n3001), .A2(\DataP/B_s[18] ), .ZN(n3281) );
  INV_X1 U2838 ( .A(n2245), .ZN(n2439) );
  AOI21_X1 U2839 ( .B1(n2354), .B2(n3611), .A(n2308), .ZN(n3441) );
  OAI211_X1 U2840 ( .C1(n2494), .C2(n2492), .A(n2489), .B(n2491), .ZN(n2299)
         );
  OR2_X1 U2841 ( .A1(n3437), .A2(n2490), .ZN(n2489) );
  NAND2_X1 U2842 ( .A1(n2538), .A2(n3424), .ZN(n2490) );
  INV_X1 U2843 ( .A(n2538), .ZN(n2492) );
  OAI21_X1 U2844 ( .B1(n3422), .B2(n2383), .A(n2465), .ZN(n3611) );
  NOR2_X1 U2845 ( .A1(n2563), .A2(n2219), .ZN(n3174) );
  OAI21_X1 U2846 ( .B1(n2999), .B2(n61), .A(n3173), .ZN(n3175) );
  AOI22_X1 U2847 ( .A1(n2997), .A2(\DataP/alu_out_M[16] ), .B1(n2991), .B2(
        \DataP/alu_out_W[16] ), .ZN(n3173) );
  XNOR2_X1 U2848 ( .A(n1563), .B(\DataP/alu_b_in[16] ), .ZN(n3422) );
  NOR2_X1 U2849 ( .A1(n1539), .A2(n2195), .ZN(n3171) );
  NAND3_X1 U2850 ( .A1(n2488), .A2(n2494), .A3(n2463), .ZN(n2462) );
  NAND2_X1 U2851 ( .A1(n1848), .A2(\DataP/IMM_s[16] ), .ZN(n3314) );
  OR2_X1 U2852 ( .A1(n3002), .A2(n2167), .ZN(n3313) );
  NAND2_X1 U2853 ( .A1(n3005), .A2(\DataP/alu_out_W[16] ), .ZN(n2520) );
  NAND2_X1 U2854 ( .A1(n1839), .A2(\DataP/B_s[16] ), .ZN(n3315) );
  NAND2_X1 U2855 ( .A1(n1905), .A2(\DataP/IMM_s[17] ), .ZN(n3304) );
  OR2_X1 U2856 ( .A1(n2566), .A2(n2170), .ZN(n3303) );
  NAND2_X1 U2857 ( .A1(n3005), .A2(\DataP/alu_out_W[17] ), .ZN(n2519) );
  NAND2_X1 U2858 ( .A1(n1839), .A2(\DataP/B_s[17] ), .ZN(n3305) );
  AND2_X1 U2859 ( .A1(n3417), .A2(n3418), .ZN(n2390) );
  INV_X1 U2860 ( .A(n3413), .ZN(n2541) );
  XNOR2_X1 U2861 ( .A(\DataP/alu_a_in[15] ), .B(n3417), .ZN(n3402) );
  NAND2_X1 U2862 ( .A1(n3392), .A2(n1842), .ZN(n3391) );
  NOR2_X1 U2863 ( .A1(n2561), .A2(n2196), .ZN(n3177) );
  OAI21_X1 U2864 ( .B1(n3000), .B2(n65), .A(n3176), .ZN(n3178) );
  AOI22_X1 U2865 ( .A1(n2997), .A2(\DataP/alu_out_M[15] ), .B1(n2992), .B2(
        \DataP/alu_out_W[15] ), .ZN(n3176) );
  INV_X1 U2866 ( .A(n1881), .ZN(n2482) );
  INV_X1 U2867 ( .A(n3417), .ZN(\DataP/alu_b_in[15] ) );
  NAND2_X1 U2868 ( .A1(n2564), .A2(\DataP/ir_E[15] ), .ZN(n3302) );
  NAND2_X1 U2869 ( .A1(n3004), .A2(\DataP/alu_out_W[15] ), .ZN(n3300) );
  OR2_X1 U2870 ( .A1(n3002), .A2(n2166), .ZN(n3301) );
  NOR2_X1 U2871 ( .A1(n1881), .A2(n1932), .ZN(n2487) );
  AND2_X1 U2872 ( .A1(n3411), .A2(n3410), .ZN(n3631) );
  INV_X1 U2873 ( .A(n3510), .ZN(n2543) );
  NAND2_X1 U2874 ( .A1(n3398), .A2(n1927), .ZN(n3408) );
  AOI21_X1 U2875 ( .B1(n3397), .B2(n3510), .A(n2546), .ZN(n3398) );
  INV_X1 U2876 ( .A(n3411), .ZN(n3414) );
  NAND2_X1 U2877 ( .A1(n3401), .A2(\DataP/alu_a_in[14] ), .ZN(n3411) );
  NOR2_X1 U2878 ( .A1(n1539), .A2(n2203), .ZN(n3180) );
  OAI21_X1 U2879 ( .B1(n3000), .B2(n69), .A(n3179), .ZN(n3181) );
  AOI22_X1 U2880 ( .A1(n2997), .A2(\DataP/alu_out_M[14] ), .B1(n2992), .B2(
        \DataP/alu_out_W[14] ), .ZN(n3179) );
  OAI21_X1 U2881 ( .B1(n2375), .B2(n2376), .A(n2373), .ZN(n2372) );
  NAND2_X1 U2882 ( .A1(n1881), .A2(n2374), .ZN(n2373) );
  NOR2_X1 U2883 ( .A1(n1932), .A2(n2375), .ZN(n2374) );
  NAND2_X1 U2884 ( .A1(n2482), .A2(n1932), .ZN(n2376) );
  INV_X1 U2885 ( .A(n3510), .ZN(n2375) );
  OR2_X1 U2886 ( .A1(n3002), .A2(n2171), .ZN(n3312) );
  NAND2_X1 U2887 ( .A1(n3004), .A2(\DataP/alu_out_W[14] ), .ZN(n3311) );
  INV_X1 U2888 ( .A(n3409), .ZN(n3645) );
  OAI21_X1 U2889 ( .B1(n2546), .B2(n3397), .A(n2149), .ZN(n3409) );
  NAND2_X1 U2890 ( .A1(n2548), .A2(n2545), .ZN(n2544) );
  INV_X1 U2891 ( .A(n3510), .ZN(n2545) );
  NOR2_X1 U2892 ( .A1(n1539), .A2(n2210), .ZN(n3183) );
  OAI21_X1 U2893 ( .B1(n3000), .B2(n73), .A(n3182), .ZN(n3184) );
  AOI22_X1 U2894 ( .A1(n2997), .A2(\DataP/alu_out_M[13] ), .B1(n2991), .B2(
        \DataP/alu_out_W[13] ), .ZN(n3182) );
  NAND2_X1 U2895 ( .A1(n2006), .A2(\DataP/alu_out_W[13] ), .ZN(n3307) );
  OR2_X1 U2896 ( .A1(n2566), .A2(n2176), .ZN(n3308) );
  NAND2_X1 U2897 ( .A1(n1848), .A2(\DataP/ir_E[13] ), .ZN(n3309) );
  NAND2_X1 U2898 ( .A1(n1839), .A2(\DataP/B_s[13] ), .ZN(n3310) );
  AND2_X1 U2899 ( .A1(n1903), .A2(n2442), .ZN(n2504) );
  NAND2_X1 U2900 ( .A1(n2294), .A2(n1938), .ZN(n2289) );
  NOR2_X1 U2901 ( .A1(n2561), .A2(n2197), .ZN(n3186) );
  OAI21_X1 U2902 ( .B1(n3000), .B2(n77), .A(n3185), .ZN(n3187) );
  AOI22_X1 U2903 ( .A1(n2997), .A2(\DataP/alu_out_M[12] ), .B1(n2992), .B2(
        \DataP/alu_out_W[12] ), .ZN(n3185) );
  NAND2_X1 U2904 ( .A1(n3005), .A2(\DataP/alu_out_W[12] ), .ZN(n3261) );
  AND2_X1 U2905 ( .A1(n1889), .A2(n2142), .ZN(n3400) );
  INV_X1 U2906 ( .A(\DataP/alu_a_in[10] ), .ZN(n3236) );
  NAND2_X1 U2907 ( .A1(n3232), .A2(n3656), .ZN(n3267) );
  NAND2_X1 U2908 ( .A1(n3658), .A2(n1921), .ZN(n3656) );
  NAND2_X1 U2909 ( .A1(n3220), .A2(n1922), .ZN(n3232) );
  INV_X1 U2910 ( .A(n1572), .ZN(n3254) );
  NOR2_X1 U2911 ( .A1(n2561), .A2(n2204), .ZN(n3189) );
  OAI21_X1 U2912 ( .B1(n1837), .B2(n81), .A(n3188), .ZN(n3190) );
  AOI22_X1 U2913 ( .A1(n2997), .A2(DRAM_ADDRESS[11]), .B1(n2992), .B2(
        \DataP/alu_out_W[11] ), .ZN(n3188) );
  INV_X1 U2914 ( .A(n3251), .ZN(n3250) );
  NAND2_X1 U2915 ( .A1(n3004), .A2(\DataP/alu_out_W[11] ), .ZN(n3244) );
  OR2_X1 U2916 ( .A1(n2566), .A2(n2164), .ZN(n3245) );
  AND4_X1 U2917 ( .A1(n3265), .A2(n2450), .A3(n3266), .A4(n3657), .ZN(n2319)
         );
  NOR2_X1 U2918 ( .A1(n2999), .A2(n93), .ZN(n3127) );
  OAI21_X1 U2919 ( .B1(n2561), .B2(n2220), .A(n3126), .ZN(n3128) );
  NAND2_X1 U2920 ( .A1(n3215), .A2(n2508), .ZN(n2509) );
  AND2_X1 U2921 ( .A1(\DataP/alu_b_in[8] ), .A2(n3510), .ZN(n2508) );
  NAND2_X1 U2922 ( .A1(n3219), .A2(\DataP/alu_a_in[9] ), .ZN(n3266) );
  NOR2_X1 U2923 ( .A1(n2562), .A2(n2190), .ZN(n3075) );
  OAI21_X1 U2924 ( .B1(n1837), .B2(n89), .A(n3074), .ZN(n3076) );
  INV_X1 U2925 ( .A(n3220), .ZN(n3219) );
  AND2_X1 U2926 ( .A1(\DataP/alu_b_in[9] ), .A2(n3510), .ZN(n2329) );
  NAND2_X1 U2927 ( .A1(n3218), .A2(n2545), .ZN(n2549) );
  NOR2_X1 U2928 ( .A1(n2561), .A2(n2211), .ZN(n3195) );
  OAI21_X1 U2929 ( .B1(n2999), .B2(n85), .A(n3192), .ZN(n3196) );
  AOI22_X1 U2930 ( .A1(n2997), .A2(DRAM_ADDRESS[10]), .B1(n2991), .B2(
        \DataP/alu_out_W[10] ), .ZN(n3192) );
  OR2_X1 U2931 ( .A1(n1846), .A2(n2334), .ZN(n2333) );
  INV_X1 U2932 ( .A(n2336), .ZN(n2334) );
  NAND2_X1 U2933 ( .A1(n2564), .A2(\DataP/ir_E[9] ), .ZN(n2391) );
  NOR2_X1 U2934 ( .A1(n2561), .A2(n2205), .ZN(n3078) );
  OAI21_X1 U2935 ( .B1(n3000), .B2(n97), .A(n3077), .ZN(n3079) );
  XNOR2_X1 U2936 ( .A(n3208), .B(\DataP/alu_b_in[7] ), .ZN(n3209) );
  INV_X1 U2937 ( .A(n3214), .ZN(\DataP/alu_b_in[7] ) );
  NAND2_X1 U2938 ( .A1(n3207), .A2(n1611), .ZN(n3208) );
  NAND2_X1 U2939 ( .A1(n3666), .A2(n3384), .ZN(n3211) );
  INV_X1 U2940 ( .A(\DataP/alu_a_in[6] ), .ZN(n3667) );
  NAND2_X1 U2941 ( .A1(n3206), .A2(n1920), .ZN(n3381) );
  INV_X1 U2942 ( .A(\DataP/alu_a_in[4] ), .ZN(n3204) );
  NAND2_X1 U2943 ( .A1(n2420), .A2(\DataP/alu_a_in[2] ), .ZN(n3370) );
  OR2_X1 U2944 ( .A1(n1996), .A2(n2337), .ZN(n3359) );
  OAI21_X1 U2945 ( .B1(n125), .B2(n3193), .A(n3112), .ZN(n3114) );
  NOR2_X1 U2946 ( .A1(n2560), .A2(n2214), .ZN(n3113) );
  NOR2_X1 U2947 ( .A1(n2561), .A2(n2215), .ZN(n3116) );
  AND2_X1 U2948 ( .A1(n3376), .A2(n3375), .ZN(n3205) );
  NOR2_X1 U2949 ( .A1(n2563), .A2(n2212), .ZN(n3109) );
  OAI21_X1 U2950 ( .B1(n1837), .B2(n113), .A(n3108), .ZN(n3110) );
  NOR2_X1 U2951 ( .A1(n2506), .A2(n2505), .ZN(n3203) );
  NOR2_X1 U2952 ( .A1(n1837), .A2(n109), .ZN(n3118) );
  OAI21_X1 U2953 ( .B1(n2562), .B2(n2221), .A(n3117), .ZN(n3119) );
  NAND2_X1 U2954 ( .A1(n1888), .A2(n3382), .ZN(n3212) );
  NOR2_X1 U2955 ( .A1(n2563), .A2(n2198), .ZN(n3121) );
  OAI21_X1 U2956 ( .B1(n3000), .B2(n105), .A(n3120), .ZN(n3122) );
  NAND2_X1 U2957 ( .A1(n3210), .A2(\DataP/alu_a_in[6] ), .ZN(n3384) );
  NOR2_X1 U2958 ( .A1(n1539), .A2(n2216), .ZN(n3124) );
  OAI21_X1 U2959 ( .B1(n3000), .B2(n101), .A(n3123), .ZN(n3125) );
  NOR2_X1 U2960 ( .A1(n3031), .A2(n3682), .ZN(n3068) );
  NAND4_X1 U2961 ( .A1(n520), .A2(n149), .A3(n145), .A4(n147), .ZN(n3682) );
  NAND2_X1 U2962 ( .A1(n3710), .A2(n3061), .ZN(n3067) );
  INV_X1 U2963 ( .A(n3073), .ZN(n3061) );
  XNOR2_X1 U2964 ( .A(n1871), .B(n2156), .ZN(n3058) );
  XNOR2_X1 U2965 ( .A(n529), .B(\DataP/Rs1[1] ), .ZN(n3054) );
  NOR2_X1 U2966 ( .A1(ALU_OPCODE_i[2]), .A2(n2134), .ZN(n3198) );
  XNOR2_X1 U2967 ( .A(n3207), .B(n1611), .ZN(n2522) );
  OR2_X1 U2968 ( .A1(n3002), .A2(n2182), .ZN(n2499) );
  AND2_X1 U2969 ( .A1(n3045), .A2(n3044), .ZN(n2314) );
  NOR2_X1 U2970 ( .A1(n3043), .A2(n3042), .ZN(n3044) );
  XNOR2_X1 U2971 ( .A(\DataP/Rs2[3] ), .B(n2570), .ZN(n3043) );
  NOR2_X1 U2972 ( .A1(n3041), .A2(n3040), .ZN(n3045) );
  XNOR2_X1 U2973 ( .A(\DataP/Rs2[1] ), .B(n529), .ZN(n3040) );
  OAI21_X1 U2974 ( .B1(n3018), .B2(n2479), .A(n2355), .ZN(n3050) );
  NAND4_X1 U2975 ( .A1(n1546), .A2(n1532), .A3(\DataP/opcode_W[4] ), .A4(n2159), .ZN(n2355) );
  XNOR2_X1 U2976 ( .A(\DataP/Rs2[2] ), .B(\DataP/add_D[2] ), .ZN(n3020) );
  XNOR2_X1 U2977 ( .A(\DataP/Rs2[4] ), .B(\DataP/add_D[4] ), .ZN(n3027) );
  INV_X1 U2978 ( .A(\DataP/alu_b_in[9] ), .ZN(n3218) );
  INV_X1 U2979 ( .A(n1537), .ZN(n2838) );
  AND3_X1 U2980 ( .A1(n1867), .A2(n3691), .A3(n3505), .ZN(n2138) );
  AND2_X1 U2981 ( .A1(n1948), .A2(n3689), .ZN(n2139) );
  NAND2_X1 U2982 ( .A1(n2181), .A2(n1995), .ZN(n3215) );
  XOR2_X1 U2983 ( .A(\DataP/dest_M[4] ), .B(n540), .Z(n2140) );
  NAND2_X1 U2984 ( .A1(n3067), .A2(n3066), .ZN(n3191) );
  INV_X1 U2985 ( .A(n2434), .ZN(n2349) );
  AND2_X1 U2986 ( .A1(n1897), .A2(n1898), .ZN(n2142) );
  AND2_X1 U2987 ( .A1(n3005), .A2(\DataP/alu_out_W[18] ), .ZN(n2145) );
  INV_X1 U2988 ( .A(n1880), .ZN(n3395) );
  OR2_X1 U2989 ( .A1(n3523), .A2(n1811), .ZN(n2147) );
  AND2_X1 U2990 ( .A1(n3347), .A2(n2433), .ZN(n2148) );
  AND2_X1 U2991 ( .A1(\DataP/alu_a_in[13] ), .A2(n2544), .ZN(n2149) );
  INV_X1 U2992 ( .A(n2407), .ZN(n2281) );
  INV_X1 U2993 ( .A(n2548), .ZN(n2546) );
  INV_X1 U2994 ( .A(n3353), .ZN(n3356) );
  OR2_X1 U2995 ( .A1(n3555), .A2(n3554), .ZN(n2158) );
  NAND2_X1 U2996 ( .A1(n2146), .A2(ALU_OPCODE_i[0]), .ZN(n3345) );
  INV_X1 U2997 ( .A(n3345), .ZN(n3223) );
  XOR2_X1 U2998 ( .A(\DataP/add_D[1] ), .B(n2160), .Z(n2163) );
  INV_X1 U2999 ( .A(n3660), .ZN(n3679) );
  AND2_X1 U3000 ( .A1(n1603), .A2(n3214), .ZN(n2181) );
  AND2_X1 U3001 ( .A1(\DataP/alu_b_in[19] ), .A2(n2545), .ZN(n2183) );
  AND2_X1 U3002 ( .A1(n3005), .A2(\DataP/alu_out_W[19] ), .ZN(n2184) );
  NAND2_X1 U3003 ( .A1(n3474), .A2(\DataP/alu_a_in[26] ), .ZN(n3505) );
  AND2_X1 U3004 ( .A1(n3580), .A2(n2011), .ZN(n2188) );
  INV_X1 U3005 ( .A(n3191), .ZN(n2994) );
  XNOR2_X1 U3006 ( .A(n3400), .B(n3395), .ZN(n3264) );
  NOR2_X1 U3007 ( .A1(n3910), .A2(n4020), .ZN(n2223) );
  XNOR2_X1 U3008 ( .A(\DataP/alu_a_in[11] ), .B(n3254), .ZN(n3318) );
  AND2_X1 U3009 ( .A1(n2550), .A2(n2428), .ZN(n2224) );
  AND2_X1 U3010 ( .A1(n2136), .A2(n1556), .ZN(n2235) );
  AND2_X1 U3011 ( .A1(n2130), .A2(n1948), .ZN(n2236) );
  AND3_X1 U3012 ( .A1(n2469), .A2(n2470), .A3(DRAM_ADDRESS[0]), .ZN(n2237) );
  AND3_X1 U3013 ( .A1(n2469), .A2(n2470), .A3(DRAM_ADDRESS[1]), .ZN(n2238) );
  AND2_X1 U3014 ( .A1(n1878), .A2(n3611), .ZN(n2239) );
  AND2_X1 U3015 ( .A1(\DataP/alu_a_in[4] ), .A2(n2461), .ZN(n2240) );
  INV_X1 U3016 ( .A(n2312), .ZN(n3496) );
  AND2_X1 U3017 ( .A1(\DataP/alu_a_in[17] ), .A2(n2538), .ZN(n2242) );
  NAND2_X1 U3018 ( .A1(n3272), .A2(n3271), .ZN(n2244) );
  INV_X1 U3019 ( .A(Rst), .ZN(n3012) );
  AOI22_X1 U3020 ( .A1(n2149), .A2(n2546), .B1(n2542), .B2(n2481), .ZN(n2282)
         );
  NAND2_X1 U3021 ( .A1(n3397), .A2(n2149), .ZN(n2283) );
  NAND2_X1 U3022 ( .A1(n3264), .A2(n2542), .ZN(n2284) );
  XNOR2_X1 U3023 ( .A(n2447), .B(n3396), .ZN(n3397) );
  NAND2_X1 U3024 ( .A1(n3272), .A2(n2285), .ZN(n3639) );
  AOI21_X1 U3025 ( .B1(n2287), .B2(n2294), .A(n2286), .ZN(n2285) );
  NAND2_X1 U3026 ( .A1(n2289), .A2(n3271), .ZN(n2286) );
  INV_X1 U3027 ( .A(n3264), .ZN(n2287) );
  NAND2_X1 U3028 ( .A1(n2290), .A2(n2225), .ZN(n2425) );
  NAND2_X1 U3029 ( .A1(n2291), .A2(n2370), .ZN(n3576) );
  NAND2_X1 U3030 ( .A1(n1992), .A2(n3510), .ZN(n2291) );
  XNOR2_X1 U3031 ( .A(n2293), .B(n2292), .ZN(n2577) );
  INV_X1 U3032 ( .A(n3442), .ZN(n2292) );
  NAND2_X1 U3033 ( .A1(n3437), .A2(n2235), .ZN(n2293) );
  AND2_X1 U3034 ( .A1(\DataP/alu_a_in[12] ), .A2(n2547), .ZN(n2294) );
  NAND2_X1 U3035 ( .A1(n2295), .A2(n3631), .ZN(n3412) );
  NAND2_X1 U3036 ( .A1(n3647), .A2(n3409), .ZN(n2295) );
  NAND2_X1 U3037 ( .A1(n2296), .A2(\DataP/alu_a_in[18] ), .ZN(n2304) );
  NAND2_X1 U3038 ( .A1(n2298), .A2(n2297), .ZN(n2296) );
  NAND2_X1 U3039 ( .A1(\DataP/alu_b_in[18] ), .A2(n2321), .ZN(n2297) );
  NAND2_X1 U3040 ( .A1(n3427), .A2(n3510), .ZN(n2298) );
  INV_X1 U3041 ( .A(n2000), .ZN(n2308) );
  AND2_X1 U3042 ( .A1(n2354), .A2(n2299), .ZN(n3612) );
  NOR2_X1 U3043 ( .A1(n3426), .A2(n1918), .ZN(n2301) );
  NAND2_X1 U3044 ( .A1(n3281), .A2(n1521), .ZN(n2302) );
  OAI22_X1 U3045 ( .A1(n2305), .A2(n2303), .B1(n1610), .B2(n2381), .ZN(n3459)
         );
  NAND4_X1 U3046 ( .A1(n2304), .A2(n3612), .A3(n1552), .A4(n3611), .ZN(n2303)
         );
  NAND4_X1 U3047 ( .A1(n3577), .A2(n2378), .A3(n3458), .A4(n1557), .ZN(n2305)
         );
  NOR2_X1 U3048 ( .A1(n2184), .A2(n2307), .ZN(n2306) );
  NAND2_X1 U3049 ( .A1(n2403), .A2(n2461), .ZN(n3669) );
  NAND2_X1 U3050 ( .A1(n2309), .A2(n3510), .ZN(n2403) );
  XNOR2_X1 U3051 ( .A(n3216), .B(\sra_131/SH[4] ), .ZN(n2309) );
  NAND2_X1 U3052 ( .A1(n1904), .A2(n2310), .ZN(n3070) );
  NOR2_X1 U3053 ( .A1(n2311), .A2(n3056), .ZN(n2310) );
  OR2_X1 U3054 ( .A1(n3054), .A2(n3055), .ZN(n2311) );
  NAND2_X1 U3055 ( .A1(n1839), .A2(\DataP/B_s[12] ), .ZN(n2387) );
  XNOR2_X1 U3056 ( .A(n2317), .B(n2316), .ZN(n3455) );
  INV_X1 U3057 ( .A(n3495), .ZN(n2316) );
  OAI21_X1 U3058 ( .B1(n3565), .B2(n1516), .A(n3463), .ZN(n2317) );
  NAND2_X1 U3059 ( .A1(n2318), .A2(n3460), .ZN(n3565) );
  NAND2_X1 U3060 ( .A1(n3592), .A2(n2188), .ZN(n2318) );
  NAND2_X1 U3061 ( .A1(n3269), .A2(n2319), .ZN(n2449) );
  NAND2_X1 U3062 ( .A1(n1866), .A2(\DataP/alu_a_in[7] ), .ZN(n3265) );
  NAND2_X1 U3063 ( .A1(n2322), .A2(n2320), .ZN(n3213) );
  NAND2_X1 U3064 ( .A1(n1950), .A2(n2321), .ZN(n2320) );
  INV_X1 U3065 ( .A(n3510), .ZN(n2321) );
  NAND2_X1 U3066 ( .A1(n3209), .A2(n3510), .ZN(n2322) );
  NAND4_X1 U3067 ( .A1(n2323), .A2(n2549), .A3(n2326), .A4(n2327), .ZN(n3220)
         );
  NAND2_X1 U3068 ( .A1(n2324), .A2(n2329), .ZN(n2323) );
  NAND2_X1 U3069 ( .A1(n3663), .A2(n2325), .ZN(n2324) );
  INV_X1 U3070 ( .A(n3216), .ZN(n2325) );
  NAND2_X1 U3071 ( .A1(n3215), .A2(n2329), .ZN(n2326) );
  NAND4_X1 U3072 ( .A1(n2510), .A2(n3218), .A3(n2328), .A4(n3663), .ZN(n2327)
         );
  NOR2_X1 U3073 ( .A1(n2543), .A2(n2003), .ZN(n2328) );
  INV_X1 U3074 ( .A(\DataP/alu_b_in[3] ), .ZN(n2330) );
  INV_X1 U3075 ( .A(n3002), .ZN(n2331) );
  NAND2_X1 U3076 ( .A1(n2564), .A2(\DataP/ir_E[8] ), .ZN(n2332) );
  NOR2_X1 U3077 ( .A1(\DataP/alu_b_in[10] ), .A2(n1572), .ZN(n3262) );
  NAND2_X1 U3078 ( .A1(n2331), .A2(DRAM_ADDRESS[10]), .ZN(n2335) );
  NAND2_X1 U3079 ( .A1(n2006), .A2(\DataP/alu_out_W[8] ), .ZN(n2336) );
  NAND2_X1 U3080 ( .A1(n2337), .A2(n1996), .ZN(n3358) );
  NAND2_X1 U3081 ( .A1(n2339), .A2(n2338), .ZN(n2337) );
  NAND2_X1 U3082 ( .A1(n1907), .A2(n3689), .ZN(n2338) );
  INV_X1 U3083 ( .A(n2148), .ZN(n2345) );
  OAI211_X1 U3084 ( .C1(n1984), .C2(n2348), .A(n2341), .B(n2340), .ZN(
        \DataP/PC_reg/N2 ) );
  NAND2_X1 U3085 ( .A1(n2148), .A2(n2347), .ZN(n2340) );
  AOI21_X1 U3086 ( .B1(n2431), .B2(n2347), .A(n2346), .ZN(n2341) );
  NAND3_X1 U3087 ( .A1(n2436), .A2(n2434), .A3(n443), .ZN(n2342) );
  NAND2_X1 U3088 ( .A1(n1919), .A2(n443), .ZN(n2348) );
  NAND2_X1 U3089 ( .A1(n3498), .A2(n2353), .ZN(n3499) );
  OAI21_X1 U3090 ( .B1(n2351), .B2(n2352), .A(n2350), .ZN(n3498) );
  INV_X1 U3091 ( .A(n3564), .ZN(n2350) );
  OAI21_X1 U3092 ( .B1(n3462), .B2(n3461), .A(n3460), .ZN(n2351) );
  NAND2_X1 U3093 ( .A1(n2462), .A2(n2242), .ZN(n2354) );
  NAND2_X1 U3094 ( .A1(n2358), .A2(n2321), .ZN(n2357) );
  INV_X1 U3095 ( .A(n1879), .ZN(n2358) );
  XNOR2_X1 U3096 ( .A(n3249), .B(n1879), .ZN(n3233) );
  INV_X1 U3097 ( .A(n2359), .ZN(n2550) );
  OAI211_X1 U3098 ( .C1(n3532), .C2(n2361), .A(n2360), .B(n3508), .ZN(n2359)
         );
  NAND2_X1 U3099 ( .A1(n2553), .A2(n3506), .ZN(n2360) );
  NAND2_X1 U3100 ( .A1(n3504), .A2(n3505), .ZN(n3532) );
  NAND2_X1 U3101 ( .A1(n3506), .A2(n3544), .ZN(n2361) );
  NAND2_X1 U3102 ( .A1(\DataP/alu_b_in[20] ), .A2(n2321), .ZN(n2364) );
  XNOR2_X1 U3103 ( .A(n3445), .B(\DataP/alu_b_in[20] ), .ZN(n2365) );
  INV_X1 U3104 ( .A(\DataP/alu_b_in[2] ), .ZN(n3011) );
  NAND2_X1 U3105 ( .A1(n3011), .A2(n3689), .ZN(n2366) );
  OR2_X1 U3106 ( .A1(n2503), .A2(n2467), .ZN(n2367) );
  OAI21_X1 U3107 ( .B1(n2467), .B2(n1550), .A(n3510), .ZN(n2368) );
  NAND2_X1 U3108 ( .A1(n3669), .A2(n3204), .ZN(n3377) );
  INV_X1 U3109 ( .A(n1638), .ZN(n2381) );
  NAND2_X1 U3110 ( .A1(n3442), .A2(n2383), .ZN(n2382) );
  INV_X1 U3111 ( .A(n3510), .ZN(n2383) );
  NAND2_X1 U3112 ( .A1(n1889), .A2(n1592), .ZN(n3249) );
  OR2_X1 U3113 ( .A1(n1988), .A2(n2394), .ZN(n2392) );
  INV_X1 U3114 ( .A(n2401), .ZN(n2394) );
  NAND3_X1 U3115 ( .A1(n2422), .A2(n1988), .A3(n2138), .ZN(n2395) );
  OAI22_X1 U3116 ( .A1(n300), .A2(n3911), .B1(n3910), .B2(n4018), .ZN(
        \DataP/PC_reg/N30 ) );
  NAND2_X1 U3117 ( .A1(n2424), .A2(n2523), .ZN(n3592) );
  NAND2_X1 U3118 ( .A1(n1528), .A2(n2240), .ZN(n3376) );
  OAI211_X1 U3119 ( .C1(n3488), .C2(n2406), .A(n2404), .B(n3510), .ZN(n2474)
         );
  NAND2_X1 U3120 ( .A1(n3488), .A2(n2405), .ZN(n2404) );
  XNOR2_X1 U3121 ( .A(n2497), .B(n2406), .ZN(n2405) );
  INV_X1 U3122 ( .A(\DataP/alu_b_in[27] ), .ZN(n2406) );
  NAND2_X1 U3123 ( .A1(n2474), .A2(n2445), .ZN(n2444) );
  NAND2_X1 U3124 ( .A1(n1934), .A2(n2383), .ZN(n2407) );
  NAND3_X1 U3125 ( .A1(n2503), .A2(n2133), .A3(n2241), .ZN(n2409) );
  NAND2_X1 U3126 ( .A1(n2408), .A2(n3510), .ZN(n2457) );
  XNOR2_X1 U3127 ( .A(n2409), .B(n1936), .ZN(n2408) );
  XNOR2_X1 U3128 ( .A(n1908), .B(n3511), .ZN(n2413) );
  NAND2_X1 U3129 ( .A1(n2410), .A2(n2411), .ZN(\DataP/PC_reg/N32 ) );
  NAND2_X1 U3130 ( .A1(n2413), .A2(n2412), .ZN(n2410) );
  NAND3_X1 U3131 ( .A1(n3466), .A2(n2131), .A3(n3467), .ZN(n2422) );
  AOI21_X1 U3132 ( .B1(n2551), .B2(n2224), .A(n2427), .ZN(n3685) );
  NAND2_X1 U3133 ( .A1(n1906), .A2(n2552), .ZN(n2551) );
  OAI21_X1 U3134 ( .B1(n2144), .B2(n2432), .A(n3351), .ZN(n2431) );
  AOI22_X1 U3135 ( .A1(n3342), .A2(n1876), .B1(n3343), .B2(n3356), .ZN(n2432)
         );
  NOR2_X1 U3136 ( .A1(n3356), .A2(n2132), .ZN(n2433) );
  NOR2_X1 U3137 ( .A1(n3357), .A2(n2435), .ZN(n2434) );
  AND2_X1 U3138 ( .A1(\DataP/ALU_C/shifter/N82 ), .A2(n3675), .ZN(n2435) );
  AOI21_X1 U3139 ( .B1(n3354), .B2(n2438), .A(n2437), .ZN(n2436) );
  NOR2_X1 U3140 ( .A1(n3356), .A2(n3355), .ZN(n2437) );
  NOR2_X1 U3141 ( .A1(ALU_OPCODE_i[2]), .A2(n2146), .ZN(n2438) );
  NOR2_X1 U3142 ( .A1(n2440), .A2(n2439), .ZN(n2441) );
  XNOR2_X1 U3143 ( .A(n3426), .B(n1928), .ZN(n3427) );
  NAND2_X1 U3144 ( .A1(n2441), .A2(n1598), .ZN(n3426) );
  OAI211_X1 U3145 ( .C1(n2474), .C2(\DataP/alu_a_in[27] ), .A(n2444), .B(n2443), .ZN(n3506) );
  NAND2_X1 U3146 ( .A1(n1912), .A2(n2446), .ZN(n2443) );
  NOR2_X1 U3147 ( .A1(n1912), .A2(n2446), .ZN(n2445) );
  INV_X1 U3148 ( .A(n2473), .ZN(n2446) );
  NAND4_X1 U3149 ( .A1(n2142), .A2(n2504), .A3(n1995), .A4(n3395), .ZN(n2447)
         );
  NAND2_X1 U3150 ( .A1(n2455), .A2(n2450), .ZN(n2448) );
  NAND2_X1 U3151 ( .A1(n2452), .A2(n2478), .ZN(n2451) );
  INV_X1 U3152 ( .A(n3318), .ZN(n2452) );
  NAND2_X1 U3153 ( .A1(n3250), .A2(n2454), .ZN(n2453) );
  AND2_X1 U3154 ( .A1(n1863), .A2(n3510), .ZN(n2454) );
  NAND2_X1 U3155 ( .A1(n2456), .A2(n3268), .ZN(n2455) );
  NAND2_X1 U3156 ( .A1(n3267), .A2(n3266), .ZN(n2456) );
  NAND2_X1 U3157 ( .A1(n2457), .A2(n2502), .ZN(n3474) );
  NAND2_X1 U3158 ( .A1(n2459), .A2(n2458), .ZN(n3206) );
  AOI21_X1 U3159 ( .B1(n2460), .B2(n2236), .A(n2139), .ZN(n2458) );
  NAND2_X1 U3160 ( .A1(n1574), .A2(n2460), .ZN(n2459) );
  AOI21_X1 U3161 ( .B1(n2003), .B2(n1948), .A(n2375), .ZN(n2460) );
  NAND2_X1 U3162 ( .A1(n3072), .A2(n3073), .ZN(n2470) );
  AOI21_X1 U3163 ( .B1(n2993), .B2(\DataP/alu_out_W[0] ), .A(n2237), .ZN(n3112) );
  NOR2_X1 U3164 ( .A1(n2464), .A2(n1938), .ZN(n2463) );
  INV_X1 U3165 ( .A(n2493), .ZN(n2464) );
  AND2_X1 U3166 ( .A1(\DataP/alu_a_in[16] ), .A2(n2466), .ZN(n2465) );
  OR2_X1 U3167 ( .A1(\DataP/alu_b_in[16] ), .A2(n3510), .ZN(n2466) );
  AND2_X1 U3168 ( .A1(n3470), .A2(\DataP/alu_a_in[25] ), .ZN(n3544) );
  INV_X1 U3169 ( .A(\DataP/alu_b_in[25] ), .ZN(n2467) );
  INV_X1 U3170 ( .A(Rst), .ZN(n2468) );
  AOI21_X1 U3171 ( .B1(n2993), .B2(\DataP/alu_out_W[1] ), .A(n2238), .ZN(n3115) );
  NAND2_X1 U3172 ( .A1(\DataP/alu_b_in[27] ), .A2(n2478), .ZN(n2473) );
  XNOR2_X1 U3173 ( .A(n2568), .B(n523), .ZN(n2476) );
  AND2_X1 U3174 ( .A1(n3059), .A2(n3057), .ZN(n2477) );
  NOR2_X1 U3175 ( .A1(n1581), .A2(\DataP/alu_b_in[2] ), .ZN(n2501) );
  INV_X1 U3176 ( .A(n3510), .ZN(n2478) );
  NAND2_X1 U3177 ( .A1(n2571), .A2(n2162), .ZN(n2479) );
  NAND4_X1 U3178 ( .A1(n2480), .A2(n2186), .A3(n3023), .A4(n2140), .ZN(n3063)
         );
  INV_X1 U3179 ( .A(n2547), .ZN(n2481) );
  OR2_X1 U3180 ( .A1(n3206), .A2(n1920), .ZN(n3382) );
  NAND4_X1 U3181 ( .A1(n1889), .A2(n2142), .A3(n2390), .A4(n2482), .ZN(n2483)
         );
  NAND3_X1 U3182 ( .A1(n2485), .A2(n2484), .A3(n2483), .ZN(n3392) );
  OR2_X1 U3183 ( .A1(n1889), .A2(n3417), .ZN(n2484) );
  NAND2_X1 U3184 ( .A1(n2486), .A2(\DataP/alu_b_in[15] ), .ZN(n2485) );
  NAND2_X1 U3185 ( .A1(n2142), .A2(n2487), .ZN(n2486) );
  OR2_X1 U3186 ( .A1(n1563), .A2(\DataP/alu_b_in[17] ), .ZN(n2488) );
  NAND2_X1 U3187 ( .A1(\DataP/alu_b_in[16] ), .A2(n3424), .ZN(n2493) );
  NAND2_X1 U3188 ( .A1(n3437), .A2(n2495), .ZN(n2494) );
  NOR2_X1 U3189 ( .A1(\DataP/alu_b_in[16] ), .A2(n1580), .ZN(n2495) );
  NAND2_X1 U3190 ( .A1(n2564), .A2(\DataP/ir_E[6] ), .ZN(n2500) );
  NAND3_X1 U3191 ( .A1(n1598), .A2(n2136), .A3(n3421), .ZN(n3445) );
  OAI21_X1 U3192 ( .B1(n2522), .B2(n3689), .A(n2521), .ZN(n3210) );
  NAND2_X1 U3193 ( .A1(n3384), .A2(n3385), .ZN(n3666) );
  OR2_X1 U3194 ( .A1(n3210), .A2(\DataP/alu_a_in[6] ), .ZN(n3385) );
  NAND3_X1 U3195 ( .A1(n3087), .A2(n3090), .A3(n3089), .ZN(n2505) );
  NAND3_X1 U3196 ( .A1(n2511), .A2(n2510), .A3(n3510), .ZN(n2507) );
  INV_X1 U3197 ( .A(n3215), .ZN(n2510) );
  NOR2_X1 U3198 ( .A1(n2003), .A2(\DataP/alu_b_in[8] ), .ZN(n2511) );
  NAND2_X1 U3199 ( .A1(n3425), .A2(n2478), .ZN(n2512) );
  NAND2_X1 U3200 ( .A1(\DataP/alu_b_in[6] ), .A2(n3689), .ZN(n2521) );
  NOR2_X1 U3201 ( .A1(n2529), .A2(n2528), .ZN(n297) );
  NOR2_X1 U3202 ( .A1(n1609), .A2(n1909), .ZN(n2528) );
  NAND2_X1 U3203 ( .A1(n2530), .A2(n1990), .ZN(n2529) );
  NAND2_X1 U3204 ( .A1(n3708), .A2(n2153), .ZN(n2530) );
  OAI211_X1 U3205 ( .C1(n1991), .C2(n2533), .A(n2531), .B(n2537), .ZN(
        \DataP/PC_reg/N33 ) );
  NAND2_X1 U3206 ( .A1(n1909), .A2(n2532), .ZN(n2531) );
  NOR2_X1 U3207 ( .A1(n2534), .A2(n3911), .ZN(n2532) );
  NAND2_X1 U3208 ( .A1(n2536), .A2(n1919), .ZN(n2533) );
  NOR2_X1 U3209 ( .A1(n2535), .A2(n2153), .ZN(n2534) );
  INV_X1 U3210 ( .A(n3707), .ZN(n2535) );
  NAND2_X1 U3211 ( .A1(n1990), .A2(n1609), .ZN(n2536) );
  OR2_X1 U3212 ( .A1(n3910), .A2(n4023), .ZN(n2537) );
  AND2_X1 U3213 ( .A1(\DataP/ALU_C/shifter/N48 ), .A2(n3007), .ZN(n2539) );
  NAND2_X1 U3214 ( .A1(n3395), .A2(n2545), .ZN(n2547) );
  NAND2_X1 U3215 ( .A1(n1860), .A2(n2543), .ZN(n2548) );
  INV_X1 U3216 ( .A(n3505), .ZN(n2553) );
  INV_X1 U3217 ( .A(n3543), .ZN(n2556) );
  OAI211_X1 U3218 ( .C1(n1841), .C2(n3697), .A(\DataP/alu_b_in[15] ), .B(n3660), .ZN(n3403) );
  NAND2_X1 U3219 ( .A1(n2564), .A2(\DataP/ir_E[7] ), .ZN(n3082) );
  NAND2_X1 U3220 ( .A1(n1905), .A2(\DataP/IMM_s[19] ), .ZN(n3290) );
  XNOR2_X1 U3221 ( .A(\DataP/alu_a_in[3] ), .B(n1963), .ZN(n3681) );
  OAI21_X1 U3222 ( .B1(\DataP/alu_a_in[13] ), .B2(n1860), .A(n3697), .ZN(n3650) );
  XNOR2_X1 U3223 ( .A(\DataP/alu_a_in[13] ), .B(n1860), .ZN(n3651) );
  INV_X1 U3224 ( .A(\DataP/alu_b_in[13] ), .ZN(n3396) );
  AOI22_X1 U3225 ( .A1(n2996), .A2(\DataP/alu_out_M[30] ), .B1(n2992), .B2(
        \DataP/alu_out_W[30] ), .ZN(n3132) );
  AOI22_X1 U3226 ( .A1(n2996), .A2(DRAM_ADDRESS[7]), .B1(n2991), .B2(
        \DataP/alu_out_W[7] ), .ZN(n3077) );
  AOI22_X1 U3227 ( .A1(n2996), .A2(\DataP/alu_out_M[31] ), .B1(n2992), .B2(
        \DataP/alu_out_W[31] ), .ZN(n3129) );
  AOI22_X1 U3228 ( .A1(n2995), .A2(DRAM_ADDRESS[9]), .B1(n2992), .B2(
        \DataP/alu_out_W[9] ), .ZN(n3074) );
  AOI22_X1 U3229 ( .A1(n2996), .A2(DRAM_ADDRESS[5]), .B1(n2991), .B2(
        \DataP/alu_out_W[5] ), .ZN(n3120) );
  AOI22_X1 U3230 ( .A1(n2996), .A2(DRAM_ADDRESS[6]), .B1(n2991), .B2(
        \DataP/alu_out_W[6] ), .ZN(n3123) );
  AOI22_X1 U3231 ( .A1(n2995), .A2(DRAM_ADDRESS[4]), .B1(n2991), .B2(
        \DataP/alu_out_W[4] ), .ZN(n3117) );
  AOI22_X1 U3232 ( .A1(n2995), .A2(DRAM_ADDRESS[3]), .B1(n2992), .B2(
        \DataP/alu_out_W[3] ), .ZN(n3108) );
  AOI22_X1 U3233 ( .A1(n2996), .A2(DRAM_ADDRESS[8]), .B1(n2991), .B2(
        \DataP/alu_out_W[8] ), .ZN(n3126) );
  AOI22_X1 U3234 ( .A1(n2995), .A2(DRAM_ADDRESS[2]), .B1(n2993), .B2(
        \DataP/alu_out_W[2] ), .ZN(n3111) );
  NAND3_X1 U3235 ( .A1(n1568), .A2(n432), .A3(n2998), .ZN(n2560) );
  NAND2_X1 U3236 ( .A1(n2006), .A2(\DataP/alu_out_W[2] ), .ZN(n3096) );
  NAND2_X1 U3237 ( .A1(n2006), .A2(\DataP/alu_out_W[9] ), .ZN(n3047) );
  NAND2_X1 U3238 ( .A1(n2006), .A2(\DataP/alu_out_W[4] ), .ZN(n3100) );
  NAND2_X1 U3239 ( .A1(n2006), .A2(\DataP/alu_out_W[7] ), .ZN(n3080) );
  NAND2_X1 U3240 ( .A1(n3330), .A2(\DataP/alu_out_W[0] ), .ZN(n3088) );
  NAND2_X1 U3241 ( .A1(n2006), .A2(\DataP/alu_out_W[3] ), .ZN(n3092) );
  NAND2_X1 U3242 ( .A1(n3330), .A2(\DataP/alu_out_W[1] ), .ZN(n3084) );
  NAND2_X1 U3243 ( .A1(n3327), .A2(\DataP/B_s[11] ), .ZN(n3247) );
  NAND2_X1 U3244 ( .A1(n1518), .A2(\DataP/B_s[2] ), .ZN(n3099) );
  NAND2_X1 U3245 ( .A1(n1839), .A2(\DataP/B_s[10] ), .ZN(n3231) );
  NAND2_X1 U3246 ( .A1(n1635), .A2(\DataP/B_s[4] ), .ZN(n3103) );
  NAND2_X1 U3247 ( .A1(n1518), .A2(\DataP/B_s[7] ), .ZN(n3083) );
  NAND2_X1 U3248 ( .A1(n1518), .A2(\DataP/B_s[0] ), .ZN(n3091) );
  NAND2_X1 U3249 ( .A1(n1518), .A2(\DataP/B_s[3] ), .ZN(n3095) );
  NAND2_X1 U3250 ( .A1(n1635), .A2(\DataP/B_s[5] ), .ZN(n3107) );
  XNOR2_X1 U3251 ( .A(n536), .B(n2154), .ZN(n3059) );
  INV_X1 U3252 ( .A(n2005), .ZN(n2566) );
  NAND2_X1 U3253 ( .A1(n2011), .A2(n3576), .ZN(n3582) );
  NAND2_X1 U3254 ( .A1(n3593), .A2(n2011), .ZN(n3461) );
  NAND2_X1 U3255 ( .A1(n3443), .A2(n2011), .ZN(n3460) );
  XNOR2_X1 U3256 ( .A(n1999), .B(\DataP/Rs1[2] ), .ZN(n3055) );
  XNOR2_X1 U3257 ( .A(\DataP/Rs2[2] ), .B(n1999), .ZN(n3042) );
  XNOR2_X1 U3258 ( .A(n530), .B(n538), .ZN(n3022) );
  NOR2_X1 U3259 ( .A1(\DataP/dest_M[4] ), .A2(\DataP/dest_M[3] ), .ZN(n3037)
         );
  INV_X1 U3260 ( .A(n2574), .ZN(n2575) );
  XNOR2_X1 U3261 ( .A(n528), .B(n2154), .ZN(n3053) );
  XNOR2_X1 U3262 ( .A(n528), .B(\DataP/Rs2[0] ), .ZN(n3041) );
  XNOR2_X1 U3263 ( .A(n528), .B(n536), .ZN(n3021) );
  XNOR2_X1 U3264 ( .A(n540), .B(n524), .ZN(n3057) );
  NAND2_X1 U3265 ( .A1(n3034), .A2(n2161), .ZN(n3035) );
  XNOR2_X1 U3266 ( .A(n1987), .B(n2572), .ZN(n3609) );
  XNOR2_X1 U3267 ( .A(\DataP/add_D[1] ), .B(\DataP/Rs2[1] ), .ZN(n3019) );
  XNOR2_X1 U3268 ( .A(\DataP/dest_M[1] ), .B(\DataP/add_D[1] ), .ZN(n3023) );
  XNOR2_X1 U3269 ( .A(\DataP/opcode_W[2] ), .B(n2151), .ZN(n3018) );
  XNOR2_X1 U3270 ( .A(n3428), .B(n1559), .ZN(n3436) );
  NAND2_X1 U3271 ( .A1(n521), .A2(n520), .ZN(n3060) );
  OAI21_X1 U3272 ( .B1(n1948), .B2(n3671), .A(n3694), .ZN(n3379) );
  XNOR2_X1 U3273 ( .A(\DataP/alu_a_in[5] ), .B(\lt_x_134/B[5] ), .ZN(n3380) );
  NAND2_X1 U3274 ( .A1(n1518), .A2(\DataP/B_s[1] ), .ZN(n3087) );
  XNOR2_X1 U3275 ( .A(n2568), .B(\DataP/Rs2[3] ), .ZN(n3024) );
  NAND4_X1 U3276 ( .A1(n1862), .A2(n1871), .A3(n540), .A4(n2568), .ZN(n3026)
         );
  OAI21_X1 U3277 ( .B1(n2575), .B2(n3682), .A(Rst), .ZN(
        \DataP/FORWARDING_BR/N12 ) );
  NAND2_X1 U3278 ( .A1(n1850), .A2(n3502), .ZN(n3545) );
  INV_X1 U3279 ( .A(n3445), .ZN(n3438) );
  OAI211_X1 U3280 ( .C1(\DataP/opcode_M[4] ), .C2(\DataP/opcode_M[0] ), .A(
        \DataP/opcode_M[1] ), .B(n1895), .ZN(n3034) );
  OAI22_X1 U3281 ( .A1(n1996), .A2(n3362), .B1(n1916), .B2(n3694), .ZN(n3363)
         );
  XNOR2_X1 U3282 ( .A(\DataP/alu_a_in[1] ), .B(n1916), .ZN(n3364) );
  NAND2_X1 U3283 ( .A1(n3069), .A2(n3068), .ZN(n3072) );
  OR2_X1 U3284 ( .A1(n3069), .A2(n3065), .ZN(n3066) );
  AOI21_X1 U3285 ( .B1(n3498), .B2(n3496), .A(n3495), .ZN(n3466) );
  AOI21_X1 U3286 ( .B1(\sra_131/SH[1] ), .B2(n3693), .A(n3697), .ZN(n3362) );
  NAND2_X1 U3287 ( .A1(n2564), .A2(\DataP/ir_E[11] ), .ZN(n3246) );
  NAND2_X1 U3288 ( .A1(n2565), .A2(\DataP/ir_E[10] ), .ZN(n3230) );
  OR2_X1 U3289 ( .A1(n2228), .A2(n3002), .ZN(n3048) );
  NAND2_X1 U3290 ( .A1(n2564), .A2(\DataP/ir_E[4] ), .ZN(n3102) );
  OR2_X1 U3291 ( .A1(n3002), .A2(n2230), .ZN(n3081) );
  NAND2_X1 U3292 ( .A1(n2564), .A2(\DataP/ir_E[2] ), .ZN(n3098) );
  NAND2_X1 U3293 ( .A1(n2564), .A2(\DataP/ir_E[3] ), .ZN(n3094) );
  NAND2_X1 U3294 ( .A1(n3328), .A2(\DataP/ir_E[5] ), .ZN(n3106) );
  NAND2_X1 U3295 ( .A1(n3328), .A2(\DataP/ir_E[0] ), .ZN(n3090) );
  NAND2_X1 U3296 ( .A1(n3328), .A2(\DataP/ir_E[1] ), .ZN(n3086) );
  NAND4_X1 U3297 ( .A1(n2711), .A2(n1913), .A3(n1916), .A4(n1605), .ZN(n2642)
         );
  NOR2_X1 U3298 ( .A1(n2846), .A2(n2642), .ZN(n2602) );
  NAND2_X1 U3299 ( .A1(n1605), .A2(n2711), .ZN(n2578) );
  AOI22_X1 U3300 ( .A1(n2709), .A2(\DataP/alu_a_in[1] ), .B1(
        \DataP/alu_a_in[2] ), .B2(n2711), .ZN(n2580) );
  AOI22_X1 U3301 ( .A1(n2839), .A2(n2578), .B1(n2580), .B2(n2988), .ZN(n2591)
         );
  NAND2_X1 U3302 ( .A1(n1913), .A2(n2591), .ZN(n2612) );
  AOI22_X1 U3303 ( .A1(n2709), .A2(\DataP/alu_a_in[3] ), .B1(
        \DataP/alu_a_in[4] ), .B2(n2711), .ZN(n2579) );
  AOI22_X1 U3304 ( .A1(n2709), .A2(\DataP/alu_a_in[5] ), .B1(
        \DataP/alu_a_in[6] ), .B2(n2711), .ZN(n2582) );
  AOI22_X1 U3305 ( .A1(n2713), .A2(n2579), .B1(n2582), .B2(n1916), .ZN(n2590)
         );
  AOI22_X1 U3306 ( .A1(n2709), .A2(\DataP/alu_a_in[7] ), .B1(
        \DataP/alu_a_in[8] ), .B2(n2711), .ZN(n2581) );
  AOI22_X1 U3307 ( .A1(n2709), .A2(\DataP/alu_a_in[9] ), .B1(
        \DataP/alu_a_in[10] ), .B2(n2711), .ZN(n2583) );
  AOI22_X1 U3308 ( .A1(n2713), .A2(n2581), .B1(n2583), .B2(n2988), .ZN(n2593)
         );
  AOI22_X1 U3309 ( .A1(n2842), .A2(n2590), .B1(n2593), .B2(n1913), .ZN(n2611)
         );
  AOI22_X1 U3310 ( .A1(n1915), .A2(n2612), .B1(n2611), .B2(n2064), .ZN(n2654)
         );
  NOR2_X1 U3311 ( .A1(\lt_x_135/B[4] ), .A2(n2697), .ZN(
        \DataP/ALU_C/shifter/N28 ) );
  AOI22_X1 U3312 ( .A1(n2709), .A2(n1605), .B1(\DataP/alu_a_in[1] ), .B2(n2711), .ZN(n2584) );
  AOI22_X1 U3313 ( .A1(n2709), .A2(\DataP/alu_a_in[2] ), .B1(
        \DataP/alu_a_in[3] ), .B2(n2710), .ZN(n2586) );
  AOI22_X1 U3314 ( .A1(n2713), .A2(n2584), .B1(n2586), .B2(n1916), .ZN(n2595)
         );
  NAND2_X1 U3315 ( .A1(n1913), .A2(n2595), .ZN(n2616) );
  INV_X1 U3316 ( .A(n1907), .ZN(n2713) );
  NAND2_X1 U3317 ( .A1(n1930), .A2(n2763), .ZN(n2780) );
  NOR2_X1 U3318 ( .A1(n1915), .A2(n2780), .ZN(n2792) );
  MUX2_X1 U3319 ( .A(n2748), .B(n2792), .S(\lt_x_134/B[4] ), .Z(
        \DataP/ALU_C/shifter/N63 ) );
  NAND3_X1 U3320 ( .A1(n2781), .A2(n2845), .A3(n2844), .ZN(n2801) );
  AOI22_X1 U3321 ( .A1(n2842), .A2(n2750), .B1(n2749), .B2(n1930), .ZN(n2782)
         );
  AOI22_X1 U3322 ( .A1(n2842), .A2(n2752), .B1(n2751), .B2(n1930), .ZN(n2823)
         );
  AOI22_X1 U3323 ( .A1(n1915), .A2(n2782), .B1(n2823), .B2(n2845), .ZN(n2753)
         );
  NAND2_X1 U3324 ( .A1(n2847), .A2(n2753), .ZN(n2754) );
  OAI21_X1 U3325 ( .B1(n2065), .B2(n2801), .A(n2754), .ZN(
        \DataP/ALU_C/shifter/N64 ) );
  NAND3_X1 U3326 ( .A1(n2784), .A2(n2127), .A3(n2844), .ZN(n2802) );
  AOI22_X1 U3327 ( .A1(n2842), .A2(n2756), .B1(n2755), .B2(n1930), .ZN(n2785)
         );
  AOI22_X1 U3328 ( .A1(n2842), .A2(n2758), .B1(n2757), .B2(n1930), .ZN(n2827)
         );
  AOI22_X1 U3329 ( .A1(n2846), .A2(n2785), .B1(n2827), .B2(n2064), .ZN(n2759)
         );
  NAND2_X1 U3330 ( .A1(n2065), .A2(n2759), .ZN(n2760) );
  OAI21_X1 U3331 ( .B1(n2065), .B2(n2802), .A(n2760), .ZN(
        \DataP/ALU_C/shifter/N65 ) );
  AND2_X1 U3332 ( .A1(n2065), .A2(n2761), .ZN(\DataP/ALU_C/shifter/N66 ) );
  AOI22_X1 U3333 ( .A1(n2842), .A2(n2763), .B1(n2762), .B2(n1930), .ZN(n2788)
         );
  AOI22_X1 U3334 ( .A1(n2842), .A2(n2765), .B1(n2764), .B2(n1930), .ZN(n2835)
         );
  AOI22_X1 U3335 ( .A1(n2846), .A2(n2788), .B1(n2835), .B2(n2127), .ZN(n2774)
         );
  AND2_X1 U3336 ( .A1(n2847), .A2(n2774), .ZN(\DataP/ALU_C/shifter/N67 ) );
  AOI22_X1 U3337 ( .A1(n2846), .A2(n2767), .B1(n2766), .B2(n2064), .ZN(n2800)
         );
  AND2_X1 U3338 ( .A1(n2847), .A2(n2800), .ZN(\DataP/ALU_C/shifter/N68 ) );
  AOI22_X1 U3339 ( .A1(n2846), .A2(n2769), .B1(n2768), .B2(n2845), .ZN(n2808)
         );
  AND2_X1 U3340 ( .A1(n2847), .A2(n2808), .ZN(\DataP/ALU_C/shifter/N69 ) );
  AOI22_X1 U3341 ( .A1(n1914), .A2(\DataP/alu_a_in[10] ), .B1(
        \DataP/alu_a_in[9] ), .B2(n1931), .ZN(n2804) );
  AOI22_X1 U3342 ( .A1(\sra_131/SH[1] ), .A2(n2770), .B1(n2804), .B2(n1916), 
        .ZN(n2816) );
  AOI22_X1 U3343 ( .A1(n2842), .A2(n2771), .B1(n2816), .B2(n1930), .ZN(n2834)
         );
  AOI22_X1 U3344 ( .A1(n1914), .A2(\DataP/alu_a_in[8] ), .B1(
        \DataP/alu_a_in[7] ), .B2(n1931), .ZN(n2803) );
  AOI22_X1 U3345 ( .A1(n1914), .A2(\DataP/alu_a_in[6] ), .B1(
        \DataP/alu_a_in[5] ), .B2(n1931), .ZN(n2806) );
  AOI22_X1 U3346 ( .A1(\sra_131/SH[1] ), .A2(n2803), .B1(n2806), .B2(n1916), 
        .ZN(n2815) );
  AOI22_X1 U3347 ( .A1(n1914), .A2(\DataP/alu_a_in[4] ), .B1(
        \DataP/alu_a_in[3] ), .B2(n1931), .ZN(n2805) );
  AOI22_X1 U3348 ( .A1(n2842), .A2(n2815), .B1(n2772), .B2(n1930), .ZN(n2773)
         );
  AOI22_X1 U3349 ( .A1(n2846), .A2(n2834), .B1(n2773), .B2(n2845), .ZN(n2775)
         );
  MUX2_X1 U3350 ( .A(n2775), .B(n2774), .S(\lt_x_134/B[4] ), .Z(
        \DataP/ALU_C/shifter/N51 ) );
  NAND2_X1 U3351 ( .A1(n1930), .A2(n2776), .ZN(n2778) );
  AOI22_X1 U3352 ( .A1(n2846), .A2(n2778), .B1(n2777), .B2(n2064), .ZN(n2813)
         );
  AND2_X1 U3353 ( .A1(n2065), .A2(n2813), .ZN(\DataP/ALU_C/shifter/N70 ) );
  AOI22_X1 U3354 ( .A1(n2846), .A2(n2780), .B1(n2779), .B2(n2064), .ZN(n2819)
         );
  AND2_X1 U3355 ( .A1(n2065), .A2(n2819), .ZN(\DataP/ALU_C/shifter/N71 ) );
  NAND2_X1 U3356 ( .A1(n2781), .A2(n2844), .ZN(n2783) );
  AOI22_X1 U3357 ( .A1(n2846), .A2(n2783), .B1(n2782), .B2(n2127), .ZN(n2824)
         );
  AND2_X1 U3358 ( .A1(n2065), .A2(n2824), .ZN(\DataP/ALU_C/shifter/N72 ) );
  NAND2_X1 U3359 ( .A1(n2784), .A2(n2844), .ZN(n2786) );
  AOI22_X1 U3360 ( .A1(n2846), .A2(n2786), .B1(n2785), .B2(n2127), .ZN(n2828)
         );
  AND2_X1 U3361 ( .A1(n2847), .A2(n2828), .ZN(\DataP/ALU_C/shifter/N73 ) );
  NOR2_X1 U3362 ( .A1(n1915), .A2(n2787), .ZN(n2832) );
  AND2_X1 U3363 ( .A1(n2832), .A2(n2847), .ZN(\DataP/ALU_C/shifter/N74 ) );
  NOR2_X1 U3364 ( .A1(n1915), .A2(n2788), .ZN(n2836) );
  INV_X1 U3365 ( .A(n2126), .ZN(n2840) );
  AOI22_X1 U3366 ( .A1(n2713), .A2(n2853), .B1(n2856), .B2(n2126), .ZN(n2867)
         );
  AOI22_X1 U3367 ( .A1(n2841), .A2(n2865), .B1(n2867), .B2(n1913), .ZN(n2918)
         );
  AOI22_X1 U3368 ( .A1(n2986), .A2(\DataP/alu_a_in[23] ), .B1(
        \DataP/alu_a_in[22] ), .B2(n2985), .ZN(n2855) );
  AOI22_X1 U3369 ( .A1(n2986), .A2(\DataP/alu_a_in[19] ), .B1(
        \DataP/alu_a_in[18] ), .B2(n2985), .ZN(n2857) );
  AOI22_X1 U3370 ( .A1(n2709), .A2(\DataP/alu_a_in[17] ), .B1(
        \DataP/alu_a_in[16] ), .B2(n2985), .ZN(n2860) );
  AOI22_X1 U3371 ( .A1(n2841), .A2(n2866), .B1(n2869), .B2(n1930), .ZN(n2976)
         );
  AOI22_X1 U3372 ( .A1(n1915), .A2(n2918), .B1(n2976), .B2(n2127), .ZN(n2893)
         );
  AOI22_X1 U3373 ( .A1(n2709), .A2(n1841), .B1(\DataP/alu_a_in[14] ), .B2(
        n2710), .ZN(n2859) );
  AOI22_X1 U3374 ( .A1(n2709), .A2(\DataP/alu_a_in[13] ), .B1(
        \DataP/alu_a_in[12] ), .B2(n2985), .ZN(n2862) );
  AOI22_X1 U3375 ( .A1(n2713), .A2(n2859), .B1(n2862), .B2(n2988), .ZN(n2868)
         );
  AOI22_X1 U3376 ( .A1(n2709), .A2(\DataP/alu_a_in[11] ), .B1(
        \DataP/alu_a_in[10] ), .B2(n2711), .ZN(n2861) );
  AOI22_X1 U3377 ( .A1(n2709), .A2(\DataP/alu_a_in[9] ), .B1(
        \DataP/alu_a_in[8] ), .B2(n2985), .ZN(n2932) );
  AOI22_X1 U3378 ( .A1(n2713), .A2(n2861), .B1(n2932), .B2(n2988), .ZN(n2951)
         );
  AOI22_X1 U3379 ( .A1(n2841), .A2(n2868), .B1(n2951), .B2(n1913), .ZN(n2975)
         );
  AOI22_X1 U3380 ( .A1(n2709), .A2(\DataP/alu_a_in[7] ), .B1(
        \DataP/alu_a_in[6] ), .B2(n2985), .ZN(n2931) );
  AOI22_X1 U3381 ( .A1(n2709), .A2(\DataP/alu_a_in[5] ), .B1(
        \DataP/alu_a_in[4] ), .B2(n2710), .ZN(n2934) );
  AOI22_X1 U3382 ( .A1(n2840), .A2(n2931), .B1(n2934), .B2(n2988), .ZN(n2950)
         );
  AOI22_X1 U3383 ( .A1(n2709), .A2(\DataP/alu_a_in[3] ), .B1(
        \DataP/alu_a_in[2] ), .B2(n2711), .ZN(n2933) );
  AOI22_X1 U3384 ( .A1(n2987), .A2(\DataP/alu_a_in[1] ), .B1(n1605), .B2(n2711), .ZN(n2848) );
  AOI221_X1 U3385 ( .B1(n2933), .B2(n2839), .C1(n2848), .C2(n2988), .A(n2842), 
        .ZN(n2849) );
  AOI21_X1 U3386 ( .B1(n2842), .B2(n2950), .A(n2849), .ZN(n2850) );
  AOI22_X1 U3387 ( .A1(n2846), .A2(n2975), .B1(n2850), .B2(n2064), .ZN(n2851)
         );
  MUX2_X1 U3388 ( .A(n2893), .B(n2851), .S(n2847), .Z(
        \DataP/ALU_C/shifter/N82 ) );
  AOI22_X1 U3389 ( .A1(\sra_131/SH[1] ), .A2(n1923), .B1(n2852), .B2(n2988), 
        .ZN(n2882) );
  AOI22_X1 U3390 ( .A1(\sra_131/SH[1] ), .A2(n2854), .B1(n2853), .B2(n2988), 
        .ZN(n2884) );
  AOI22_X1 U3391 ( .A1(n2841), .A2(n2882), .B1(n2884), .B2(n2989), .ZN(n2900)
         );
  NAND2_X1 U3392 ( .A1(n2846), .A2(\DataP/alu_a_in[31] ), .ZN(n2920) );
  OAI21_X1 U3393 ( .B1(n1915), .B2(n2900), .A(n2920), .ZN(n2924) );
  AOI22_X1 U3394 ( .A1(\sra_131/SH[1] ), .A2(n2856), .B1(n2855), .B2(n2988), 
        .ZN(n2883) );
  AOI22_X1 U3395 ( .A1(\sra_131/SH[1] ), .A2(n2858), .B1(n2857), .B2(n2988), 
        .ZN(n2886) );
  AOI22_X1 U3396 ( .A1(n2841), .A2(n2883), .B1(n2886), .B2(n2989), .ZN(n2899)
         );
  AOI22_X1 U3397 ( .A1(\sra_131/SH[1] ), .A2(n2860), .B1(n2859), .B2(n2988), 
        .ZN(n2885) );
  AOI22_X1 U3398 ( .A1(n2839), .A2(n2862), .B1(n2861), .B2(n2988), .ZN(n2965)
         );
  AOI22_X1 U3399 ( .A1(n2841), .A2(n2885), .B1(n2965), .B2(n2989), .ZN(n2936)
         );
  AOI22_X1 U3400 ( .A1(n2846), .A2(n2899), .B1(n2936), .B2(n2127), .ZN(n2863)
         );
  MUX2_X1 U3401 ( .A(n2924), .B(n2863), .S(n2847), .Z(
        \DataP/ALU_C/shifter/N92 ) );
  AOI22_X1 U3402 ( .A1(n2987), .A2(\DataP/alu_a_in[30] ), .B1(
        \DataP/alu_a_in[29] ), .B2(n2985), .ZN(n2871) );
  AOI22_X1 U3403 ( .A1(n2987), .A2(\DataP/alu_a_in[28] ), .B1(
        \DataP/alu_a_in[27] ), .B2(n2985), .ZN(n2873) );
  AOI22_X1 U3404 ( .A1(n2839), .A2(n2871), .B1(n2873), .B2(n2988), .ZN(n2889)
         );
  NOR2_X1 U3405 ( .A1(n1913), .A2(n1923), .ZN(n2881) );
  AOI21_X1 U3406 ( .B1(n1913), .B2(n2889), .A(n2881), .ZN(n2902) );
  OAI21_X1 U3407 ( .B1(n2846), .B2(n2902), .A(n2920), .ZN(n2925) );
  AOI22_X1 U3408 ( .A1(n2709), .A2(\DataP/alu_a_in[26] ), .B1(
        \DataP/alu_a_in[25] ), .B2(n2711), .ZN(n2872) );
  AOI22_X1 U3409 ( .A1(n2987), .A2(\DataP/alu_a_in[24] ), .B1(
        \DataP/alu_a_in[23] ), .B2(n2710), .ZN(n2875) );
  AOI22_X1 U3410 ( .A1(n2839), .A2(n2872), .B1(n2875), .B2(n2988), .ZN(n2888)
         );
  AOI22_X1 U3411 ( .A1(n2987), .A2(\DataP/alu_a_in[22] ), .B1(
        \DataP/alu_a_in[21] ), .B2(n2985), .ZN(n2874) );
  AOI22_X1 U3412 ( .A1(n2987), .A2(\DataP/alu_a_in[20] ), .B1(n1553), .B2(
        n2985), .ZN(n2877) );
  AOI22_X1 U3413 ( .A1(\sra_131/SH[1] ), .A2(n2874), .B1(n2877), .B2(n2988), 
        .ZN(n2891) );
  AOI22_X1 U3414 ( .A1(n2841), .A2(n2888), .B1(n2891), .B2(n2989), .ZN(n2901)
         );
  AOI22_X1 U3415 ( .A1(n2987), .A2(\DataP/alu_a_in[18] ), .B1(
        \DataP/alu_a_in[17] ), .B2(n2985), .ZN(n2876) );
  AOI22_X1 U3416 ( .A1(n2987), .A2(\DataP/alu_a_in[16] ), .B1(n1841), .B2(
        n2985), .ZN(n2879) );
  AOI22_X1 U3417 ( .A1(\sra_131/SH[1] ), .A2(n2876), .B1(n2879), .B2(n2988), 
        .ZN(n2890) );
  AOI22_X1 U3418 ( .A1(n2987), .A2(\DataP/alu_a_in[14] ), .B1(
        \DataP/alu_a_in[13] ), .B2(n2985), .ZN(n2878) );
  AOI22_X1 U3419 ( .A1(n2987), .A2(\DataP/alu_a_in[12] ), .B1(
        \DataP/alu_a_in[11] ), .B2(n2711), .ZN(n2903) );
  AOI22_X1 U3420 ( .A1(\sra_131/SH[1] ), .A2(n2878), .B1(n2903), .B2(n2988), 
        .ZN(n2970) );
  AOI22_X1 U3421 ( .A1(n2841), .A2(n2890), .B1(n2970), .B2(n1913), .ZN(n2946)
         );
  AOI22_X1 U3422 ( .A1(n1915), .A2(n2901), .B1(n2946), .B2(n2127), .ZN(n2864)
         );
  MUX2_X1 U3423 ( .A(n2925), .B(n2864), .S(n2065), .Z(
        \DataP/ALU_C/shifter/N93 ) );
  AOI21_X1 U3424 ( .B1(n2989), .B2(n2865), .A(n2881), .ZN(n2911) );
  OAI21_X1 U3425 ( .B1(n1915), .B2(n2911), .A(n2920), .ZN(n2927) );
  AOI22_X1 U3426 ( .A1(n2841), .A2(n2867), .B1(n2866), .B2(n1913), .ZN(n2910)
         );
  AOI22_X1 U3427 ( .A1(n2841), .A2(n2869), .B1(n2868), .B2(n1913), .ZN(n2953)
         );
  AOI22_X1 U3428 ( .A1(n1915), .A2(n2910), .B1(n2953), .B2(n2064), .ZN(n2870)
         );
  MUX2_X1 U3429 ( .A(n2927), .B(n2870), .S(n2847), .Z(
        \DataP/ALU_C/shifter/N94 ) );
  AOI22_X1 U3430 ( .A1(\sra_131/SH[1] ), .A2(n1923), .B1(n2871), .B2(n2988), 
        .ZN(n2896) );
  AOI21_X1 U3431 ( .B1(n1913), .B2(n2896), .A(n2881), .ZN(n2913) );
  OAI21_X1 U3432 ( .B1(n2846), .B2(n2913), .A(n2920), .ZN(n2929) );
  AOI22_X1 U3433 ( .A1(n2840), .A2(n2873), .B1(n2872), .B2(n2988), .ZN(n2895)
         );
  AOI22_X1 U3434 ( .A1(n2839), .A2(n2875), .B1(n2874), .B2(n2988), .ZN(n2898)
         );
  AOI22_X1 U3435 ( .A1(n2841), .A2(n2895), .B1(n2898), .B2(n1913), .ZN(n2912)
         );
  AOI22_X1 U3436 ( .A1(n2839), .A2(n2877), .B1(n2876), .B2(n2988), .ZN(n2897)
         );
  AOI22_X1 U3437 ( .A1(\sra_131/SH[1] ), .A2(n2879), .B1(n2878), .B2(n2988), 
        .ZN(n2904) );
  AOI22_X1 U3438 ( .A1(n2841), .A2(n2897), .B1(n2904), .B2(n1913), .ZN(n2960)
         );
  AOI22_X1 U3439 ( .A1(n1915), .A2(n2912), .B1(n2960), .B2(n2064), .ZN(n2880)
         );
  MUX2_X1 U3440 ( .A(n2929), .B(n2880), .S(n2065), .Z(
        \DataP/ALU_C/shifter/N95 ) );
  AOI21_X1 U3441 ( .B1(n1913), .B2(n2882), .A(n2881), .ZN(n2915) );
  OAI21_X1 U3442 ( .B1(n1915), .B2(n2915), .A(n2920), .ZN(n2938) );
  AOI22_X1 U3443 ( .A1(n2841), .A2(n2884), .B1(n2883), .B2(n1913), .ZN(n2914)
         );
  AOI22_X1 U3444 ( .A1(n2841), .A2(n2886), .B1(n2885), .B2(n1913), .ZN(n2966)
         );
  AOI22_X1 U3445 ( .A1(n2846), .A2(n2914), .B1(n2966), .B2(n2127), .ZN(n2887)
         );
  MUX2_X1 U3446 ( .A(n2938), .B(n2887), .S(n2847), .Z(
        \DataP/ALU_C/shifter/N96 ) );
  NAND2_X1 U3447 ( .A1(\lt_x_134/B[4] ), .A2(\DataP/alu_a_in[31] ), .ZN(n2923)
         );
  AOI22_X1 U3448 ( .A1(n2841), .A2(n2889), .B1(n2888), .B2(n1913), .ZN(n2916)
         );
  AOI22_X1 U3449 ( .A1(n2841), .A2(n2891), .B1(n2890), .B2(n1913), .ZN(n2972)
         );
  AOI221_X1 U3450 ( .B1(n2916), .B2(n2846), .C1(n2972), .C2(n2064), .A(
        \lt_x_134/B[4] ), .ZN(n2892) );
  OR2_X1 U3451 ( .A1(n2981), .A2(n2892), .ZN(\DataP/ALU_C/shifter/N97 ) );
  AOI21_X1 U3452 ( .B1(n2847), .B2(n2893), .A(n2981), .ZN(n2894) );
  AOI22_X1 U3453 ( .A1(n2841), .A2(n2896), .B1(n2895), .B2(n1913), .ZN(n2921)
         );
  AOI22_X1 U3454 ( .A1(n2841), .A2(n2898), .B1(n2897), .B2(n1913), .ZN(n2979)
         );
  MUX2_X1 U3455 ( .A(n2921), .B(n2979), .S(n2064), .Z(n2909) );
  OAI21_X1 U3456 ( .B1(\lt_x_134/B[4] ), .B2(n2909), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N99 ) );
  MUX2_X1 U3457 ( .A(n2900), .B(n2899), .S(n2127), .Z(n2937) );
  OAI21_X1 U3458 ( .B1(\lt_x_134/B[4] ), .B2(n2937), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N100 ) );
  MUX2_X1 U3459 ( .A(n2902), .B(n2901), .S(n2064), .Z(n2949) );
  OAI21_X1 U3460 ( .B1(\lt_x_135/B[4] ), .B2(n2949), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N101 ) );
  AOI22_X1 U3461 ( .A1(n2987), .A2(\DataP/alu_a_in[10] ), .B1(
        \DataP/alu_a_in[9] ), .B2(n2710), .ZN(n2941) );
  AOI22_X1 U3462 ( .A1(n1612), .A2(n2903), .B1(n2941), .B2(n2988), .ZN(n2958)
         );
  AOI22_X1 U3463 ( .A1(n2841), .A2(n2904), .B1(n2958), .B2(n2989), .ZN(n2978)
         );
  AOI22_X1 U3464 ( .A1(n2987), .A2(\DataP/alu_a_in[8] ), .B1(
        \DataP/alu_a_in[7] ), .B2(n2710), .ZN(n2940) );
  AOI22_X1 U3465 ( .A1(n2987), .A2(\DataP/alu_a_in[6] ), .B1(
        \DataP/alu_a_in[5] ), .B2(n2985), .ZN(n2943) );
  AOI22_X1 U3466 ( .A1(n2839), .A2(n2940), .B1(n2943), .B2(n2988), .ZN(n2957)
         );
  AOI22_X1 U3467 ( .A1(n2987), .A2(\DataP/alu_a_in[4] ), .B1(
        \DataP/alu_a_in[3] ), .B2(n2711), .ZN(n2942) );
  AOI22_X1 U3468 ( .A1(n2841), .A2(n2957), .B1(n2905), .B2(n2989), .ZN(n2906)
         );
  AOI22_X1 U3469 ( .A1(n1915), .A2(n2978), .B1(n2906), .B2(n2845), .ZN(n2907)
         );
  NAND2_X1 U3470 ( .A1(n2847), .A2(n2907), .ZN(n2908) );
  OAI21_X1 U3471 ( .B1(n2847), .B2(n2909), .A(n2908), .ZN(
        \DataP/ALU_C/shifter/N83 ) );
  MUX2_X1 U3472 ( .A(n2911), .B(n2910), .S(n2127), .Z(n2956) );
  OAI21_X1 U3473 ( .B1(\lt_x_135/B[4] ), .B2(n2956), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N102 ) );
  MUX2_X1 U3474 ( .A(n2913), .B(n2912), .S(n2064), .Z(n2963) );
  OAI21_X1 U3475 ( .B1(\lt_x_134/B[4] ), .B2(n2963), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N103 ) );
  MUX2_X1 U3476 ( .A(n2915), .B(n2914), .S(n2127), .Z(n2968) );
  OAI21_X1 U3477 ( .B1(\lt_x_134/B[4] ), .B2(n2968), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N104 ) );
  OAI21_X1 U3478 ( .B1(n1915), .B2(n2916), .A(n2920), .ZN(n2917) );
  OAI21_X1 U3479 ( .B1(\lt_x_135/B[4] ), .B2(n2982), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N105 ) );
  OAI21_X1 U3480 ( .B1(n1915), .B2(n2918), .A(n2920), .ZN(n2919) );
  OAI21_X1 U3481 ( .B1(\lt_x_134/B[4] ), .B2(n2983), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N106 ) );
  OAI21_X1 U3482 ( .B1(n2846), .B2(n2921), .A(n2920), .ZN(n2922) );
  OAI21_X1 U3483 ( .B1(\lt_x_134/B[4] ), .B2(n2984), .A(n2923), .ZN(
        \DataP/ALU_C/shifter/N107 ) );
  AOI21_X1 U3484 ( .B1(n2065), .B2(n2927), .A(n2981), .ZN(n2928) );
  AOI22_X1 U3485 ( .A1(\sra_131/SH[1] ), .A2(n2932), .B1(n2931), .B2(n2988), 
        .ZN(n2964) );
  AOI22_X1 U3486 ( .A1(n1612), .A2(n2934), .B1(n2933), .B2(n2988), .ZN(n2935)
         );
  AOI21_X1 U3487 ( .B1(n2847), .B2(n2938), .A(n2981), .ZN(n2939) );
  AOI22_X1 U3488 ( .A1(n2840), .A2(n2941), .B1(n2940), .B2(n2988), .ZN(n2969)
         );
  AOI22_X1 U3489 ( .A1(n2839), .A2(n2943), .B1(n2942), .B2(n2988), .ZN(n2944)
         );
  AOI22_X1 U3490 ( .A1(n2841), .A2(n2969), .B1(n2944), .B2(n2989), .ZN(n2945)
         );
  AOI22_X1 U3491 ( .A1(n2846), .A2(n2946), .B1(n2945), .B2(n2064), .ZN(n2947)
         );
  NAND2_X1 U3492 ( .A1(n2065), .A2(n2947), .ZN(n2948) );
  AOI22_X1 U3493 ( .A1(n2841), .A2(n2951), .B1(n2950), .B2(n2989), .ZN(n2952)
         );
  AOI22_X1 U3494 ( .A1(n2846), .A2(n2953), .B1(n2952), .B2(n2845), .ZN(n2954)
         );
  NAND2_X1 U3495 ( .A1(n2847), .A2(n2954), .ZN(n2955) );
  AOI22_X1 U3496 ( .A1(n2842), .A2(n2958), .B1(n2957), .B2(n2989), .ZN(n2959)
         );
  AOI22_X1 U3497 ( .A1(n1915), .A2(n2960), .B1(n2959), .B2(n2845), .ZN(n2961)
         );
  NAND2_X1 U3498 ( .A1(n2065), .A2(n2961), .ZN(n2962) );
  AOI22_X1 U3499 ( .A1(n2841), .A2(n2970), .B1(n2969), .B2(n2989), .ZN(n2971)
         );
  AOI22_X1 U3500 ( .A1(n1915), .A2(n2972), .B1(n2971), .B2(n2845), .ZN(n2973)
         );
  NAND2_X1 U3501 ( .A1(n2847), .A2(n2973), .ZN(n2974) );
  OAI21_X1 U3502 ( .B1(n2065), .B2(n2982), .A(n2974), .ZN(
        \DataP/ALU_C/shifter/N89 ) );
  INV_X1 U3503 ( .A(n2985), .ZN(n2986) );
  INV_X1 U3504 ( .A(n2841), .ZN(n2989) );
  INV_X1 U3505 ( .A(n2994), .ZN(n2993) );
  INV_X1 U3506 ( .A(n1845), .ZN(n2997) );
  XOR2_X1 U3507 ( .A(\DataP/dest_M[4] ), .B(n524), .Z(n3052) );
  XOR2_X1 U3508 ( .A(\DataP/dest_M[3] ), .B(n523), .Z(n3051) );
  NAND3_X1 U3509 ( .A1(n3053), .A2(n3052), .A3(n3051), .ZN(n3056) );
  NAND3_X1 U3510 ( .A1(n2994), .A2(n432), .A3(n1844), .ZN(n3194) );
  NAND3_X1 U3511 ( .A1(n3199), .A2(n443), .A3(ALU_OPCODE_i[3]), .ZN(n3200) );
  NAND3_X1 U3512 ( .A1(ALU_OPCODE_i[0]), .A2(ALU_OPCODE_i[3]), .A3(n3222), 
        .ZN(n3695) );
  NAND3_X1 U3513 ( .A1(\DataP/alu_a_in[11] ), .A2(n3689), .A3(n1572), .ZN(
        n3271) );
  XOR2_X1 U3514 ( .A(n3273), .B(n1601), .Z(n3279) );
  NAND3_X1 U3515 ( .A1(\DataP/alu_a_in[12] ), .A2(n3693), .A3(n1880), .ZN(
        n3274) );
  MUX2_X1 U3516 ( .A(n3341), .B(n3343), .S(ALU_OPCODE_i[1]), .Z(n3342) );
  NAND3_X1 U3517 ( .A1(n1602), .A2(n3343), .A3(n2144), .ZN(n3344) );
  NAND3_X1 U3518 ( .A1(n3348), .A2(ALU_OPCODE_i[3]), .A3(n2150), .ZN(n3355) );
  XOR2_X1 U3519 ( .A(n3361), .B(n3360), .Z(n3367) );
  MUX2_X1 U3520 ( .A(n3391), .B(n3402), .S(n3689), .Z(n3393) );
  NAND3_X1 U3521 ( .A1(n1841), .A2(n3689), .A3(\DataP/alu_b_in[15] ), .ZN(
        n3415) );
  NAND3_X1 U3522 ( .A1(n3434), .A2(n3433), .A3(n3432), .ZN(n3435) );
  NAND3_X1 U3523 ( .A1(n3438), .A2(n3468), .A3(n1933), .ZN(n3439) );
  MUX2_X1 U3524 ( .A(\DataP/alu_b_in[23] ), .B(n3440), .S(n3510), .Z(n3464) );
  MUX2_X1 U3525 ( .A(n3446), .B(n1933), .S(n3689), .Z(n3447) );
  MUX2_X1 U3526 ( .A(n3469), .B(\DataP/alu_b_in[24] ), .S(n3689), .Z(n3471) );
  MUX2_X1 U3527 ( .A(n3492), .B(n3491), .S(n3510), .Z(n3493) );
  NAND3_X1 U3528 ( .A1(n1849), .A2(n3499), .A3(n3500), .ZN(n3503) );
  NAND3_X1 U3529 ( .A1(n3540), .A2(n3539), .A3(n3538), .ZN(n3541) );
  XOR2_X1 U3530 ( .A(n3545), .B(n3546), .Z(n3553) );
  NAND3_X1 U3531 ( .A1(n3551), .A2(n3550), .A3(n3549), .ZN(n3552) );
  NAND3_X1 U3532 ( .A1(n3561), .A2(n3560), .A3(n3559), .ZN(n3562) );
  XOR2_X1 U3533 ( .A(n3582), .B(n3581), .Z(n3591) );
  XOR2_X1 U3534 ( .A(n1533), .B(n1989), .Z(n3601) );
  NAND3_X1 U3535 ( .A1(n3599), .A2(n3598), .A3(n3597), .ZN(n3600) );
  NAND3_X1 U3536 ( .A1(n3619), .A2(n3618), .A3(n3617), .ZN(n3620) );
  XOR2_X1 U3537 ( .A(n2239), .B(n1986), .Z(n3630) );
  NAND3_X1 U3538 ( .A1(\DataP/alu_a_in[16] ), .A2(n3693), .A3(
        \DataP/alu_b_in[16] ), .ZN(n3623) );
  NAND3_X1 U3539 ( .A1(n3628), .A2(n3627), .A3(n3626), .ZN(n3629) );
  NAND3_X1 U3540 ( .A1(\DataP/alu_a_in[13] ), .A2(n3693), .A3(n1860), .ZN(
        n3649) );
  MUX2_X1 U3541 ( .A(n3661), .B(n3679), .S(\DataP/alu_a_in[8] ), .Z(n3664) );
  NAND3_X1 U3542 ( .A1(n3696), .A2(n3695), .A3(n3694), .ZN(n3698) );
  AOI22_X1 U3543 ( .A1(n1940), .A2(\DataP/npc_pre[30] ), .B1(
        \DataP/pc_out[30] ), .B2(n3010), .ZN(n3769) );
  AOI22_X1 U3544 ( .A1(n1940), .A2(\DataP/npc_pre[28] ), .B1(
        \DataP/pc_out[28] ), .B2(n3010), .ZN(n3753) );
  AOI22_X1 U3545 ( .A1(n1940), .A2(\DataP/npc_pre[26] ), .B1(
        \DataP/pc_out[26] ), .B2(n3010), .ZN(n3754) );
  AOI22_X1 U3546 ( .A1(n1940), .A2(\DataP/npc_pre[24] ), .B1(
        \DataP/pc_out[24] ), .B2(n3010), .ZN(n3764) );
  AOI22_X1 U3547 ( .A1(n1940), .A2(\DataP/npc_pre[22] ), .B1(
        \DataP/pc_out[22] ), .B2(n3010), .ZN(n3763) );
  AOI22_X1 U3548 ( .A1(n1940), .A2(\DataP/npc_pre[20] ), .B1(
        \DataP/pc_out[20] ), .B2(n3010), .ZN(n3760) );
  AOI22_X1 U3549 ( .A1(n1940), .A2(\DataP/npc_pre[18] ), .B1(
        \DataP/pc_out[18] ), .B2(n3010), .ZN(n3765) );
  AOI22_X1 U3550 ( .A1(n1940), .A2(\DataP/npc_pre[16] ), .B1(
        \DataP/pc_out[16] ), .B2(n3010), .ZN(n3759) );
  AOI22_X1 U3551 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[14] ), .B1(
        \DataP/pc_out[14] ), .B2(n3010), .ZN(n3758) );
  AOI22_X1 U3552 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[12] ), .B1(
        \DataP/pc_out[12] ), .B2(n3010), .ZN(n3766) );
  AOI22_X1 U3553 ( .A1(n1940), .A2(\DataP/npc_pre[10] ), .B1(
        \DataP/pc_out[10] ), .B2(n3010), .ZN(n3774) );
  AOI22_X1 U3554 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[8] ), .B1(
        IRAM_ADDRESS[6]), .B2(n3010), .ZN(n3736) );
  AOI22_X1 U3555 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[6] ), .B1(
        IRAM_ADDRESS[4]), .B2(n3010), .ZN(n3742) );
  AOI22_X1 U3556 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[4] ), .B1(
        IRAM_ADDRESS[2]), .B2(n3010), .ZN(n3749) );
  AOI22_X1 U3557 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[2] ), .B1(
        IRAM_ADDRESS[0]), .B2(n3010), .ZN(\DataP/NPC_add/N3 ) );
  AOI22_X1 U3558 ( .A1(\DataP/npc_mux_sel ), .A2(\DataP/npc_pre[3] ), .B1(
        IRAM_ADDRESS[1]), .B2(n3010), .ZN(n3751) );
  NOR2_X1 U3559 ( .A1(\DataP/NPC_add/N3 ), .A2(n3751), .ZN(n3750) );
  INV_X1 U3560 ( .A(n3750), .ZN(n3748) );
  NOR2_X1 U3561 ( .A1(n3749), .A2(n3748), .ZN(n3747) );
  OAI221_X1 U3562 ( .B1(n1940), .B2(IRAM_ADDRESS[3]), .C1(n3010), .C2(
        \DataP/npc_pre[5] ), .A(n3747), .ZN(n3743) );
  NOR2_X1 U3563 ( .A1(n3742), .A2(n3743), .ZN(n3741) );
  OAI221_X1 U3564 ( .B1(n1940), .B2(IRAM_ADDRESS[5]), .C1(n3010), .C2(
        \DataP/npc_pre[7] ), .A(n3741), .ZN(n3737) );
  NOR2_X1 U3565 ( .A1(n3736), .A2(n3737), .ZN(n3735) );
  OAI221_X1 U3566 ( .B1(n1940), .B2(IRAM_ADDRESS[7]), .C1(n3010), .C2(
        \DataP/npc_pre[9] ), .A(n3735), .ZN(n3773) );
  NOR2_X1 U3567 ( .A1(n3774), .A2(n3773), .ZN(n3731) );
  MUX2_X1 U3568 ( .A(\DataP/pc_out[11] ), .B(\DataP/npc_pre[11] ), .S(n1940), 
        .Z(n3770) );
  NAND2_X1 U3569 ( .A1(n3731), .A2(n3770), .ZN(n3730) );
  NOR2_X1 U3570 ( .A1(n3766), .A2(n3730), .ZN(n3729) );
  MUX2_X1 U3571 ( .A(\DataP/pc_out[13] ), .B(\DataP/npc_pre[13] ), .S(n1940), 
        .Z(n3761) );
  NAND2_X1 U3572 ( .A1(n3729), .A2(n3761), .ZN(n3728) );
  NOR2_X1 U3573 ( .A1(n3758), .A2(n3728), .ZN(n3727) );
  MUX2_X1 U3574 ( .A(\DataP/pc_out[15] ), .B(\DataP/npc_pre[15] ), .S(n1940), 
        .Z(n3757) );
  NAND2_X1 U3575 ( .A1(n3727), .A2(n3757), .ZN(n3726) );
  NOR2_X1 U3576 ( .A1(n3759), .A2(n3726), .ZN(n3725) );
  MUX2_X1 U3577 ( .A(\DataP/pc_out[17] ), .B(\DataP/npc_pre[17] ), .S(n1940), 
        .Z(n3767) );
  NAND2_X1 U3578 ( .A1(n3725), .A2(n3767), .ZN(n3724) );
  NOR2_X1 U3579 ( .A1(n3765), .A2(n3724), .ZN(n3723) );
  MUX2_X1 U3580 ( .A(\DataP/pc_out[19] ), .B(\DataP/npc_pre[19] ), .S(n1940), 
        .Z(n3762) );
  NAND2_X1 U3581 ( .A1(n3723), .A2(n3762), .ZN(n3722) );
  NOR2_X1 U3582 ( .A1(n3760), .A2(n3722), .ZN(n3721) );
  MUX2_X1 U3583 ( .A(\DataP/pc_out[21] ), .B(\DataP/npc_pre[21] ), .S(n1940), 
        .Z(n3771) );
  NAND2_X1 U3584 ( .A1(n3721), .A2(n3771), .ZN(n3720) );
  NOR2_X1 U3585 ( .A1(n3763), .A2(n3720), .ZN(n3719) );
  MUX2_X1 U3586 ( .A(\DataP/pc_out[23] ), .B(\DataP/npc_pre[23] ), .S(n1940), 
        .Z(n3772) );
  NAND2_X1 U3587 ( .A1(n3719), .A2(n3772), .ZN(n3718) );
  NOR2_X1 U3588 ( .A1(n3764), .A2(n3718), .ZN(n3717) );
  MUX2_X1 U3589 ( .A(\DataP/pc_out[25] ), .B(\DataP/npc_pre[25] ), .S(n1940), 
        .Z(n3755) );
  NAND2_X1 U3590 ( .A1(n3717), .A2(n3755), .ZN(n3716) );
  NOR2_X1 U3591 ( .A1(n3754), .A2(n3716), .ZN(n3715) );
  MUX2_X1 U3592 ( .A(\DataP/pc_out[27] ), .B(\DataP/npc_pre[27] ), .S(n1940), 
        .Z(n3756) );
  NAND2_X1 U3593 ( .A1(n3715), .A2(n3756), .ZN(n3714) );
  NOR2_X1 U3594 ( .A1(n3753), .A2(n3714), .ZN(n3713) );
  MUX2_X1 U3595 ( .A(\DataP/pc_out[29] ), .B(\DataP/npc_pre[29] ), .S(n1940), 
        .Z(n3768) );
  NAND2_X1 U3596 ( .A1(n3713), .A2(n3768), .ZN(n3712) );
  NOR2_X1 U3597 ( .A1(n3769), .A2(n3712), .ZN(n3752) );
  AOI21_X1 U3598 ( .B1(n3769), .B2(n3712), .A(n3752), .ZN(\DataP/NPC_add/N31 )
         );
  XOR2_X1 U3599 ( .A(n3713), .B(n3768), .Z(\DataP/NPC_add/N30 ) );
  AOI21_X1 U3600 ( .B1(n3753), .B2(n3714), .A(n3713), .ZN(\DataP/NPC_add/N29 )
         );
  XOR2_X1 U3601 ( .A(n3715), .B(n3756), .Z(\DataP/NPC_add/N28 ) );
  AOI21_X1 U3602 ( .B1(n3754), .B2(n3716), .A(n3715), .ZN(\DataP/NPC_add/N27 )
         );
  XOR2_X1 U3603 ( .A(n3717), .B(n3755), .Z(\DataP/NPC_add/N26 ) );
  AOI21_X1 U3604 ( .B1(n3764), .B2(n3718), .A(n3717), .ZN(\DataP/NPC_add/N25 )
         );
  XOR2_X1 U3605 ( .A(n3719), .B(n3772), .Z(\DataP/NPC_add/N24 ) );
  AOI21_X1 U3606 ( .B1(n3763), .B2(n3720), .A(n3719), .ZN(\DataP/NPC_add/N23 )
         );
  XOR2_X1 U3607 ( .A(n3721), .B(n3771), .Z(\DataP/NPC_add/N22 ) );
  AOI21_X1 U3608 ( .B1(n3760), .B2(n3722), .A(n3721), .ZN(\DataP/NPC_add/N21 )
         );
  XOR2_X1 U3609 ( .A(n3723), .B(n3762), .Z(\DataP/NPC_add/N20 ) );
  AOI21_X1 U3610 ( .B1(n3765), .B2(n3724), .A(n3723), .ZN(\DataP/NPC_add/N19 )
         );
  XOR2_X1 U3611 ( .A(n3725), .B(n3767), .Z(\DataP/NPC_add/N18 ) );
  AOI21_X1 U3612 ( .B1(n3759), .B2(n3726), .A(n3725), .ZN(\DataP/NPC_add/N17 )
         );
  XOR2_X1 U3613 ( .A(n3727), .B(n3757), .Z(\DataP/NPC_add/N16 ) );
  AOI21_X1 U3614 ( .B1(n3758), .B2(n3728), .A(n3727), .ZN(\DataP/NPC_add/N15 )
         );
  XOR2_X1 U3615 ( .A(n3729), .B(n3761), .Z(\DataP/NPC_add/N14 ) );
  AOI21_X1 U3616 ( .B1(n3766), .B2(n3730), .A(n3729), .ZN(\DataP/NPC_add/N13 )
         );
  XOR2_X1 U3617 ( .A(n3731), .B(n3770), .Z(\DataP/NPC_add/N12 ) );
  AOI21_X1 U3618 ( .B1(n3774), .B2(n3773), .A(n3731), .ZN(\DataP/NPC_add/N11 )
         );
  AOI22_X1 U3619 ( .A1(n1940), .A2(\DataP/npc_pre[9] ), .B1(IRAM_ADDRESS[7]), 
        .B2(n3010), .ZN(n3734) );
  INV_X1 U3620 ( .A(n3735), .ZN(n3733) );
  INV_X1 U3621 ( .A(n3773), .ZN(n3732) );
  AOI21_X1 U3622 ( .B1(n3734), .B2(n3733), .A(n3732), .ZN(\DataP/NPC_add/N10 )
         );
  AOI21_X1 U3623 ( .B1(n3736), .B2(n3737), .A(n3735), .ZN(\DataP/NPC_add/N9 )
         );
  AOI22_X1 U3624 ( .A1(n1940), .A2(\DataP/npc_pre[7] ), .B1(IRAM_ADDRESS[5]), 
        .B2(n3010), .ZN(n3740) );
  INV_X1 U3625 ( .A(n3741), .ZN(n3739) );
  INV_X1 U3626 ( .A(n3737), .ZN(n3738) );
  AOI21_X1 U3627 ( .B1(n3740), .B2(n3739), .A(n3738), .ZN(\DataP/NPC_add/N8 )
         );
  AOI21_X1 U3628 ( .B1(n3742), .B2(n3743), .A(n3741), .ZN(\DataP/NPC_add/N7 )
         );
  AOI22_X1 U3629 ( .A1(n1940), .A2(\DataP/npc_pre[5] ), .B1(IRAM_ADDRESS[3]), 
        .B2(n3010), .ZN(n3746) );
  INV_X1 U3630 ( .A(n3747), .ZN(n3745) );
  INV_X1 U3631 ( .A(n3743), .ZN(n3744) );
  AOI21_X1 U3632 ( .B1(n3746), .B2(n3745), .A(n3744), .ZN(\DataP/NPC_add/N6 )
         );
  AOI21_X1 U3633 ( .B1(n3749), .B2(n3748), .A(n3747), .ZN(\DataP/NPC_add/N5 )
         );
  AOI21_X1 U3634 ( .B1(n3751), .B2(\DataP/NPC_add/N3 ), .A(n3750), .ZN(
        \DataP/NPC_add/N4 ) );
  AOI22_X1 U3635 ( .A1(n1940), .A2(\DataP/npc_pre[31] ), .B1(
        \DataP/pc_out[31] ), .B2(n3010), .ZN(n3775) );
  XNOR2_X1 U3636 ( .A(n3775), .B(n3752), .ZN(\DataP/NPC_add/N32 ) );
  NAND2_X1 U3639 ( .A1(IR_CU_28), .A2(n516), .ZN(n3781) );
  NOR2_X1 U3640 ( .A1(n3955), .A2(n3781), .ZN(n606) );
  NAND2_X1 U3641 ( .A1(IR_CU_27), .A2(n497), .ZN(n3951) );
  NOR2_X1 U3642 ( .A1(n514), .A2(n515), .ZN(n3976) );
  NAND3_X1 U3643 ( .A1(IR_CU_31), .A2(n3976), .A3(n510), .ZN(n3813) );
  NOR2_X1 U3644 ( .A1(IR_CU_27), .A2(n497), .ZN(n3797) );
  INV_X1 U3645 ( .A(n3976), .ZN(n3977) );
  NOR2_X1 U3646 ( .A1(n3781), .A2(n3977), .ZN(n3814) );
  NOR3_X1 U3647 ( .A1(IR_CU_27), .A2(n3955), .A3(n516), .ZN(n3847) );
  AOI22_X1 U3648 ( .A1(IR_CU_31), .A2(n3966), .B1(n2141), .B2(n504), .ZN(n3776) );
  NAND2_X1 U3649 ( .A1(n515), .A2(n510), .ZN(n3845) );
  NOR3_X1 U3650 ( .A1(n514), .A2(n2129), .A3(n3781), .ZN(n3796) );
  AOI22_X1 U3651 ( .A1(n3856), .A2(n606), .B1(n3853), .B2(n3796), .ZN(n3798)
         );
  OAI211_X1 U3652 ( .C1(n3776), .C2(n3845), .A(n3798), .B(n3956), .ZN(n3777)
         );
  AOI211_X1 U3653 ( .C1(n3797), .C2(n3814), .A(n3847), .B(n3777), .ZN(n3788)
         );
  NOR4_X1 U3654 ( .A1(IR_CU[8]), .A2(IR_CU[6]), .A3(IR_CU[7]), .A4(IR_CU[9]), 
        .ZN(n3778) );
  NAND3_X1 U3655 ( .A1(n3953), .A2(n484), .A3(n3778), .ZN(n3790) );
  NOR2_X1 U3656 ( .A1(n479), .A2(n3790), .ZN(n3824) );
  NAND2_X1 U3657 ( .A1(IR_CU[5]), .A2(n3824), .ZN(n3802) );
  NOR3_X1 U3658 ( .A1(n477), .A2(n2128), .A3(n3802), .ZN(n3786) );
  NOR3_X1 U3659 ( .A1(n478), .A2(n3790), .A3(n2135), .ZN(n3804) );
  NAND2_X1 U3660 ( .A1(n3804), .A2(n476), .ZN(n3806) );
  OAI21_X1 U3661 ( .B1(n476), .B2(n479), .A(n2128), .ZN(n3779) );
  OAI211_X1 U3662 ( .C1(n479), .C2(n2128), .A(n3779), .B(n477), .ZN(n3780) );
  NAND2_X1 U3663 ( .A1(IR_CU[5]), .A2(n480), .ZN(n3836) );
  AOI221_X1 U3664 ( .B1(n3790), .B2(n3806), .C1(n3780), .C2(n3806), .A(n3836), 
        .ZN(n3785) );
  INV_X1 U3665 ( .A(n3786), .ZN(n3833) );
  NOR3_X1 U3666 ( .A1(n3795), .A2(n3955), .A3(n3951), .ZN(n3821) );
  INV_X1 U3667 ( .A(n3781), .ZN(n3782) );
  NAND3_X1 U3668 ( .A1(n514), .A2(n3782), .A3(n2129), .ZN(n3817) );
  NAND4_X1 U3669 ( .A1(n3804), .A2(IR_CU[1]), .A3(n480), .A4(n482), .ZN(n3827)
         );
  OAI21_X1 U3670 ( .B1(n504), .B2(n3817), .A(n3827), .ZN(n3801) );
  AOI211_X1 U3671 ( .C1(n3856), .C2(n3796), .A(n3821), .B(n3801), .ZN(n3784)
         );
  NAND3_X1 U3672 ( .A1(n3966), .A2(n3976), .A3(n510), .ZN(n3783) );
  OAI211_X1 U3673 ( .C1(n3833), .C2(n476), .A(n3784), .B(n3783), .ZN(n3792) );
  AOI211_X1 U3674 ( .C1(n3786), .C2(IR_CU[4]), .A(n3785), .B(n3792), .ZN(n3787) );
  OAI211_X1 U3675 ( .C1(n3951), .C2(n3813), .A(n3788), .B(n3787), .ZN(
        \CU_I/aluOpcode_i[0] ) );
  INV_X1 U3676 ( .A(n3795), .ZN(n3968) );
  NAND2_X1 U3677 ( .A1(n3968), .A2(IR_CU_27), .ZN(n3954) );
  NOR2_X1 U3678 ( .A1(IR_CU[1]), .A2(n478), .ZN(n3789) );
  AOI22_X1 U3679 ( .A1(IR_CU[1]), .A2(n478), .B1(n3789), .B2(n476), .ZN(n3803)
         );
  NOR3_X1 U3680 ( .A1(n3803), .A2(n3836), .A3(n3790), .ZN(n3791) );
  AOI21_X1 U3681 ( .B1(n3814), .B2(n3856), .A(n3791), .ZN(n3794) );
  NOR3_X1 U3682 ( .A1(IR_CU[1]), .A2(n478), .A3(n3802), .ZN(n3832) );
  NOR2_X1 U3683 ( .A1(n516), .A2(n510), .ZN(n3974) );
  NAND2_X1 U3684 ( .A1(n3976), .A2(n3974), .ZN(n3828) );
  AOI211_X1 U3685 ( .C1(n3832), .C2(n476), .A(n3792), .B(n3807), .ZN(n3793) );
  OAI211_X1 U3686 ( .C1(n514), .C2(n3954), .A(n3794), .B(n3793), .ZN(
        \CU_I/aluOpcode_i[1] ) );
  INV_X1 U3687 ( .A(n3966), .ZN(n3849) );
  NOR3_X1 U3688 ( .A1(n3795), .A2(n3955), .A3(n3849), .ZN(n3820) );
  NOR3_X1 U3689 ( .A1(n3795), .A2(n3837), .A3(n3977), .ZN(n3831) );
  INV_X1 U3690 ( .A(n3796), .ZN(n3799) );
  INV_X1 U3691 ( .A(n3797), .ZN(n3970) );
  OAI21_X1 U3692 ( .B1(n3799), .B2(n3970), .A(n3798), .ZN(n3800) );
  NOR4_X1 U3693 ( .A1(n3820), .A2(n3831), .A3(n3801), .A4(n3800), .ZN(n3812)
         );
  NOR3_X1 U3694 ( .A1(n3803), .A2(n3802), .A3(n480), .ZN(n3810) );
  NAND3_X1 U3695 ( .A1(n478), .A2(n3824), .A3(n476), .ZN(n3835) );
  NAND2_X1 U3696 ( .A1(n3804), .A2(IR_CU[0]), .ZN(n3805) );
  AOI211_X1 U3697 ( .C1(n3835), .C2(n3805), .A(IR_CU[1]), .B(n3836), .ZN(n3809) );
  NOR3_X1 U3698 ( .A1(IR_CU[4]), .A2(n477), .A3(n3806), .ZN(n3808) );
  NOR4_X1 U3699 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  OAI211_X1 U3700 ( .C1(n504), .C2(n3813), .A(n3812), .B(n3811), .ZN(
        \CU_I/aluOpcode_i[2] ) );
  AOI211_X1 U3701 ( .C1(IR_CU_31), .C2(n510), .A(n3977), .B(n3970), .ZN(n3819)
         );
  NAND2_X1 U3702 ( .A1(n3856), .A2(n3814), .ZN(n3816) );
  NAND2_X1 U3703 ( .A1(n606), .A2(n504), .ZN(n3815) );
  OAI211_X1 U3704 ( .C1(n3849), .C2(n3817), .A(n3816), .B(n3815), .ZN(n3818)
         );
  NOR4_X1 U3705 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3826)
         );
  OAI211_X1 U3706 ( .C1(n2128), .C2(n480), .A(IR_CU[5]), .B(IR_CU[0]), .ZN(
        n3822) );
  OAI21_X1 U3707 ( .B1(n478), .B2(n3836), .A(n3822), .ZN(n3823) );
  NAND3_X1 U3708 ( .A1(n3824), .A2(n477), .A3(n3823), .ZN(n3825) );
  OAI211_X1 U3709 ( .C1(n476), .C2(n3827), .A(n3826), .B(n3825), .ZN(
        \CU_I/aluOpcode_i[3] ) );
  OAI211_X1 U3710 ( .C1(n516), .C2(n2141), .A(n510), .B(n2129), .ZN(n3829) );
  AOI22_X1 U3711 ( .A1(IR_CU_27), .A2(n3829), .B1(n3828), .B2(n504), .ZN(n3830) );
  AOI211_X1 U3712 ( .C1(n3832), .C2(IR_CU[4]), .A(n3831), .B(n3830), .ZN(n3834) );
  OAI211_X1 U3713 ( .C1(n3836), .C2(n3835), .A(n3834), .B(n3833), .ZN(
        \CU_I/aluOpcode_i[4] ) );
  OAI211_X1 U3714 ( .C1(IR_CU_26), .C2(n2129), .A(IR_CU_28), .B(IR_CU_27), 
        .ZN(n3839) );
  NOR3_X1 U3715 ( .A1(n515), .A2(n510), .A3(n3837), .ZN(n3838) );
  AOI21_X1 U3716 ( .B1(n2141), .B2(n3839), .A(n3838), .ZN(n3857) );
  NOR3_X1 U3717 ( .A1(n515), .A2(n2141), .A3(n504), .ZN(n3859) );
  INV_X1 U3718 ( .A(n3845), .ZN(n3840) );
  AOI22_X1 U3719 ( .A1(IR_CU_28), .A2(n3859), .B1(n3856), .B2(n3840), .ZN(
        n3841) );
  AOI22_X1 U3720 ( .A1(IR_CU_28), .A2(IR_CU_27), .B1(n504), .B2(n510), .ZN(
        n3844) );
  NAND2_X1 U3721 ( .A1(n3976), .A2(n3844), .ZN(n3860) );
  OAI221_X1 U3722 ( .B1(IR_CU_31), .B2(n3857), .C1(IR_CU_31), .C2(n3841), .A(
        n3860), .ZN(n3846) );
  AOI21_X1 U3723 ( .B1(n3968), .B2(n3966), .A(n3846), .ZN(n1371) );
  AOI21_X1 U3724 ( .B1(IR_CU_26), .B2(n510), .A(n504), .ZN(n3843) );
  INV_X1 U3725 ( .A(n3955), .ZN(n3973) );
  NAND2_X1 U3726 ( .A1(IR_CU_31), .A2(n3973), .ZN(n3842) );
  OAI21_X1 U3727 ( .B1(n3843), .B2(n3842), .A(n1371), .ZN(\CU_I/cw[0] ) );
  AND3_X1 U3728 ( .A1(n3973), .A2(n3844), .A3(n516), .ZN(\CU_I/cw[10] ) );
  NOR2_X1 U3729 ( .A1(n516), .A2(n3845), .ZN(n3850) );
  AOI21_X1 U3730 ( .B1(n3951), .B2(n3850), .A(n3847), .ZN(n3862) );
  INV_X1 U3731 ( .A(n3862), .ZN(\CU_I/cw[6] ) );
  OR2_X1 U3732 ( .A1(n3846), .A2(\CU_I/cw[6] ), .ZN(\CU_I/cw[1] ) );
  NAND2_X1 U3733 ( .A1(n3850), .A2(n2141), .ZN(n3852) );
  AOI22_X1 U3734 ( .A1(n3850), .A2(n3856), .B1(n3847), .B2(n510), .ZN(n3848)
         );
  OAI21_X1 U3735 ( .B1(n3849), .B2(n3852), .A(n3848), .ZN(\CU_I/cw[3] ) );
  NAND2_X1 U3736 ( .A1(n3973), .A2(n3974), .ZN(n3854) );
  OAI211_X1 U3737 ( .C1(n2141), .C2(n497), .A(n3850), .B(n504), .ZN(n3851) );
  OAI21_X1 U3738 ( .B1(n3970), .B2(n3854), .A(n3851), .ZN(\CU_I/cw[4] ) );
  INV_X1 U3739 ( .A(n3854), .ZN(n3855) );
  AOI21_X1 U3740 ( .B1(n3856), .B2(n3855), .A(\CU_I/cw[7] ), .ZN(n1357) );
  INV_X1 U3741 ( .A(n3857), .ZN(n3858) );
  AOI221_X1 U3742 ( .B1(n3859), .B2(n516), .C1(n3858), .C2(n516), .A(
        \CU_I/cw[10] ), .ZN(n3861) );
  NAND3_X1 U3743 ( .A1(n3862), .A2(n3861), .A3(n3860), .ZN(\CU_I/cw[9] ) );
  NAND3_X1 U3744 ( .A1(n443), .A2(ALU_OPCODE_i[2]), .A3(ALU_OPCODE_i[1]), .ZN(
        n3903) );
  OR2_X1 U3745 ( .A1(n3903), .A2(ALU_OPCODE_i[0]), .ZN(n3984) );
  NOR4_X1 U3746 ( .A1(\DataP/alu_out_W[12] ), .A2(\DataP/alu_out_W[11] ), .A3(
        \DataP/alu_out_W[10] ), .A4(\DataP/alu_out_W[0] ), .ZN(n3866) );
  NOR4_X1 U3747 ( .A1(\DataP/alu_out_W[15] ), .A2(\DataP/alu_out_W[14] ), .A3(
        \DataP/alu_out_W[13] ), .A4(\DataP/alu_out_W[16] ), .ZN(n3865) );
  NOR4_X1 U3748 ( .A1(\DataP/alu_out_W[17] ), .A2(\DataP/alu_out_W[19] ), .A3(
        \DataP/alu_out_W[18] ), .A4(\DataP/alu_out_W[1] ), .ZN(n3864) );
  NOR4_X1 U3749 ( .A1(\DataP/alu_out_W[23] ), .A2(\DataP/alu_out_W[21] ), .A3(
        \DataP/alu_out_W[20] ), .A4(\DataP/alu_out_W[22] ), .ZN(n3863) );
  NAND4_X1 U3750 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3899)
         );
  INV_X1 U3751 ( .A(\DataP/FWD_MUX_BR_S[0] ), .ZN(n3871) );
  NAND2_X1 U3752 ( .A1(n3871), .A2(\DataP/FWD_MUX_BR_S[1] ), .ZN(n3880) );
  INV_X1 U3753 ( .A(n3880), .ZN(n3898) );
  NOR4_X1 U3754 ( .A1(\DataP/alu_out_W[27] ), .A2(\DataP/alu_out_W[26] ), .A3(
        \DataP/alu_out_W[25] ), .A4(\DataP/alu_out_W[24] ), .ZN(n3870) );
  NOR4_X1 U3755 ( .A1(\DataP/alu_out_W[30] ), .A2(\DataP/alu_out_W[29] ), .A3(
        \DataP/alu_out_W[28] ), .A4(\DataP/alu_out_W[2] ), .ZN(n3869) );
  NOR4_X1 U3756 ( .A1(\DataP/alu_out_W[31] ), .A2(\DataP/alu_out_W[5] ), .A3(
        \DataP/alu_out_W[4] ), .A4(\DataP/alu_out_W[3] ), .ZN(n3868) );
  NOR4_X1 U3757 ( .A1(\DataP/alu_out_W[9] ), .A2(\DataP/alu_out_W[8] ), .A3(
        \DataP/alu_out_W[7] ), .A4(\DataP/alu_out_W[6] ), .ZN(n3867) );
  NAND4_X1 U3758 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3897)
         );
  NOR2_X1 U3759 ( .A1(\DataP/FWD_MUX_BR_S[1] ), .A2(n3871), .ZN(n3895) );
  NOR4_X1 U3760 ( .A1(\DataP/A_s[27] ), .A2(\DataP/A_s[26] ), .A3(
        \DataP/A_s[25] ), .A4(\DataP/A_s[24] ), .ZN(n3875) );
  NOR4_X1 U3761 ( .A1(\DataP/A_s[30] ), .A2(\DataP/A_s[29] ), .A3(
        \DataP/A_s[28] ), .A4(\DataP/A_s[2] ), .ZN(n3874) );
  NOR4_X1 U3762 ( .A1(\DataP/A_s[31] ), .A2(\DataP/A_s[5] ), .A3(
        \DataP/A_s[4] ), .A4(\DataP/A_s[3] ), .ZN(n3873) );
  NOR4_X1 U3763 ( .A1(\DataP/A_s[9] ), .A2(\DataP/A_s[8] ), .A3(\DataP/A_s[7] ), .A4(\DataP/A_s[6] ), .ZN(n3872) );
  NAND4_X1 U3764 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3882)
         );
  NOR4_X1 U3765 ( .A1(\DataP/A_s[12] ), .A2(\DataP/A_s[11] ), .A3(
        \DataP/A_s[10] ), .A4(\DataP/A_s[0] ), .ZN(n3879) );
  NOR4_X1 U3766 ( .A1(\DataP/A_s[15] ), .A2(\DataP/A_s[14] ), .A3(
        \DataP/A_s[13] ), .A4(\DataP/A_s[16] ), .ZN(n3878) );
  NOR4_X1 U3767 ( .A1(\DataP/A_s[17] ), .A2(\DataP/A_s[19] ), .A3(
        \DataP/A_s[18] ), .A4(\DataP/A_s[1] ), .ZN(n3877) );
  NOR4_X1 U3768 ( .A1(\DataP/A_s[23] ), .A2(\DataP/A_s[21] ), .A3(
        \DataP/A_s[20] ), .A4(\DataP/A_s[22] ), .ZN(n3876) );
  NAND4_X1 U3769 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3881)
         );
  OAI21_X1 U3770 ( .B1(n3882), .B2(n3881), .A(n3880), .ZN(n3894) );
  NOR4_X1 U3771 ( .A1(DRAM_ADDRESS[11]), .A2(DRAM_ADDRESS[10]), .A3(
        DRAM_ADDRESS[1]), .A4(DRAM_ADDRESS[0]), .ZN(n3886) );
  NOR4_X1 U3772 ( .A1(DRAM_ADDRESS[5]), .A2(DRAM_ADDRESS[4]), .A3(
        DRAM_ADDRESS[3]), .A4(DRAM_ADDRESS[2]), .ZN(n3885) );
  NOR4_X1 U3773 ( .A1(DRAM_ADDRESS[9]), .A2(DRAM_ADDRESS[8]), .A3(
        DRAM_ADDRESS[7]), .A4(DRAM_ADDRESS[6]), .ZN(n3884) );
  NOR4_X1 U3774 ( .A1(\DataP/alu_out_M[15] ), .A2(\DataP/alu_out_M[14] ), .A3(
        \DataP/alu_out_M[13] ), .A4(\DataP/alu_out_M[12] ), .ZN(n3883) );
  NAND4_X1 U3775 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3892)
         );
  NOR4_X1 U3776 ( .A1(\DataP/alu_out_M[16] ), .A2(\DataP/alu_out_M[17] ), .A3(
        \DataP/alu_out_M[19] ), .A4(\DataP/alu_out_M[18] ), .ZN(n3890) );
  NOR4_X1 U3777 ( .A1(\DataP/alu_out_M[23] ), .A2(\DataP/alu_out_M[21] ), .A3(
        \DataP/alu_out_M[20] ), .A4(\DataP/alu_out_M[22] ), .ZN(n3889) );
  NOR4_X1 U3778 ( .A1(\DataP/alu_out_M[27] ), .A2(\DataP/alu_out_M[26] ), .A3(
        \DataP/alu_out_M[25] ), .A4(\DataP/alu_out_M[24] ), .ZN(n3888) );
  NOR4_X1 U3779 ( .A1(\DataP/alu_out_M[31] ), .A2(\DataP/alu_out_M[30] ), .A3(
        \DataP/alu_out_M[29] ), .A4(\DataP/alu_out_M[28] ), .ZN(n3887) );
  NAND4_X1 U3780 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  OAI21_X1 U3781 ( .B1(n3892), .B2(n3891), .A(n3895), .ZN(n3893) );
  OAI21_X1 U3782 ( .B1(n3895), .B2(n3894), .A(n3893), .ZN(n3896) );
  AOI221_X1 U3783 ( .B1(n3899), .B2(n3898), .C1(n3897), .C2(n3898), .A(n3896), 
        .ZN(n3900) );
  XNOR2_X1 U3784 ( .A(\DataP/pr_E ), .B(n3900), .ZN(n3983) );
  NAND2_X1 U3785 ( .A1(BR_EN_i), .A2(ALU_OPCODE_i[3]), .ZN(n3982) );
  NAND2_X1 U3786 ( .A1(ALU_OPCODE_i[1]), .A2(ALU_OPCODE_i[0]), .ZN(n3902) );
  INV_X1 U3787 ( .A(\DataP/npc[8] ), .ZN(n3998) );
  INV_X1 U3788 ( .A(\DataP/npc[9] ), .ZN(n3999) );
  OAI22_X1 U3789 ( .A1(n341), .A2(n3911), .B1(n3910), .B2(n3999), .ZN(
        \DataP/PC_reg/N11 ) );
  INV_X1 U3790 ( .A(\DataP/npc[10] ), .ZN(n4000) );
  OAI22_X1 U3791 ( .A1(n340), .A2(n3911), .B1(n3910), .B2(n4000), .ZN(
        \DataP/PC_reg/N12 ) );
  INV_X1 U3792 ( .A(\DataP/npc[11] ), .ZN(n4001) );
  OAI22_X1 U3793 ( .A1(n2137), .A2(n3911), .B1(n3910), .B2(n4001), .ZN(
        \DataP/PC_reg/N13 ) );
  INV_X1 U3794 ( .A(\DataP/npc[12] ), .ZN(n4002) );
  OAI22_X1 U3795 ( .A1(n337), .A2(n3911), .B1(n3910), .B2(n4002), .ZN(
        \DataP/PC_reg/N14 ) );
  NAND3_X1 U3796 ( .A1(n2222), .A2(n3907), .A3(n3906), .ZN(n3905) );
  INV_X1 U3797 ( .A(\DataP/npc[0] ), .ZN(n3990) );
  INV_X1 U3798 ( .A(\DataP/npc[1] ), .ZN(n3991) );
  OAI22_X1 U3799 ( .A1(n358), .A2(n3911), .B1(n3910), .B2(n3991), .ZN(
        \DataP/PC_reg/N3 ) );
  INV_X1 U3800 ( .A(\DataP/npc[2] ), .ZN(n3992) );
  OAI22_X1 U3801 ( .A1(n357), .A2(n3911), .B1(n3910), .B2(n3992), .ZN(
        \DataP/PC_reg/N4 ) );
  INV_X1 U3802 ( .A(\DataP/npc[3] ), .ZN(n3993) );
  INV_X1 U3803 ( .A(\DataP/npc[4] ), .ZN(n3994) );
  INV_X1 U3804 ( .A(\DataP/npc[5] ), .ZN(n3995) );
  OAI22_X1 U3805 ( .A1(n354), .A2(n3911), .B1(n3910), .B2(n3995), .ZN(
        \DataP/PC_reg/N7 ) );
  INV_X1 U3806 ( .A(\DataP/npc[6] ), .ZN(n3996) );
  INV_X1 U3807 ( .A(\DataP/npc[7] ), .ZN(n3997) );
  OAI22_X1 U3808 ( .A1(n350), .A2(n3911), .B1(n3910), .B2(n3997), .ZN(
        \DataP/PC_reg/N9 ) );
  AOI22_X1 U3809 ( .A1(n3008), .A2(\DataP/LMD_out[0] ), .B1(n3943), .B2(
        \DataP/link_addr_W[0] ), .ZN(n3912) );
  OAI21_X1 U3810 ( .B1(n2272), .B2(n3946), .A(n3912), .ZN(\DataP/WB[0] ) );
  AOI22_X1 U3811 ( .A1(n3008), .A2(\DataP/LMD_out[10] ), .B1(n3943), .B2(
        \DataP/link_addr_W[10] ), .ZN(n3913) );
  OAI21_X1 U3812 ( .B1(n2257), .B2(n3946), .A(n3913), .ZN(\DataP/WB[10] ) );
  AOI22_X1 U3813 ( .A1(n3008), .A2(\DataP/LMD_out[11] ), .B1(n3943), .B2(
        \DataP/link_addr_W[11] ), .ZN(n3914) );
  OAI21_X1 U3814 ( .B1(n2251), .B2(n3946), .A(n3914), .ZN(\DataP/WB[11] ) );
  AOI22_X1 U3815 ( .A1(n3008), .A2(\DataP/LMD_out[12] ), .B1(n3943), .B2(
        \DataP/link_addr_W[12] ), .ZN(n3915) );
  OAI21_X1 U3816 ( .B1(n2246), .B2(n3946), .A(n3915), .ZN(\DataP/WB[12] ) );
  AOI22_X1 U3817 ( .A1(n3008), .A2(\DataP/LMD_out[13] ), .B1(n3943), .B2(
        \DataP/link_addr_W[13] ), .ZN(n3916) );
  OAI21_X1 U3818 ( .B1(n2258), .B2(n3946), .A(n3916), .ZN(\DataP/WB[13] ) );
  AOI22_X1 U3819 ( .A1(n3008), .A2(\DataP/LMD_out[14] ), .B1(n3943), .B2(
        \DataP/link_addr_W[14] ), .ZN(n3917) );
  OAI21_X1 U3820 ( .B1(n2252), .B2(n3946), .A(n3917), .ZN(\DataP/WB[14] ) );
  AOI22_X1 U3821 ( .A1(n3008), .A2(\DataP/LMD_out[15] ), .B1(n3943), .B2(
        \DataP/link_addr_W[15] ), .ZN(n3918) );
  OAI21_X1 U3822 ( .B1(n2247), .B2(n3946), .A(n3918), .ZN(\DataP/WB[15] ) );
  AOI22_X1 U3823 ( .A1(n3008), .A2(\DataP/LMD_out[16] ), .B1(n3943), .B2(
        \DataP/link_addr_W[16] ), .ZN(n3919) );
  OAI21_X1 U3824 ( .B1(n2263), .B2(n3946), .A(n3919), .ZN(\DataP/WB[16] ) );
  AOI22_X1 U3825 ( .A1(n3944), .A2(\DataP/LMD_out[17] ), .B1(n3943), .B2(
        \DataP/link_addr_W[17] ), .ZN(n3920) );
  OAI21_X1 U3826 ( .B1(n2248), .B2(n3946), .A(n3920), .ZN(\DataP/WB[17] ) );
  AOI22_X1 U3827 ( .A1(n3944), .A2(\DataP/LMD_out[18] ), .B1(n3943), .B2(
        \DataP/link_addr_W[18] ), .ZN(n3921) );
  OAI21_X1 U3828 ( .B1(n2259), .B2(n3946), .A(n3921), .ZN(\DataP/WB[18] ) );
  AOI22_X1 U3829 ( .A1(n3008), .A2(\DataP/LMD_out[19] ), .B1(n3943), .B2(
        \DataP/link_addr_W[19] ), .ZN(n3922) );
  OAI21_X1 U3830 ( .B1(n2253), .B2(n3946), .A(n3922), .ZN(\DataP/WB[19] ) );
  AOI22_X1 U3831 ( .A1(n3008), .A2(\DataP/LMD_out[1] ), .B1(n3943), .B2(
        \DataP/link_addr_W[1] ), .ZN(n3923) );
  OAI21_X1 U3832 ( .B1(n2273), .B2(n3946), .A(n3923), .ZN(\DataP/WB[1] ) );
  AOI22_X1 U3833 ( .A1(n3008), .A2(\DataP/LMD_out[20] ), .B1(n3943), .B2(
        \DataP/link_addr_W[20] ), .ZN(n3924) );
  OAI21_X1 U3834 ( .B1(n2260), .B2(n3946), .A(n3924), .ZN(\DataP/WB[20] ) );
  AOI22_X1 U3835 ( .A1(n3008), .A2(\DataP/LMD_out[21] ), .B1(n3943), .B2(
        \DataP/link_addr_W[21] ), .ZN(n3925) );
  OAI21_X1 U3836 ( .B1(n2254), .B2(n3946), .A(n3925), .ZN(\DataP/WB[21] ) );
  AOI22_X1 U3837 ( .A1(n3008), .A2(\DataP/LMD_out[22] ), .B1(n3943), .B2(
        \DataP/link_addr_W[22] ), .ZN(n3926) );
  OAI21_X1 U3838 ( .B1(n2264), .B2(n3946), .A(n3926), .ZN(\DataP/WB[22] ) );
  AOI22_X1 U3839 ( .A1(n3008), .A2(\DataP/LMD_out[23] ), .B1(n3943), .B2(
        \DataP/link_addr_W[23] ), .ZN(n3927) );
  OAI21_X1 U3840 ( .B1(n2249), .B2(n3946), .A(n3927), .ZN(\DataP/WB[23] ) );
  AOI22_X1 U3841 ( .A1(n3008), .A2(\DataP/LMD_out[24] ), .B1(n3943), .B2(
        \DataP/link_addr_W[24] ), .ZN(n3928) );
  OAI21_X1 U3842 ( .B1(n2265), .B2(n3946), .A(n3928), .ZN(\DataP/WB[24] ) );
  AOI22_X1 U3843 ( .A1(n3008), .A2(\DataP/LMD_out[25] ), .B1(n3943), .B2(
        \DataP/link_addr_W[25] ), .ZN(n3929) );
  OAI21_X1 U3844 ( .B1(n2261), .B2(n3946), .A(n3929), .ZN(\DataP/WB[25] ) );
  AOI22_X1 U3845 ( .A1(n3008), .A2(\DataP/LMD_out[26] ), .B1(n3943), .B2(
        \DataP/link_addr_W[26] ), .ZN(n3930) );
  OAI21_X1 U3846 ( .B1(n2255), .B2(n3946), .A(n3930), .ZN(\DataP/WB[26] ) );
  AOI22_X1 U3847 ( .A1(n3008), .A2(\DataP/LMD_out[27] ), .B1(n3943), .B2(
        \DataP/link_addr_W[27] ), .ZN(n3931) );
  OAI21_X1 U3848 ( .B1(n2250), .B2(n3946), .A(n3931), .ZN(\DataP/WB[27] ) );
  AOI22_X1 U3849 ( .A1(n3944), .A2(\DataP/LMD_out[28] ), .B1(n3943), .B2(
        \DataP/link_addr_W[28] ), .ZN(n3932) );
  OAI21_X1 U3850 ( .B1(n2262), .B2(n3946), .A(n3932), .ZN(\DataP/WB[28] ) );
  AOI22_X1 U3851 ( .A1(n3944), .A2(\DataP/LMD_out[29] ), .B1(n3943), .B2(
        \DataP/link_addr_W[29] ), .ZN(n3933) );
  OAI21_X1 U3852 ( .B1(n2256), .B2(n3946), .A(n3933), .ZN(\DataP/WB[29] ) );
  AOI22_X1 U3853 ( .A1(n3944), .A2(\DataP/LMD_out[2] ), .B1(n3943), .B2(
        \DataP/link_addr_W[2] ), .ZN(n3934) );
  OAI21_X1 U3854 ( .B1(n2276), .B2(n3946), .A(n3934), .ZN(\DataP/WB[2] ) );
  AOI22_X1 U3855 ( .A1(n3944), .A2(\DataP/LMD_out[30] ), .B1(n3943), .B2(
        \DataP/link_addr_W[30] ), .ZN(n3935) );
  OAI21_X1 U3856 ( .B1(n2266), .B2(n3946), .A(n3935), .ZN(\DataP/WB[30] ) );
  AOI22_X1 U3857 ( .A1(n3944), .A2(\DataP/LMD_out[31] ), .B1(n3943), .B2(
        \DataP/link_addr_W[31] ), .ZN(n3936) );
  OAI21_X1 U3858 ( .B1(n2267), .B2(n3946), .A(n3936), .ZN(\DataP/WB[31] ) );
  AOI22_X1 U3859 ( .A1(n3944), .A2(\DataP/LMD_out[3] ), .B1(n3943), .B2(
        \DataP/link_addr_W[3] ), .ZN(n3937) );
  OAI21_X1 U3860 ( .B1(n2277), .B2(n3946), .A(n3937), .ZN(\DataP/WB[3] ) );
  AOI22_X1 U3861 ( .A1(n3944), .A2(\DataP/LMD_out[4] ), .B1(n3943), .B2(
        \DataP/link_addr_W[4] ), .ZN(n3938) );
  OAI21_X1 U3862 ( .B1(n2274), .B2(n3946), .A(n3938), .ZN(\DataP/WB[4] ) );
  AOI22_X1 U3863 ( .A1(n3008), .A2(\DataP/LMD_out[5] ), .B1(n3943), .B2(
        \DataP/link_addr_W[5] ), .ZN(n3939) );
  OAI21_X1 U3864 ( .B1(n2270), .B2(n3946), .A(n3939), .ZN(\DataP/WB[5] ) );
  AOI22_X1 U3865 ( .A1(n3944), .A2(\DataP/LMD_out[6] ), .B1(n3943), .B2(
        \DataP/link_addr_W[6] ), .ZN(n3940) );
  OAI21_X1 U3866 ( .B1(n2268), .B2(n3946), .A(n3940), .ZN(\DataP/WB[6] ) );
  AOI22_X1 U3867 ( .A1(n3008), .A2(\DataP/LMD_out[7] ), .B1(n3943), .B2(
        \DataP/link_addr_W[7] ), .ZN(n3941) );
  OAI21_X1 U3868 ( .B1(n2275), .B2(n3946), .A(n3941), .ZN(\DataP/WB[7] ) );
  AOI22_X1 U3869 ( .A1(n3944), .A2(\DataP/LMD_out[8] ), .B1(n3943), .B2(
        \DataP/link_addr_W[8] ), .ZN(n3942) );
  OAI21_X1 U3870 ( .B1(n2271), .B2(n3946), .A(n3942), .ZN(\DataP/WB[8] ) );
  AOI22_X1 U3871 ( .A1(n3008), .A2(\DataP/LMD_out[9] ), .B1(n3943), .B2(
        \DataP/link_addr_W[9] ), .ZN(n3945) );
  OAI21_X1 U3872 ( .B1(n2269), .B2(n3946), .A(n3945), .ZN(\DataP/WB[9] ) );
  INV_X1 U3873 ( .A(n144), .ZN(n3952) );
  AOI211_X1 U3874 ( .C1(n606), .C2(n504), .A(\CU_I/cw[7] ), .B(n3953), .ZN(
        n3950) );
  OAI211_X1 U3875 ( .C1(n3952), .C2(n3951), .A(Rst), .B(n3950), .ZN(n3964) );
  AND2_X1 U3876 ( .A1(Rst), .A2(n3953), .ZN(n3962) );
  NOR2_X1 U3877 ( .A1(n3955), .A2(n3954), .ZN(n3965) );
  NAND2_X1 U3878 ( .A1(Rst), .A2(n3965), .ZN(n3979) );
  OAI22_X1 U3879 ( .A1(n497), .A2(n3979), .B1(n3956), .B2(n3964), .ZN(n3961)
         );
  AOI21_X1 U3880 ( .B1(n3962), .B2(\DataP/IR1[11] ), .A(n3961), .ZN(n3957) );
  OAI21_X1 U3881 ( .B1(n485), .B2(n3964), .A(n3957), .ZN(\DataP/dest_D[0] ) );
  AOI21_X1 U3882 ( .B1(n3962), .B2(\DataP/IR1[12] ), .A(n3961), .ZN(n3958) );
  OAI21_X1 U3883 ( .B1(n486), .B2(n3964), .A(n3958), .ZN(\DataP/dest_D[1] ) );
  AOI21_X1 U3884 ( .B1(n3962), .B2(\DataP/IR1[13] ), .A(n3961), .ZN(n3959) );
  OAI21_X1 U3885 ( .B1(n487), .B2(n3964), .A(n3959), .ZN(\DataP/dest_D[2] ) );
  AOI21_X1 U3886 ( .B1(n3962), .B2(\DataP/IR1[14] ), .A(n3961), .ZN(n3960) );
  OAI21_X1 U3887 ( .B1(n488), .B2(n3964), .A(n3960), .ZN(\DataP/dest_D[3] ) );
  AOI21_X1 U3888 ( .B1(n3962), .B2(\DataP/IR1[15] ), .A(n3961), .ZN(n3963) );
  OAI21_X1 U3889 ( .B1(n489), .B2(n3964), .A(n3963), .ZN(\DataP/dest_D[4] ) );
  NAND2_X1 U3890 ( .A1(IR_CU_28), .A2(n3966), .ZN(n3971) );
  OAI21_X1 U3891 ( .B1(n515), .B2(IR_CU_27), .A(n2141), .ZN(n3967) );
  AOI22_X1 U3892 ( .A1(n3968), .A2(n497), .B1(n510), .B2(n3967), .ZN(n3969) );
  OAI221_X1 U3893 ( .B1(n514), .B2(n3971), .C1(n2141), .C2(n3970), .A(n3969), 
        .ZN(n3972) );
  AOI211_X1 U3894 ( .C1(IR_CU_27), .C2(n3974), .A(n3973), .B(n3972), .ZN(n3975) );
  OAI221_X1 U3895 ( .B1(IR_CU_31), .B2(n3977), .C1(n516), .C2(n3976), .A(n3975), .ZN(n3978) );
  NAND4_X1 U3896 ( .A1(Rst), .A2(\DataP/IR1[15] ), .A3(n3981), .A4(n3978), 
        .ZN(n3980) );
  OAI21_X1 U3897 ( .B1(n485), .B2(n3979), .A(n3980), .ZN(\DataP/imm_out[16] )
         );
  OAI21_X1 U3898 ( .B1(n486), .B2(n3979), .A(n3980), .ZN(\DataP/imm_out[17] )
         );
  OAI21_X1 U3899 ( .B1(n487), .B2(n3979), .A(n3980), .ZN(\DataP/imm_out[18] )
         );
  OAI21_X1 U3900 ( .B1(n488), .B2(n3979), .A(n3980), .ZN(\DataP/imm_out[19] )
         );
  OAI21_X1 U3901 ( .B1(n489), .B2(n3979), .A(n3980), .ZN(\DataP/imm_out[20] )
         );
  NAND2_X1 U3902 ( .A1(Rst), .A2(\DataP/IR1[21] ), .ZN(n3989) );
  OAI21_X1 U3903 ( .B1(n3981), .B2(n3989), .A(n3980), .ZN(\DataP/imm_out[21] )
         );
  NAND2_X1 U3904 ( .A1(Rst), .A2(\DataP/IR1[22] ), .ZN(n3988) );
  OAI21_X1 U3905 ( .B1(n3981), .B2(n3988), .A(n3980), .ZN(\DataP/imm_out[22] )
         );
  NAND2_X1 U3906 ( .A1(Rst), .A2(\DataP/IR1[23] ), .ZN(n3987) );
  OAI21_X1 U3907 ( .B1(n3981), .B2(n3987), .A(n3980), .ZN(\DataP/imm_out[23] )
         );
  NAND2_X1 U3908 ( .A1(Rst), .A2(\DataP/IR1[24] ), .ZN(n3986) );
  OAI21_X1 U3909 ( .B1(n3981), .B2(n3986), .A(n3980), .ZN(\DataP/imm_out[24] )
         );
  NAND2_X1 U3910 ( .A1(Rst), .A2(\DataP/IR1[25] ), .ZN(n3985) );
  OAI21_X1 U3911 ( .B1(n3981), .B2(n3985), .A(n3980), .ZN(\DataP/imm_out[31] )
         );
  MUX2_X1 U3912 ( .A(\DataP/pc_out_0 ), .B(\DataP/npc_pre[0] ), .S(n1940), .Z(
        \DataP/NPC_add/N1 ) );
  MUX2_X1 U3913 ( .A(\DataP/pc_out_1 ), .B(\DataP/npc_pre[1] ), .S(n1940), .Z(
        \DataP/NPC_add/N2 ) );
  NAND2_X1 U3914 ( .A1(\DataP/npc[0] ), .A2(n3009), .ZN(n127) );
  AOI21_X1 U3915 ( .B1(n3990), .B2(n4022), .A(n3013), .ZN(n126) );
  NAND2_X1 U3916 ( .A1(\DataP/npc[1] ), .A2(n4021), .ZN(n123) );
  AOI21_X1 U3917 ( .B1(n3991), .B2(n4022), .A(n3013), .ZN(n122) );
  NAND2_X1 U3918 ( .A1(\DataP/npc[2] ), .A2(n3009), .ZN(n119) );
  AOI21_X1 U3919 ( .B1(n3992), .B2(n4022), .A(n3013), .ZN(n118) );
  NAND2_X1 U3920 ( .A1(\DataP/npc[3] ), .A2(n4021), .ZN(n115) );
  AOI21_X1 U3921 ( .B1(n3993), .B2(n4022), .A(n3013), .ZN(n114) );
  NAND2_X1 U3922 ( .A1(\DataP/npc[4] ), .A2(n3009), .ZN(n111) );
  AOI21_X1 U3923 ( .B1(n3994), .B2(n4022), .A(n3013), .ZN(n110) );
  NAND2_X1 U3924 ( .A1(\DataP/npc[5] ), .A2(n4021), .ZN(n107) );
  AOI21_X1 U3925 ( .B1(n3995), .B2(n4022), .A(n3013), .ZN(n106) );
  NAND2_X1 U3926 ( .A1(\DataP/npc[6] ), .A2(n4021), .ZN(n103) );
  AOI21_X1 U3927 ( .B1(n3996), .B2(n4022), .A(n3013), .ZN(n102) );
  NAND2_X1 U3928 ( .A1(\DataP/npc[7] ), .A2(n4021), .ZN(n99) );
  AOI21_X1 U3929 ( .B1(n3997), .B2(n4022), .A(n3013), .ZN(n98) );
  NAND2_X1 U3930 ( .A1(\DataP/npc[8] ), .A2(n4021), .ZN(n95) );
  AOI21_X1 U3931 ( .B1(n3998), .B2(n4022), .A(n3013), .ZN(n94) );
  NAND2_X1 U3932 ( .A1(\DataP/npc[9] ), .A2(n4021), .ZN(n91) );
  AOI21_X1 U3933 ( .B1(n3999), .B2(n4022), .A(n3013), .ZN(n90) );
  NAND2_X1 U3934 ( .A1(\DataP/npc[10] ), .A2(n4021), .ZN(n87) );
  AOI21_X1 U3935 ( .B1(n4000), .B2(n4022), .A(n3014), .ZN(n86) );
  NAND2_X1 U3936 ( .A1(\DataP/npc[11] ), .A2(n4021), .ZN(n83) );
  AOI21_X1 U3937 ( .B1(n4001), .B2(n4022), .A(n3013), .ZN(n82) );
  NAND2_X1 U3938 ( .A1(\DataP/npc[12] ), .A2(n3009), .ZN(n79) );
  AOI21_X1 U3939 ( .B1(n4002), .B2(n4022), .A(n3013), .ZN(n78) );
  NAND2_X1 U3940 ( .A1(\DataP/npc[13] ), .A2(n3009), .ZN(n75) );
  AOI21_X1 U3941 ( .B1(n4003), .B2(n4022), .A(n3013), .ZN(n74) );
  NAND2_X1 U3942 ( .A1(\DataP/npc[14] ), .A2(n3009), .ZN(n71) );
  AOI21_X1 U3943 ( .B1(n4004), .B2(n4022), .A(n3013), .ZN(n70) );
  NAND2_X1 U3944 ( .A1(\DataP/npc[15] ), .A2(n3009), .ZN(n67) );
  AOI21_X1 U3945 ( .B1(n4005), .B2(n4022), .A(n3014), .ZN(n66) );
  NAND2_X1 U3946 ( .A1(\DataP/npc[16] ), .A2(n3009), .ZN(n63) );
  AOI21_X1 U3947 ( .B1(n4006), .B2(n4022), .A(n3014), .ZN(n62) );
  NAND2_X1 U3948 ( .A1(\DataP/npc[17] ), .A2(n3009), .ZN(n59) );
  AOI21_X1 U3949 ( .B1(n4007), .B2(n4022), .A(n3014), .ZN(n58) );
  NAND2_X1 U3950 ( .A1(\DataP/npc[18] ), .A2(n3009), .ZN(n55) );
  AOI21_X1 U3951 ( .B1(n4008), .B2(n4022), .A(n3014), .ZN(n54) );
  NAND2_X1 U3952 ( .A1(\DataP/npc[19] ), .A2(n3009), .ZN(n51) );
  AOI21_X1 U3953 ( .B1(n4009), .B2(n4022), .A(n3014), .ZN(n50) );
  NAND2_X1 U3954 ( .A1(\DataP/npc[20] ), .A2(n3009), .ZN(n47) );
  AOI21_X1 U3955 ( .B1(n4010), .B2(n4022), .A(n3014), .ZN(n46) );
  NAND2_X1 U3956 ( .A1(\DataP/npc[21] ), .A2(n3009), .ZN(n43) );
  AOI21_X1 U3957 ( .B1(n4011), .B2(n4022), .A(n3014), .ZN(n42) );
  NAND2_X1 U3958 ( .A1(\DataP/npc[22] ), .A2(n4021), .ZN(n39) );
  AOI21_X1 U3959 ( .B1(n4012), .B2(n4022), .A(n3014), .ZN(n38) );
  NAND2_X1 U3960 ( .A1(\DataP/npc[23] ), .A2(n4021), .ZN(n35) );
  AOI21_X1 U3961 ( .B1(n4013), .B2(n4022), .A(n3014), .ZN(n34) );
  NAND2_X1 U3962 ( .A1(\DataP/npc[24] ), .A2(n3009), .ZN(n31) );
  AOI21_X1 U3963 ( .B1(n4014), .B2(n4022), .A(n3014), .ZN(n30) );
  NAND2_X1 U3964 ( .A1(\DataP/npc[25] ), .A2(n3009), .ZN(n27) );
  AOI21_X1 U3965 ( .B1(n4015), .B2(n4022), .A(n3014), .ZN(n26) );
  NAND2_X1 U3966 ( .A1(\DataP/npc[26] ), .A2(n3009), .ZN(n23) );
  AOI21_X1 U3967 ( .B1(n4016), .B2(n4022), .A(n3014), .ZN(n22) );
  NAND2_X1 U3968 ( .A1(\DataP/npc[27] ), .A2(n3009), .ZN(n19) );
  AOI21_X1 U3969 ( .B1(n4017), .B2(n4022), .A(n3014), .ZN(n18) );
  NAND2_X1 U3970 ( .A1(\DataP/npc[28] ), .A2(n3009), .ZN(n15) );
  AOI21_X1 U3971 ( .B1(n4018), .B2(n4022), .A(n3014), .ZN(n14) );
  NAND2_X1 U3972 ( .A1(\DataP/npc[29] ), .A2(n3009), .ZN(n11) );
  AOI21_X1 U3973 ( .B1(n4019), .B2(n4022), .A(n3014), .ZN(n10) );
  NAND2_X1 U3974 ( .A1(\DataP/npc[30] ), .A2(n3009), .ZN(n7) );
  AOI21_X1 U3975 ( .B1(n4020), .B2(n4022), .A(n3014), .ZN(n6) );
  NAND2_X1 U3976 ( .A1(\DataP/npc[31] ), .A2(n3009), .ZN(n3) );
  AOI21_X1 U3977 ( .B1(n4023), .B2(n4022), .A(n3013), .ZN(n2) );
endmodule

